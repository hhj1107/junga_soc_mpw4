magic
tech sky130A
magscale 1 2
timestamp 1640419346
<< obsli1 >>
rect 1104 629 163731 164305
<< obsm1 >>
rect 382 8 164022 164336
<< metal2 >>
rect 386 165957 442 166757
rect 1214 165957 1270 166757
rect 2134 165957 2190 166757
rect 3054 165957 3110 166757
rect 3974 165957 4030 166757
rect 4894 165957 4950 166757
rect 5814 165957 5870 166757
rect 6734 165957 6790 166757
rect 7654 165957 7710 166757
rect 8574 165957 8630 166757
rect 9494 165957 9550 166757
rect 10414 165957 10470 166757
rect 11334 165957 11390 166757
rect 12254 165957 12310 166757
rect 13174 165957 13230 166757
rect 14094 165957 14150 166757
rect 15014 165957 15070 166757
rect 15934 165957 15990 166757
rect 16854 165957 16910 166757
rect 17774 165957 17830 166757
rect 18694 165957 18750 166757
rect 19614 165957 19670 166757
rect 20534 165957 20590 166757
rect 21454 165957 21510 166757
rect 22374 165957 22430 166757
rect 23294 165957 23350 166757
rect 24214 165957 24270 166757
rect 25134 165957 25190 166757
rect 26054 165957 26110 166757
rect 26974 165957 27030 166757
rect 27894 165957 27950 166757
rect 28814 165957 28870 166757
rect 29734 165957 29790 166757
rect 30654 165957 30710 166757
rect 31574 165957 31630 166757
rect 32494 165957 32550 166757
rect 33414 165957 33470 166757
rect 34334 165957 34390 166757
rect 35254 165957 35310 166757
rect 36174 165957 36230 166757
rect 37094 165957 37150 166757
rect 38014 165957 38070 166757
rect 38934 165957 38990 166757
rect 39854 165957 39910 166757
rect 40774 165957 40830 166757
rect 41694 165957 41750 166757
rect 42614 165957 42670 166757
rect 43534 165957 43590 166757
rect 44454 165957 44510 166757
rect 45374 165957 45430 166757
rect 46294 165957 46350 166757
rect 47214 165957 47270 166757
rect 48134 165957 48190 166757
rect 49054 165957 49110 166757
rect 49974 165957 50030 166757
rect 50894 165957 50950 166757
rect 51814 165957 51870 166757
rect 52734 165957 52790 166757
rect 53654 165957 53710 166757
rect 54574 165957 54630 166757
rect 55494 165957 55550 166757
rect 56414 165957 56470 166757
rect 57334 165957 57390 166757
rect 58254 165957 58310 166757
rect 59174 165957 59230 166757
rect 60094 165957 60150 166757
rect 61014 165957 61070 166757
rect 61934 165957 61990 166757
rect 62854 165957 62910 166757
rect 63774 165957 63830 166757
rect 64694 165957 64750 166757
rect 65614 165957 65670 166757
rect 66534 165957 66590 166757
rect 67454 165957 67510 166757
rect 68374 165957 68430 166757
rect 69294 165957 69350 166757
rect 70214 165957 70270 166757
rect 71134 165957 71190 166757
rect 72054 165957 72110 166757
rect 72974 165957 73030 166757
rect 73894 165957 73950 166757
rect 74814 165957 74870 166757
rect 75734 165957 75790 166757
rect 76654 165957 76710 166757
rect 77574 165957 77630 166757
rect 78494 165957 78550 166757
rect 79414 165957 79470 166757
rect 80334 165957 80390 166757
rect 81254 165957 81310 166757
rect 82174 165957 82230 166757
rect 83094 165957 83150 166757
rect 84014 165957 84070 166757
rect 84934 165957 84990 166757
rect 85854 165957 85910 166757
rect 86774 165957 86830 166757
rect 87694 165957 87750 166757
rect 88614 165957 88670 166757
rect 89534 165957 89590 166757
rect 90454 165957 90510 166757
rect 91374 165957 91430 166757
rect 92294 165957 92350 166757
rect 93214 165957 93270 166757
rect 94134 165957 94190 166757
rect 95054 165957 95110 166757
rect 95974 165957 96030 166757
rect 96894 165957 96950 166757
rect 97814 165957 97870 166757
rect 98734 165957 98790 166757
rect 99654 165957 99710 166757
rect 100574 165957 100630 166757
rect 101494 165957 101550 166757
rect 102414 165957 102470 166757
rect 103334 165957 103390 166757
rect 104254 165957 104310 166757
rect 105174 165957 105230 166757
rect 106094 165957 106150 166757
rect 107014 165957 107070 166757
rect 107934 165957 107990 166757
rect 108854 165957 108910 166757
rect 109774 165957 109830 166757
rect 110694 165957 110750 166757
rect 111614 165957 111670 166757
rect 112534 165957 112590 166757
rect 113454 165957 113510 166757
rect 114374 165957 114430 166757
rect 115294 165957 115350 166757
rect 116214 165957 116270 166757
rect 117134 165957 117190 166757
rect 118054 165957 118110 166757
rect 118974 165957 119030 166757
rect 119894 165957 119950 166757
rect 120814 165957 120870 166757
rect 121734 165957 121790 166757
rect 122654 165957 122710 166757
rect 123574 165957 123630 166757
rect 124494 165957 124550 166757
rect 125414 165957 125470 166757
rect 126334 165957 126390 166757
rect 127254 165957 127310 166757
rect 128174 165957 128230 166757
rect 129094 165957 129150 166757
rect 130014 165957 130070 166757
rect 130934 165957 130990 166757
rect 131854 165957 131910 166757
rect 132774 165957 132830 166757
rect 133694 165957 133750 166757
rect 134614 165957 134670 166757
rect 135534 165957 135590 166757
rect 136454 165957 136510 166757
rect 137374 165957 137430 166757
rect 138294 165957 138350 166757
rect 139214 165957 139270 166757
rect 140134 165957 140190 166757
rect 141054 165957 141110 166757
rect 141974 165957 142030 166757
rect 142894 165957 142950 166757
rect 143814 165957 143870 166757
rect 144734 165957 144790 166757
rect 145654 165957 145710 166757
rect 146574 165957 146630 166757
rect 147494 165957 147550 166757
rect 148414 165957 148470 166757
rect 149334 165957 149390 166757
rect 150254 165957 150310 166757
rect 151174 165957 151230 166757
rect 152094 165957 152150 166757
rect 153014 165957 153070 166757
rect 153934 165957 153990 166757
rect 154854 165957 154910 166757
rect 155774 165957 155830 166757
rect 156694 165957 156750 166757
rect 157614 165957 157670 166757
rect 158534 165957 158590 166757
rect 159454 165957 159510 166757
rect 160374 165957 160430 166757
rect 161294 165957 161350 166757
rect 162214 165957 162270 166757
rect 163134 165957 163190 166757
rect 164054 165957 164110 166757
rect 478 0 534 800
rect 1490 0 1546 800
rect 2502 0 2558 800
rect 3514 0 3570 800
rect 4526 0 4582 800
rect 5538 0 5594 800
rect 6642 0 6698 800
rect 7654 0 7710 800
rect 8666 0 8722 800
rect 9678 0 9734 800
rect 10690 0 10746 800
rect 11702 0 11758 800
rect 12806 0 12862 800
rect 13818 0 13874 800
rect 14830 0 14886 800
rect 15842 0 15898 800
rect 16854 0 16910 800
rect 17958 0 18014 800
rect 18970 0 19026 800
rect 19982 0 20038 800
rect 20994 0 21050 800
rect 22006 0 22062 800
rect 23018 0 23074 800
rect 24122 0 24178 800
rect 25134 0 25190 800
rect 26146 0 26202 800
rect 27158 0 27214 800
rect 28170 0 28226 800
rect 29274 0 29330 800
rect 30286 0 30342 800
rect 31298 0 31354 800
rect 32310 0 32366 800
rect 33322 0 33378 800
rect 34334 0 34390 800
rect 35438 0 35494 800
rect 36450 0 36506 800
rect 37462 0 37518 800
rect 38474 0 38530 800
rect 39486 0 39542 800
rect 40590 0 40646 800
rect 41602 0 41658 800
rect 42614 0 42670 800
rect 43626 0 43682 800
rect 44638 0 44694 800
rect 45650 0 45706 800
rect 46754 0 46810 800
rect 47766 0 47822 800
rect 48778 0 48834 800
rect 49790 0 49846 800
rect 50802 0 50858 800
rect 51906 0 51962 800
rect 52918 0 52974 800
rect 53930 0 53986 800
rect 54942 0 54998 800
rect 55954 0 56010 800
rect 56966 0 57022 800
rect 58070 0 58126 800
rect 59082 0 59138 800
rect 60094 0 60150 800
rect 61106 0 61162 800
rect 62118 0 62174 800
rect 63222 0 63278 800
rect 64234 0 64290 800
rect 65246 0 65302 800
rect 66258 0 66314 800
rect 67270 0 67326 800
rect 68282 0 68338 800
rect 69386 0 69442 800
rect 70398 0 70454 800
rect 71410 0 71466 800
rect 72422 0 72478 800
rect 73434 0 73490 800
rect 74538 0 74594 800
rect 75550 0 75606 800
rect 76562 0 76618 800
rect 77574 0 77630 800
rect 78586 0 78642 800
rect 79598 0 79654 800
rect 80702 0 80758 800
rect 81714 0 81770 800
rect 82726 0 82782 800
rect 83738 0 83794 800
rect 84750 0 84806 800
rect 85854 0 85910 800
rect 86866 0 86922 800
rect 87878 0 87934 800
rect 88890 0 88946 800
rect 89902 0 89958 800
rect 90914 0 90970 800
rect 92018 0 92074 800
rect 93030 0 93086 800
rect 94042 0 94098 800
rect 95054 0 95110 800
rect 96066 0 96122 800
rect 97170 0 97226 800
rect 98182 0 98238 800
rect 99194 0 99250 800
rect 100206 0 100262 800
rect 101218 0 101274 800
rect 102230 0 102286 800
rect 103334 0 103390 800
rect 104346 0 104402 800
rect 105358 0 105414 800
rect 106370 0 106426 800
rect 107382 0 107438 800
rect 108486 0 108542 800
rect 109498 0 109554 800
rect 110510 0 110566 800
rect 111522 0 111578 800
rect 112534 0 112590 800
rect 113546 0 113602 800
rect 114650 0 114706 800
rect 115662 0 115718 800
rect 116674 0 116730 800
rect 117686 0 117742 800
rect 118698 0 118754 800
rect 119802 0 119858 800
rect 120814 0 120870 800
rect 121826 0 121882 800
rect 122838 0 122894 800
rect 123850 0 123906 800
rect 124862 0 124918 800
rect 125966 0 126022 800
rect 126978 0 127034 800
rect 127990 0 128046 800
rect 129002 0 129058 800
rect 130014 0 130070 800
rect 131118 0 131174 800
rect 132130 0 132186 800
rect 133142 0 133198 800
rect 134154 0 134210 800
rect 135166 0 135222 800
rect 136178 0 136234 800
rect 137282 0 137338 800
rect 138294 0 138350 800
rect 139306 0 139362 800
rect 140318 0 140374 800
rect 141330 0 141386 800
rect 142434 0 142490 800
rect 143446 0 143502 800
rect 144458 0 144514 800
rect 145470 0 145526 800
rect 146482 0 146538 800
rect 147494 0 147550 800
rect 148598 0 148654 800
rect 149610 0 149666 800
rect 150622 0 150678 800
rect 151634 0 151690 800
rect 152646 0 152702 800
rect 153750 0 153806 800
rect 154762 0 154818 800
rect 155774 0 155830 800
rect 156786 0 156842 800
rect 157798 0 157854 800
rect 158810 0 158866 800
rect 159914 0 159970 800
rect 160926 0 160982 800
rect 161938 0 161994 800
rect 162950 0 163006 800
rect 163962 0 164018 800
<< obsm2 >>
rect 498 165901 1158 165957
rect 1326 165901 2078 165957
rect 2246 165901 2998 165957
rect 3166 165901 3918 165957
rect 4086 165901 4838 165957
rect 5006 165901 5758 165957
rect 5926 165901 6678 165957
rect 6846 165901 7598 165957
rect 7766 165901 8518 165957
rect 8686 165901 9438 165957
rect 9606 165901 10358 165957
rect 10526 165901 11278 165957
rect 11446 165901 12198 165957
rect 12366 165901 13118 165957
rect 13286 165901 14038 165957
rect 14206 165901 14958 165957
rect 15126 165901 15878 165957
rect 16046 165901 16798 165957
rect 16966 165901 17718 165957
rect 17886 165901 18638 165957
rect 18806 165901 19558 165957
rect 19726 165901 20478 165957
rect 20646 165901 21398 165957
rect 21566 165901 22318 165957
rect 22486 165901 23238 165957
rect 23406 165901 24158 165957
rect 24326 165901 25078 165957
rect 25246 165901 25998 165957
rect 26166 165901 26918 165957
rect 27086 165901 27838 165957
rect 28006 165901 28758 165957
rect 28926 165901 29678 165957
rect 29846 165901 30598 165957
rect 30766 165901 31518 165957
rect 31686 165901 32438 165957
rect 32606 165901 33358 165957
rect 33526 165901 34278 165957
rect 34446 165901 35198 165957
rect 35366 165901 36118 165957
rect 36286 165901 37038 165957
rect 37206 165901 37958 165957
rect 38126 165901 38878 165957
rect 39046 165901 39798 165957
rect 39966 165901 40718 165957
rect 40886 165901 41638 165957
rect 41806 165901 42558 165957
rect 42726 165901 43478 165957
rect 43646 165901 44398 165957
rect 44566 165901 45318 165957
rect 45486 165901 46238 165957
rect 46406 165901 47158 165957
rect 47326 165901 48078 165957
rect 48246 165901 48998 165957
rect 49166 165901 49918 165957
rect 50086 165901 50838 165957
rect 51006 165901 51758 165957
rect 51926 165901 52678 165957
rect 52846 165901 53598 165957
rect 53766 165901 54518 165957
rect 54686 165901 55438 165957
rect 55606 165901 56358 165957
rect 56526 165901 57278 165957
rect 57446 165901 58198 165957
rect 58366 165901 59118 165957
rect 59286 165901 60038 165957
rect 60206 165901 60958 165957
rect 61126 165901 61878 165957
rect 62046 165901 62798 165957
rect 62966 165901 63718 165957
rect 63886 165901 64638 165957
rect 64806 165901 65558 165957
rect 65726 165901 66478 165957
rect 66646 165901 67398 165957
rect 67566 165901 68318 165957
rect 68486 165901 69238 165957
rect 69406 165901 70158 165957
rect 70326 165901 71078 165957
rect 71246 165901 71998 165957
rect 72166 165901 72918 165957
rect 73086 165901 73838 165957
rect 74006 165901 74758 165957
rect 74926 165901 75678 165957
rect 75846 165901 76598 165957
rect 76766 165901 77518 165957
rect 77686 165901 78438 165957
rect 78606 165901 79358 165957
rect 79526 165901 80278 165957
rect 80446 165901 81198 165957
rect 81366 165901 82118 165957
rect 82286 165901 83038 165957
rect 83206 165901 83958 165957
rect 84126 165901 84878 165957
rect 85046 165901 85798 165957
rect 85966 165901 86718 165957
rect 86886 165901 87638 165957
rect 87806 165901 88558 165957
rect 88726 165901 89478 165957
rect 89646 165901 90398 165957
rect 90566 165901 91318 165957
rect 91486 165901 92238 165957
rect 92406 165901 93158 165957
rect 93326 165901 94078 165957
rect 94246 165901 94998 165957
rect 95166 165901 95918 165957
rect 96086 165901 96838 165957
rect 97006 165901 97758 165957
rect 97926 165901 98678 165957
rect 98846 165901 99598 165957
rect 99766 165901 100518 165957
rect 100686 165901 101438 165957
rect 101606 165901 102358 165957
rect 102526 165901 103278 165957
rect 103446 165901 104198 165957
rect 104366 165901 105118 165957
rect 105286 165901 106038 165957
rect 106206 165901 106958 165957
rect 107126 165901 107878 165957
rect 108046 165901 108798 165957
rect 108966 165901 109718 165957
rect 109886 165901 110638 165957
rect 110806 165901 111558 165957
rect 111726 165901 112478 165957
rect 112646 165901 113398 165957
rect 113566 165901 114318 165957
rect 114486 165901 115238 165957
rect 115406 165901 116158 165957
rect 116326 165901 117078 165957
rect 117246 165901 117998 165957
rect 118166 165901 118918 165957
rect 119086 165901 119838 165957
rect 120006 165901 120758 165957
rect 120926 165901 121678 165957
rect 121846 165901 122598 165957
rect 122766 165901 123518 165957
rect 123686 165901 124438 165957
rect 124606 165901 125358 165957
rect 125526 165901 126278 165957
rect 126446 165901 127198 165957
rect 127366 165901 128118 165957
rect 128286 165901 129038 165957
rect 129206 165901 129958 165957
rect 130126 165901 130878 165957
rect 131046 165901 131798 165957
rect 131966 165901 132718 165957
rect 132886 165901 133638 165957
rect 133806 165901 134558 165957
rect 134726 165901 135478 165957
rect 135646 165901 136398 165957
rect 136566 165901 137318 165957
rect 137486 165901 138238 165957
rect 138406 165901 139158 165957
rect 139326 165901 140078 165957
rect 140246 165901 140998 165957
rect 141166 165901 141918 165957
rect 142086 165901 142838 165957
rect 143006 165901 143758 165957
rect 143926 165901 144678 165957
rect 144846 165901 145598 165957
rect 145766 165901 146518 165957
rect 146686 165901 147438 165957
rect 147606 165901 148358 165957
rect 148526 165901 149278 165957
rect 149446 165901 150198 165957
rect 150366 165901 151118 165957
rect 151286 165901 152038 165957
rect 152206 165901 152958 165957
rect 153126 165901 153878 165957
rect 154046 165901 154798 165957
rect 154966 165901 155718 165957
rect 155886 165901 156638 165957
rect 156806 165901 157558 165957
rect 157726 165901 158478 165957
rect 158646 165901 159398 165957
rect 159566 165901 160318 165957
rect 160486 165901 161238 165957
rect 161406 165901 162158 165957
rect 162326 165901 163078 165957
rect 163246 165901 163998 165957
rect 388 856 164016 165901
rect 388 2 422 856
rect 590 2 1434 856
rect 1602 2 2446 856
rect 2614 2 3458 856
rect 3626 2 4470 856
rect 4638 2 5482 856
rect 5650 2 6586 856
rect 6754 2 7598 856
rect 7766 2 8610 856
rect 8778 2 9622 856
rect 9790 2 10634 856
rect 10802 2 11646 856
rect 11814 2 12750 856
rect 12918 2 13762 856
rect 13930 2 14774 856
rect 14942 2 15786 856
rect 15954 2 16798 856
rect 16966 2 17902 856
rect 18070 2 18914 856
rect 19082 2 19926 856
rect 20094 2 20938 856
rect 21106 2 21950 856
rect 22118 2 22962 856
rect 23130 2 24066 856
rect 24234 2 25078 856
rect 25246 2 26090 856
rect 26258 2 27102 856
rect 27270 2 28114 856
rect 28282 2 29218 856
rect 29386 2 30230 856
rect 30398 2 31242 856
rect 31410 2 32254 856
rect 32422 2 33266 856
rect 33434 2 34278 856
rect 34446 2 35382 856
rect 35550 2 36394 856
rect 36562 2 37406 856
rect 37574 2 38418 856
rect 38586 2 39430 856
rect 39598 2 40534 856
rect 40702 2 41546 856
rect 41714 2 42558 856
rect 42726 2 43570 856
rect 43738 2 44582 856
rect 44750 2 45594 856
rect 45762 2 46698 856
rect 46866 2 47710 856
rect 47878 2 48722 856
rect 48890 2 49734 856
rect 49902 2 50746 856
rect 50914 2 51850 856
rect 52018 2 52862 856
rect 53030 2 53874 856
rect 54042 2 54886 856
rect 55054 2 55898 856
rect 56066 2 56910 856
rect 57078 2 58014 856
rect 58182 2 59026 856
rect 59194 2 60038 856
rect 60206 2 61050 856
rect 61218 2 62062 856
rect 62230 2 63166 856
rect 63334 2 64178 856
rect 64346 2 65190 856
rect 65358 2 66202 856
rect 66370 2 67214 856
rect 67382 2 68226 856
rect 68394 2 69330 856
rect 69498 2 70342 856
rect 70510 2 71354 856
rect 71522 2 72366 856
rect 72534 2 73378 856
rect 73546 2 74482 856
rect 74650 2 75494 856
rect 75662 2 76506 856
rect 76674 2 77518 856
rect 77686 2 78530 856
rect 78698 2 79542 856
rect 79710 2 80646 856
rect 80814 2 81658 856
rect 81826 2 82670 856
rect 82838 2 83682 856
rect 83850 2 84694 856
rect 84862 2 85798 856
rect 85966 2 86810 856
rect 86978 2 87822 856
rect 87990 2 88834 856
rect 89002 2 89846 856
rect 90014 2 90858 856
rect 91026 2 91962 856
rect 92130 2 92974 856
rect 93142 2 93986 856
rect 94154 2 94998 856
rect 95166 2 96010 856
rect 96178 2 97114 856
rect 97282 2 98126 856
rect 98294 2 99138 856
rect 99306 2 100150 856
rect 100318 2 101162 856
rect 101330 2 102174 856
rect 102342 2 103278 856
rect 103446 2 104290 856
rect 104458 2 105302 856
rect 105470 2 106314 856
rect 106482 2 107326 856
rect 107494 2 108430 856
rect 108598 2 109442 856
rect 109610 2 110454 856
rect 110622 2 111466 856
rect 111634 2 112478 856
rect 112646 2 113490 856
rect 113658 2 114594 856
rect 114762 2 115606 856
rect 115774 2 116618 856
rect 116786 2 117630 856
rect 117798 2 118642 856
rect 118810 2 119746 856
rect 119914 2 120758 856
rect 120926 2 121770 856
rect 121938 2 122782 856
rect 122950 2 123794 856
rect 123962 2 124806 856
rect 124974 2 125910 856
rect 126078 2 126922 856
rect 127090 2 127934 856
rect 128102 2 128946 856
rect 129114 2 129958 856
rect 130126 2 131062 856
rect 131230 2 132074 856
rect 132242 2 133086 856
rect 133254 2 134098 856
rect 134266 2 135110 856
rect 135278 2 136122 856
rect 136290 2 137226 856
rect 137394 2 138238 856
rect 138406 2 139250 856
rect 139418 2 140262 856
rect 140430 2 141274 856
rect 141442 2 142378 856
rect 142546 2 143390 856
rect 143558 2 144402 856
rect 144570 2 145414 856
rect 145582 2 146426 856
rect 146594 2 147438 856
rect 147606 2 148542 856
rect 148710 2 149554 856
rect 149722 2 150566 856
rect 150734 2 151578 856
rect 151746 2 152590 856
rect 152758 2 153694 856
rect 153862 2 154706 856
rect 154874 2 155718 856
rect 155886 2 156730 856
rect 156898 2 157742 856
rect 157910 2 158754 856
rect 158922 2 159858 856
rect 160026 2 160870 856
rect 161038 2 161882 856
rect 162050 2 162894 856
rect 163062 2 163906 856
<< metal3 >>
rect 163813 165520 164613 165640
rect 0 164976 800 165096
rect 163813 163344 164613 163464
rect 0 161576 800 161696
rect 163813 161168 164613 161288
rect 163813 158992 164613 159112
rect 0 158312 800 158432
rect 163813 156816 164613 156936
rect 0 154912 800 155032
rect 163813 154640 164613 154760
rect 163813 152464 164613 152584
rect 0 151648 800 151768
rect 163813 150152 164613 150272
rect 0 148248 800 148368
rect 163813 147976 164613 148096
rect 163813 145800 164613 145920
rect 0 144984 800 145104
rect 163813 143624 164613 143744
rect 0 141584 800 141704
rect 163813 141448 164613 141568
rect 163813 139272 164613 139392
rect 0 138320 800 138440
rect 163813 137096 164613 137216
rect 0 134920 800 135040
rect 163813 134920 164613 135040
rect 163813 132608 164613 132728
rect 0 131656 800 131776
rect 163813 130432 164613 130552
rect 0 128256 800 128376
rect 163813 128256 164613 128376
rect 163813 126080 164613 126200
rect 0 124992 800 125112
rect 163813 123904 164613 124024
rect 0 121592 800 121712
rect 163813 121728 164613 121848
rect 163813 119552 164613 119672
rect 0 118328 800 118448
rect 163813 117240 164613 117360
rect 0 114928 800 115048
rect 163813 115064 164613 115184
rect 163813 112888 164613 113008
rect 0 111664 800 111784
rect 163813 110712 164613 110832
rect 163813 108536 164613 108656
rect 0 108264 800 108384
rect 163813 106360 164613 106480
rect 0 105000 800 105120
rect 163813 104184 164613 104304
rect 163813 102008 164613 102128
rect 0 101600 800 101720
rect 163813 99696 164613 99816
rect 0 98336 800 98456
rect 163813 97520 164613 97640
rect 163813 95344 164613 95464
rect 0 94936 800 95056
rect 163813 93168 164613 93288
rect 0 91672 800 91792
rect 163813 90992 164613 91112
rect 163813 88816 164613 88936
rect 0 88272 800 88392
rect 163813 86640 164613 86760
rect 0 85008 800 85128
rect 163813 84464 164613 84584
rect 163813 82152 164613 82272
rect 0 81608 800 81728
rect 163813 79976 164613 80096
rect 0 78208 800 78328
rect 163813 77800 164613 77920
rect 163813 75624 164613 75744
rect 0 74944 800 75064
rect 163813 73448 164613 73568
rect 0 71544 800 71664
rect 163813 71272 164613 71392
rect 163813 69096 164613 69216
rect 0 68280 800 68400
rect 163813 66784 164613 66904
rect 0 64880 800 65000
rect 163813 64608 164613 64728
rect 163813 62432 164613 62552
rect 0 61616 800 61736
rect 163813 60256 164613 60376
rect 0 58216 800 58336
rect 163813 58080 164613 58200
rect 163813 55904 164613 56024
rect 0 54952 800 55072
rect 163813 53728 164613 53848
rect 0 51552 800 51672
rect 163813 51552 164613 51672
rect 163813 49240 164613 49360
rect 0 48288 800 48408
rect 163813 47064 164613 47184
rect 0 44888 800 45008
rect 163813 44888 164613 45008
rect 163813 42712 164613 42832
rect 0 41624 800 41744
rect 163813 40536 164613 40656
rect 0 38224 800 38344
rect 163813 38360 164613 38480
rect 163813 36184 164613 36304
rect 0 34960 800 35080
rect 163813 33872 164613 33992
rect 0 31560 800 31680
rect 163813 31696 164613 31816
rect 163813 29520 164613 29640
rect 0 28296 800 28416
rect 163813 27344 164613 27464
rect 163813 25168 164613 25288
rect 0 24896 800 25016
rect 163813 22992 164613 23112
rect 0 21632 800 21752
rect 163813 20816 164613 20936
rect 163813 18640 164613 18760
rect 0 18232 800 18352
rect 163813 16328 164613 16448
rect 0 14968 800 15088
rect 163813 14152 164613 14272
rect 163813 11976 164613 12096
rect 0 11568 800 11688
rect 163813 9800 164613 9920
rect 0 8304 800 8424
rect 163813 7624 164613 7744
rect 163813 5448 164613 5568
rect 0 4904 800 5024
rect 163813 3272 164613 3392
rect 0 1640 800 1760
rect 163813 1096 164613 1216
<< obsm3 >>
rect 422 163544 163813 164321
rect 422 163264 163733 163544
rect 422 161776 163813 163264
rect 880 161496 163813 161776
rect 422 161368 163813 161496
rect 422 161088 163733 161368
rect 422 159192 163813 161088
rect 422 158912 163733 159192
rect 422 158512 163813 158912
rect 880 158232 163813 158512
rect 422 157016 163813 158232
rect 422 156736 163733 157016
rect 422 155112 163813 156736
rect 880 154840 163813 155112
rect 880 154832 163733 154840
rect 422 154560 163733 154832
rect 422 152664 163813 154560
rect 422 152384 163733 152664
rect 422 151848 163813 152384
rect 880 151568 163813 151848
rect 422 150352 163813 151568
rect 422 150072 163733 150352
rect 422 148448 163813 150072
rect 880 148176 163813 148448
rect 880 148168 163733 148176
rect 422 147896 163733 148168
rect 422 146000 163813 147896
rect 422 145720 163733 146000
rect 422 145184 163813 145720
rect 880 144904 163813 145184
rect 422 143824 163813 144904
rect 422 143544 163733 143824
rect 422 141784 163813 143544
rect 880 141648 163813 141784
rect 880 141504 163733 141648
rect 422 141368 163733 141504
rect 422 139472 163813 141368
rect 422 139192 163733 139472
rect 422 138520 163813 139192
rect 880 138240 163813 138520
rect 422 137296 163813 138240
rect 422 137016 163733 137296
rect 422 135120 163813 137016
rect 880 134840 163733 135120
rect 422 132808 163813 134840
rect 422 132528 163733 132808
rect 422 131856 163813 132528
rect 880 131576 163813 131856
rect 422 130632 163813 131576
rect 422 130352 163733 130632
rect 422 128456 163813 130352
rect 880 128176 163733 128456
rect 422 126280 163813 128176
rect 422 126000 163733 126280
rect 422 125192 163813 126000
rect 880 124912 163813 125192
rect 422 124104 163813 124912
rect 422 123824 163733 124104
rect 422 121928 163813 123824
rect 422 121792 163733 121928
rect 880 121648 163733 121792
rect 880 121512 163813 121648
rect 422 119752 163813 121512
rect 422 119472 163733 119752
rect 422 118528 163813 119472
rect 880 118248 163813 118528
rect 422 117440 163813 118248
rect 422 117160 163733 117440
rect 422 115264 163813 117160
rect 422 115128 163733 115264
rect 880 114984 163733 115128
rect 880 114848 163813 114984
rect 422 113088 163813 114848
rect 422 112808 163733 113088
rect 422 111864 163813 112808
rect 880 111584 163813 111864
rect 422 110912 163813 111584
rect 422 110632 163733 110912
rect 422 108736 163813 110632
rect 422 108464 163733 108736
rect 880 108456 163733 108464
rect 880 108184 163813 108456
rect 422 106560 163813 108184
rect 422 106280 163733 106560
rect 422 105200 163813 106280
rect 880 104920 163813 105200
rect 422 104384 163813 104920
rect 422 104104 163733 104384
rect 422 102208 163813 104104
rect 422 101928 163733 102208
rect 422 101800 163813 101928
rect 880 101520 163813 101800
rect 422 99896 163813 101520
rect 422 99616 163733 99896
rect 422 98536 163813 99616
rect 880 98256 163813 98536
rect 422 97720 163813 98256
rect 422 97440 163733 97720
rect 422 95544 163813 97440
rect 422 95264 163733 95544
rect 422 95136 163813 95264
rect 880 94856 163813 95136
rect 422 93368 163813 94856
rect 422 93088 163733 93368
rect 422 91872 163813 93088
rect 880 91592 163813 91872
rect 422 91192 163813 91592
rect 422 90912 163733 91192
rect 422 89016 163813 90912
rect 422 88736 163733 89016
rect 422 88472 163813 88736
rect 880 88192 163813 88472
rect 422 86840 163813 88192
rect 422 86560 163733 86840
rect 422 85208 163813 86560
rect 880 84928 163813 85208
rect 422 84664 163813 84928
rect 422 84384 163733 84664
rect 422 82352 163813 84384
rect 422 82072 163733 82352
rect 422 81808 163813 82072
rect 880 81528 163813 81808
rect 422 80176 163813 81528
rect 422 79896 163733 80176
rect 422 78408 163813 79896
rect 880 78128 163813 78408
rect 422 78000 163813 78128
rect 422 77720 163733 78000
rect 422 75824 163813 77720
rect 422 75544 163733 75824
rect 422 75144 163813 75544
rect 880 74864 163813 75144
rect 422 73648 163813 74864
rect 422 73368 163733 73648
rect 422 71744 163813 73368
rect 880 71472 163813 71744
rect 880 71464 163733 71472
rect 422 71192 163733 71464
rect 422 69296 163813 71192
rect 422 69016 163733 69296
rect 422 68480 163813 69016
rect 880 68200 163813 68480
rect 422 66984 163813 68200
rect 422 66704 163733 66984
rect 422 65080 163813 66704
rect 880 64808 163813 65080
rect 880 64800 163733 64808
rect 422 64528 163733 64800
rect 422 62632 163813 64528
rect 422 62352 163733 62632
rect 422 61816 163813 62352
rect 880 61536 163813 61816
rect 422 60456 163813 61536
rect 422 60176 163733 60456
rect 422 58416 163813 60176
rect 880 58280 163813 58416
rect 880 58136 163733 58280
rect 422 58000 163733 58136
rect 422 56104 163813 58000
rect 422 55824 163733 56104
rect 422 55152 163813 55824
rect 880 54872 163813 55152
rect 422 53928 163813 54872
rect 422 53648 163733 53928
rect 422 51752 163813 53648
rect 880 51472 163733 51752
rect 422 49440 163813 51472
rect 422 49160 163733 49440
rect 422 48488 163813 49160
rect 880 48208 163813 48488
rect 422 47264 163813 48208
rect 422 46984 163733 47264
rect 422 45088 163813 46984
rect 880 44808 163733 45088
rect 422 42912 163813 44808
rect 422 42632 163733 42912
rect 422 41824 163813 42632
rect 880 41544 163813 41824
rect 422 40736 163813 41544
rect 422 40456 163733 40736
rect 422 38560 163813 40456
rect 422 38424 163733 38560
rect 880 38280 163733 38424
rect 880 38144 163813 38280
rect 422 36384 163813 38144
rect 422 36104 163733 36384
rect 422 35160 163813 36104
rect 880 34880 163813 35160
rect 422 34072 163813 34880
rect 422 33792 163733 34072
rect 422 31896 163813 33792
rect 422 31760 163733 31896
rect 880 31616 163733 31760
rect 880 31480 163813 31616
rect 422 29720 163813 31480
rect 422 29440 163733 29720
rect 422 28496 163813 29440
rect 880 28216 163813 28496
rect 422 27544 163813 28216
rect 422 27264 163733 27544
rect 422 25368 163813 27264
rect 422 25096 163733 25368
rect 880 25088 163733 25096
rect 880 24816 163813 25088
rect 422 23192 163813 24816
rect 422 22912 163733 23192
rect 422 21832 163813 22912
rect 880 21552 163813 21832
rect 422 21016 163813 21552
rect 422 20736 163733 21016
rect 422 18840 163813 20736
rect 422 18560 163733 18840
rect 422 18432 163813 18560
rect 880 18152 163813 18432
rect 422 16528 163813 18152
rect 422 16248 163733 16528
rect 422 15168 163813 16248
rect 880 14888 163813 15168
rect 422 14352 163813 14888
rect 422 14072 163733 14352
rect 422 12176 163813 14072
rect 422 11896 163733 12176
rect 422 11768 163813 11896
rect 880 11488 163813 11768
rect 422 10000 163813 11488
rect 422 9720 163733 10000
rect 422 8504 163813 9720
rect 880 8224 163813 8504
rect 422 7824 163813 8224
rect 422 7544 163733 7824
rect 422 5648 163813 7544
rect 422 5368 163733 5648
rect 422 5104 163813 5368
rect 880 4824 163813 5104
rect 422 3472 163813 4824
rect 422 3192 163733 3472
rect 422 1840 163813 3192
rect 880 1560 163813 1840
rect 422 1296 163813 1560
rect 422 1016 163733 1296
rect 422 35 163813 1016
<< metal4 >>
rect 4208 2128 4528 164336
rect 19568 2128 19888 164336
rect 34928 2128 35248 164336
rect 50288 2128 50608 164336
rect 65648 2128 65968 164336
rect 81008 2128 81328 164336
rect 96368 2128 96688 164336
rect 111728 2128 112048 164336
rect 127088 2128 127408 164336
rect 142448 2128 142768 164336
rect 157808 2128 158128 164336
<< obsm4 >>
rect 427 2048 4128 164117
rect 4608 2048 19488 164117
rect 19968 2048 34848 164117
rect 35328 2048 50208 164117
rect 50688 2048 65568 164117
rect 66048 2048 80928 164117
rect 81408 2048 96288 164117
rect 96768 2048 111648 164117
rect 112128 2048 127008 164117
rect 127488 2048 142368 164117
rect 142848 2048 148242 164117
rect 427 35 148242 2048
<< labels >>
rlabel metal2 s 107014 165957 107070 166757 6 i_dout0[0]
port 1 nsew signal input
rlabel metal2 s 130934 165957 130990 166757 6 i_dout0[10]
port 2 nsew signal input
rlabel metal2 s 141330 0 141386 800 6 i_dout0[11]
port 3 nsew signal input
rlabel metal2 s 138294 165957 138350 166757 6 i_dout0[12]
port 4 nsew signal input
rlabel metal3 s 0 78208 800 78328 6 i_dout0[13]
port 5 nsew signal input
rlabel metal3 s 0 88272 800 88392 6 i_dout0[14]
port 6 nsew signal input
rlabel metal2 s 145470 0 145526 800 6 i_dout0[15]
port 7 nsew signal input
rlabel metal3 s 0 94936 800 95056 6 i_dout0[16]
port 8 nsew signal input
rlabel metal2 s 149610 0 149666 800 6 i_dout0[17]
port 9 nsew signal input
rlabel metal2 s 144734 165957 144790 166757 6 i_dout0[18]
port 10 nsew signal input
rlabel metal3 s 163813 117240 164613 117360 6 i_dout0[19]
port 11 nsew signal input
rlabel metal3 s 163813 11976 164613 12096 6 i_dout0[1]
port 12 nsew signal input
rlabel metal3 s 0 108264 800 108384 6 i_dout0[20]
port 13 nsew signal input
rlabel metal3 s 163813 128256 164613 128376 6 i_dout0[21]
port 14 nsew signal input
rlabel metal3 s 163813 132608 164613 132728 6 i_dout0[22]
port 15 nsew signal input
rlabel metal3 s 0 124992 800 125112 6 i_dout0[23]
port 16 nsew signal input
rlabel metal2 s 152094 165957 152150 166757 6 i_dout0[24]
port 17 nsew signal input
rlabel metal3 s 0 141584 800 141704 6 i_dout0[25]
port 18 nsew signal input
rlabel metal3 s 0 151648 800 151768 6 i_dout0[26]
port 19 nsew signal input
rlabel metal2 s 155774 165957 155830 166757 6 i_dout0[27]
port 20 nsew signal input
rlabel metal2 s 158534 165957 158590 166757 6 i_dout0[28]
port 21 nsew signal input
rlabel metal3 s 163813 154640 164613 154760 6 i_dout0[29]
port 22 nsew signal input
rlabel metal3 s 163813 25168 164613 25288 6 i_dout0[2]
port 23 nsew signal input
rlabel metal2 s 161294 165957 161350 166757 6 i_dout0[30]
port 24 nsew signal input
rlabel metal2 s 164054 165957 164110 166757 6 i_dout0[31]
port 25 nsew signal input
rlabel metal2 s 113454 165957 113510 166757 6 i_dout0[3]
port 26 nsew signal input
rlabel metal2 s 118054 165957 118110 166757 6 i_dout0[4]
port 27 nsew signal input
rlabel metal3 s 0 44888 800 45008 6 i_dout0[5]
port 28 nsew signal input
rlabel metal3 s 0 48288 800 48408 6 i_dout0[6]
port 29 nsew signal input
rlabel metal3 s 163813 64608 164613 64728 6 i_dout0[7]
port 30 nsew signal input
rlabel metal2 s 126334 165957 126390 166757 6 i_dout0[8]
port 31 nsew signal input
rlabel metal2 s 139306 0 139362 800 6 i_dout0[9]
port 32 nsew signal input
rlabel metal2 s 113546 0 113602 800 6 i_dout0_1[0]
port 33 nsew signal input
rlabel metal3 s 163813 75624 164613 75744 6 i_dout0_1[10]
port 34 nsew signal input
rlabel metal2 s 134614 165957 134670 166757 6 i_dout0_1[11]
port 35 nsew signal input
rlabel metal2 s 137374 165957 137430 166757 6 i_dout0_1[12]
port 36 nsew signal input
rlabel metal3 s 0 71544 800 71664 6 i_dout0_1[13]
port 37 nsew signal input
rlabel metal3 s 0 85008 800 85128 6 i_dout0_1[14]
port 38 nsew signal input
rlabel metal2 s 144458 0 144514 800 6 i_dout0_1[15]
port 39 nsew signal input
rlabel metal2 s 146482 0 146538 800 6 i_dout0_1[16]
port 40 nsew signal input
rlabel metal2 s 148598 0 148654 800 6 i_dout0_1[17]
port 41 nsew signal input
rlabel metal3 s 163813 106360 164613 106480 6 i_dout0_1[18]
port 42 nsew signal input
rlabel metal3 s 163813 115064 164613 115184 6 i_dout0_1[19]
port 43 nsew signal input
rlabel metal2 s 119802 0 119858 800 6 i_dout0_1[1]
port 44 nsew signal input
rlabel metal3 s 163813 119552 164613 119672 6 i_dout0_1[20]
port 45 nsew signal input
rlabel metal3 s 163813 123904 164613 124024 6 i_dout0_1[21]
port 46 nsew signal input
rlabel metal2 s 149334 165957 149390 166757 6 i_dout0_1[22]
port 47 nsew signal input
rlabel metal2 s 154762 0 154818 800 6 i_dout0_1[23]
port 48 nsew signal input
rlabel metal3 s 163813 139272 164613 139392 6 i_dout0_1[24]
port 49 nsew signal input
rlabel metal2 s 153014 165957 153070 166757 6 i_dout0_1[25]
port 50 nsew signal input
rlabel metal2 s 153934 165957 153990 166757 6 i_dout0_1[26]
port 51 nsew signal input
rlabel metal3 s 163813 145800 164613 145920 6 i_dout0_1[27]
port 52 nsew signal input
rlabel metal3 s 163813 147976 164613 148096 6 i_dout0_1[28]
port 53 nsew signal input
rlabel metal3 s 163813 150152 164613 150272 6 i_dout0_1[29]
port 54 nsew signal input
rlabel metal3 s 0 14968 800 15088 6 i_dout0_1[2]
port 55 nsew signal input
rlabel metal3 s 0 158312 800 158432 6 i_dout0_1[30]
port 56 nsew signal input
rlabel metal2 s 163134 165957 163190 166757 6 i_dout0_1[31]
port 57 nsew signal input
rlabel metal2 s 112534 165957 112590 166757 6 i_dout0_1[3]
port 58 nsew signal input
rlabel metal2 s 116214 165957 116270 166757 6 i_dout0_1[4]
port 59 nsew signal input
rlabel metal3 s 163813 47064 164613 47184 6 i_dout0_1[5]
port 60 nsew signal input
rlabel metal3 s 163813 58080 164613 58200 6 i_dout0_1[6]
port 61 nsew signal input
rlabel metal3 s 0 54952 800 55072 6 i_dout0_1[7]
port 62 nsew signal input
rlabel metal2 s 135166 0 135222 800 6 i_dout0_1[8]
port 63 nsew signal input
rlabel metal2 s 138294 0 138350 800 6 i_dout0_1[9]
port 64 nsew signal input
rlabel metal3 s 163813 7624 164613 7744 6 i_dout1[0]
port 65 nsew signal input
rlabel metal2 s 131854 165957 131910 166757 6 i_dout1[10]
port 66 nsew signal input
rlabel metal3 s 163813 79976 164613 80096 6 i_dout1[11]
port 67 nsew signal input
rlabel metal2 s 139214 165957 139270 166757 6 i_dout1[12]
port 68 nsew signal input
rlabel metal2 s 141054 165957 141110 166757 6 i_dout1[13]
port 69 nsew signal input
rlabel metal2 s 143446 0 143502 800 6 i_dout1[14]
port 70 nsew signal input
rlabel metal3 s 163813 95344 164613 95464 6 i_dout1[15]
port 71 nsew signal input
rlabel metal3 s 163813 99696 164613 99816 6 i_dout1[16]
port 72 nsew signal input
rlabel metal3 s 163813 104184 164613 104304 6 i_dout1[17]
port 73 nsew signal input
rlabel metal2 s 151634 0 151690 800 6 i_dout1[18]
port 74 nsew signal input
rlabel metal3 s 0 98336 800 98456 6 i_dout1[19]
port 75 nsew signal input
rlabel metal2 s 108854 165957 108910 166757 6 i_dout1[1]
port 76 nsew signal input
rlabel metal2 s 147494 165957 147550 166757 6 i_dout1[20]
port 77 nsew signal input
rlabel metal3 s 163813 130432 164613 130552 6 i_dout1[21]
port 78 nsew signal input
rlabel metal2 s 153750 0 153806 800 6 i_dout1[22]
port 79 nsew signal input
rlabel metal2 s 150254 165957 150310 166757 6 i_dout1[23]
port 80 nsew signal input
rlabel metal3 s 0 131656 800 131776 6 i_dout1[24]
port 81 nsew signal input
rlabel metal3 s 163813 141448 164613 141568 6 i_dout1[25]
port 82 nsew signal input
rlabel metal3 s 0 154912 800 155032 6 i_dout1[26]
port 83 nsew signal input
rlabel metal2 s 156694 165957 156750 166757 6 i_dout1[27]
port 84 nsew signal input
rlabel metal2 s 159454 165957 159510 166757 6 i_dout1[28]
port 85 nsew signal input
rlabel metal3 s 163813 156816 164613 156936 6 i_dout1[29]
port 86 nsew signal input
rlabel metal3 s 0 21632 800 21752 6 i_dout1[2]
port 87 nsew signal input
rlabel metal3 s 0 161576 800 161696 6 i_dout1[30]
port 88 nsew signal input
rlabel metal3 s 0 164976 800 165096 6 i_dout1[31]
port 89 nsew signal input
rlabel metal3 s 0 34960 800 35080 6 i_dout1[3]
port 90 nsew signal input
rlabel metal2 s 123850 0 123906 800 6 i_dout1[4]
port 91 nsew signal input
rlabel metal2 s 126978 0 127034 800 6 i_dout1[5]
port 92 nsew signal input
rlabel metal2 s 130014 0 130070 800 6 i_dout1[6]
port 93 nsew signal input
rlabel metal2 s 131118 0 131174 800 6 i_dout1[7]
port 94 nsew signal input
rlabel metal2 s 127254 165957 127310 166757 6 i_dout1[8]
port 95 nsew signal input
rlabel metal2 s 140318 0 140374 800 6 i_dout1[9]
port 96 nsew signal input
rlabel metal3 s 163813 5448 164613 5568 6 i_dout1_1[0]
port 97 nsew signal input
rlabel metal3 s 0 68280 800 68400 6 i_dout1_1[10]
port 98 nsew signal input
rlabel metal3 s 163813 77800 164613 77920 6 i_dout1_1[11]
port 99 nsew signal input
rlabel metal2 s 142434 0 142490 800 6 i_dout1_1[12]
port 100 nsew signal input
rlabel metal3 s 0 74944 800 75064 6 i_dout1_1[13]
port 101 nsew signal input
rlabel metal3 s 163813 86640 164613 86760 6 i_dout1_1[14]
port 102 nsew signal input
rlabel metal3 s 163813 93168 164613 93288 6 i_dout1_1[15]
port 103 nsew signal input
rlabel metal2 s 141974 165957 142030 166757 6 i_dout1_1[16]
port 104 nsew signal input
rlabel metal3 s 163813 102008 164613 102128 6 i_dout1_1[17]
port 105 nsew signal input
rlabel metal3 s 163813 108536 164613 108656 6 i_dout1_1[18]
port 106 nsew signal input
rlabel metal2 s 145654 165957 145710 166757 6 i_dout1_1[19]
port 107 nsew signal input
rlabel metal3 s 0 8304 800 8424 6 i_dout1_1[1]
port 108 nsew signal input
rlabel metal3 s 0 105000 800 105120 6 i_dout1_1[20]
port 109 nsew signal input
rlabel metal3 s 163813 126080 164613 126200 6 i_dout1_1[21]
port 110 nsew signal input
rlabel metal3 s 0 114928 800 115048 6 i_dout1_1[22]
port 111 nsew signal input
rlabel metal3 s 0 121592 800 121712 6 i_dout1_1[23]
port 112 nsew signal input
rlabel metal2 s 151174 165957 151230 166757 6 i_dout1_1[24]
port 113 nsew signal input
rlabel metal3 s 0 138320 800 138440 6 i_dout1_1[25]
port 114 nsew signal input
rlabel metal3 s 0 148248 800 148368 6 i_dout1_1[26]
port 115 nsew signal input
rlabel metal2 s 157798 0 157854 800 6 i_dout1_1[27]
port 116 nsew signal input
rlabel metal2 s 159914 0 159970 800 6 i_dout1_1[28]
port 117 nsew signal input
rlabel metal3 s 163813 152464 164613 152584 6 i_dout1_1[29]
port 118 nsew signal input
rlabel metal3 s 0 18232 800 18352 6 i_dout1_1[2]
port 119 nsew signal input
rlabel metal3 s 163813 161168 164613 161288 6 i_dout1_1[30]
port 120 nsew signal input
rlabel metal3 s 163813 165520 164613 165640 6 i_dout1_1[31]
port 121 nsew signal input
rlabel metal3 s 163813 33872 164613 33992 6 i_dout1_1[3]
port 122 nsew signal input
rlabel metal2 s 117134 165957 117190 166757 6 i_dout1_1[4]
port 123 nsew signal input
rlabel metal2 s 119894 165957 119950 166757 6 i_dout1_1[5]
port 124 nsew signal input
rlabel metal3 s 163813 60256 164613 60376 6 i_dout1_1[6]
port 125 nsew signal input
rlabel metal2 s 124494 165957 124550 166757 6 i_dout1_1[7]
port 126 nsew signal input
rlabel metal2 s 136178 0 136234 800 6 i_dout1_1[8]
port 127 nsew signal input
rlabel metal3 s 163813 71272 164613 71392 6 i_dout1_1[9]
port 128 nsew signal input
rlabel metal2 s 386 165957 442 166757 6 io_in[0]
port 129 nsew signal input
rlabel metal2 s 27894 165957 27950 166757 6 io_in[10]
port 130 nsew signal input
rlabel metal2 s 30654 165957 30710 166757 6 io_in[11]
port 131 nsew signal input
rlabel metal2 s 33414 165957 33470 166757 6 io_in[12]
port 132 nsew signal input
rlabel metal2 s 36174 165957 36230 166757 6 io_in[13]
port 133 nsew signal input
rlabel metal2 s 38934 165957 38990 166757 6 io_in[14]
port 134 nsew signal input
rlabel metal2 s 41694 165957 41750 166757 6 io_in[15]
port 135 nsew signal input
rlabel metal2 s 44454 165957 44510 166757 6 io_in[16]
port 136 nsew signal input
rlabel metal2 s 47214 165957 47270 166757 6 io_in[17]
port 137 nsew signal input
rlabel metal2 s 49974 165957 50030 166757 6 io_in[18]
port 138 nsew signal input
rlabel metal2 s 52734 165957 52790 166757 6 io_in[19]
port 139 nsew signal input
rlabel metal2 s 3054 165957 3110 166757 6 io_in[1]
port 140 nsew signal input
rlabel metal2 s 55494 165957 55550 166757 6 io_in[20]
port 141 nsew signal input
rlabel metal2 s 58254 165957 58310 166757 6 io_in[21]
port 142 nsew signal input
rlabel metal2 s 61014 165957 61070 166757 6 io_in[22]
port 143 nsew signal input
rlabel metal2 s 63774 165957 63830 166757 6 io_in[23]
port 144 nsew signal input
rlabel metal2 s 66534 165957 66590 166757 6 io_in[24]
port 145 nsew signal input
rlabel metal2 s 69294 165957 69350 166757 6 io_in[25]
port 146 nsew signal input
rlabel metal2 s 72054 165957 72110 166757 6 io_in[26]
port 147 nsew signal input
rlabel metal2 s 74814 165957 74870 166757 6 io_in[27]
port 148 nsew signal input
rlabel metal2 s 77574 165957 77630 166757 6 io_in[28]
port 149 nsew signal input
rlabel metal2 s 80334 165957 80390 166757 6 io_in[29]
port 150 nsew signal input
rlabel metal2 s 5814 165957 5870 166757 6 io_in[2]
port 151 nsew signal input
rlabel metal2 s 83094 165957 83150 166757 6 io_in[30]
port 152 nsew signal input
rlabel metal2 s 85854 165957 85910 166757 6 io_in[31]
port 153 nsew signal input
rlabel metal2 s 88614 165957 88670 166757 6 io_in[32]
port 154 nsew signal input
rlabel metal2 s 91374 165957 91430 166757 6 io_in[33]
port 155 nsew signal input
rlabel metal2 s 94134 165957 94190 166757 6 io_in[34]
port 156 nsew signal input
rlabel metal2 s 96894 165957 96950 166757 6 io_in[35]
port 157 nsew signal input
rlabel metal2 s 99654 165957 99710 166757 6 io_in[36]
port 158 nsew signal input
rlabel metal2 s 102414 165957 102470 166757 6 io_in[37]
port 159 nsew signal input
rlabel metal2 s 8574 165957 8630 166757 6 io_in[3]
port 160 nsew signal input
rlabel metal2 s 11334 165957 11390 166757 6 io_in[4]
port 161 nsew signal input
rlabel metal2 s 14094 165957 14150 166757 6 io_in[5]
port 162 nsew signal input
rlabel metal2 s 16854 165957 16910 166757 6 io_in[6]
port 163 nsew signal input
rlabel metal2 s 19614 165957 19670 166757 6 io_in[7]
port 164 nsew signal input
rlabel metal2 s 22374 165957 22430 166757 6 io_in[8]
port 165 nsew signal input
rlabel metal2 s 25134 165957 25190 166757 6 io_in[9]
port 166 nsew signal input
rlabel metal2 s 1214 165957 1270 166757 6 io_oeb[0]
port 167 nsew signal output
rlabel metal2 s 28814 165957 28870 166757 6 io_oeb[10]
port 168 nsew signal output
rlabel metal2 s 31574 165957 31630 166757 6 io_oeb[11]
port 169 nsew signal output
rlabel metal2 s 34334 165957 34390 166757 6 io_oeb[12]
port 170 nsew signal output
rlabel metal2 s 37094 165957 37150 166757 6 io_oeb[13]
port 171 nsew signal output
rlabel metal2 s 39854 165957 39910 166757 6 io_oeb[14]
port 172 nsew signal output
rlabel metal2 s 42614 165957 42670 166757 6 io_oeb[15]
port 173 nsew signal output
rlabel metal2 s 45374 165957 45430 166757 6 io_oeb[16]
port 174 nsew signal output
rlabel metal2 s 48134 165957 48190 166757 6 io_oeb[17]
port 175 nsew signal output
rlabel metal2 s 50894 165957 50950 166757 6 io_oeb[18]
port 176 nsew signal output
rlabel metal2 s 53654 165957 53710 166757 6 io_oeb[19]
port 177 nsew signal output
rlabel metal2 s 3974 165957 4030 166757 6 io_oeb[1]
port 178 nsew signal output
rlabel metal2 s 56414 165957 56470 166757 6 io_oeb[20]
port 179 nsew signal output
rlabel metal2 s 59174 165957 59230 166757 6 io_oeb[21]
port 180 nsew signal output
rlabel metal2 s 61934 165957 61990 166757 6 io_oeb[22]
port 181 nsew signal output
rlabel metal2 s 64694 165957 64750 166757 6 io_oeb[23]
port 182 nsew signal output
rlabel metal2 s 67454 165957 67510 166757 6 io_oeb[24]
port 183 nsew signal output
rlabel metal2 s 70214 165957 70270 166757 6 io_oeb[25]
port 184 nsew signal output
rlabel metal2 s 72974 165957 73030 166757 6 io_oeb[26]
port 185 nsew signal output
rlabel metal2 s 75734 165957 75790 166757 6 io_oeb[27]
port 186 nsew signal output
rlabel metal2 s 78494 165957 78550 166757 6 io_oeb[28]
port 187 nsew signal output
rlabel metal2 s 81254 165957 81310 166757 6 io_oeb[29]
port 188 nsew signal output
rlabel metal2 s 6734 165957 6790 166757 6 io_oeb[2]
port 189 nsew signal output
rlabel metal2 s 84014 165957 84070 166757 6 io_oeb[30]
port 190 nsew signal output
rlabel metal2 s 86774 165957 86830 166757 6 io_oeb[31]
port 191 nsew signal output
rlabel metal2 s 89534 165957 89590 166757 6 io_oeb[32]
port 192 nsew signal output
rlabel metal2 s 92294 165957 92350 166757 6 io_oeb[33]
port 193 nsew signal output
rlabel metal2 s 95054 165957 95110 166757 6 io_oeb[34]
port 194 nsew signal output
rlabel metal2 s 97814 165957 97870 166757 6 io_oeb[35]
port 195 nsew signal output
rlabel metal2 s 100574 165957 100630 166757 6 io_oeb[36]
port 196 nsew signal output
rlabel metal2 s 103334 165957 103390 166757 6 io_oeb[37]
port 197 nsew signal output
rlabel metal2 s 9494 165957 9550 166757 6 io_oeb[3]
port 198 nsew signal output
rlabel metal2 s 12254 165957 12310 166757 6 io_oeb[4]
port 199 nsew signal output
rlabel metal2 s 15014 165957 15070 166757 6 io_oeb[5]
port 200 nsew signal output
rlabel metal2 s 17774 165957 17830 166757 6 io_oeb[6]
port 201 nsew signal output
rlabel metal2 s 20534 165957 20590 166757 6 io_oeb[7]
port 202 nsew signal output
rlabel metal2 s 23294 165957 23350 166757 6 io_oeb[8]
port 203 nsew signal output
rlabel metal2 s 26054 165957 26110 166757 6 io_oeb[9]
port 204 nsew signal output
rlabel metal2 s 2134 165957 2190 166757 6 io_out[0]
port 205 nsew signal output
rlabel metal2 s 29734 165957 29790 166757 6 io_out[10]
port 206 nsew signal output
rlabel metal2 s 32494 165957 32550 166757 6 io_out[11]
port 207 nsew signal output
rlabel metal2 s 35254 165957 35310 166757 6 io_out[12]
port 208 nsew signal output
rlabel metal2 s 38014 165957 38070 166757 6 io_out[13]
port 209 nsew signal output
rlabel metal2 s 40774 165957 40830 166757 6 io_out[14]
port 210 nsew signal output
rlabel metal2 s 43534 165957 43590 166757 6 io_out[15]
port 211 nsew signal output
rlabel metal2 s 46294 165957 46350 166757 6 io_out[16]
port 212 nsew signal output
rlabel metal2 s 49054 165957 49110 166757 6 io_out[17]
port 213 nsew signal output
rlabel metal2 s 51814 165957 51870 166757 6 io_out[18]
port 214 nsew signal output
rlabel metal2 s 54574 165957 54630 166757 6 io_out[19]
port 215 nsew signal output
rlabel metal2 s 4894 165957 4950 166757 6 io_out[1]
port 216 nsew signal output
rlabel metal2 s 57334 165957 57390 166757 6 io_out[20]
port 217 nsew signal output
rlabel metal2 s 60094 165957 60150 166757 6 io_out[21]
port 218 nsew signal output
rlabel metal2 s 62854 165957 62910 166757 6 io_out[22]
port 219 nsew signal output
rlabel metal2 s 65614 165957 65670 166757 6 io_out[23]
port 220 nsew signal output
rlabel metal2 s 68374 165957 68430 166757 6 io_out[24]
port 221 nsew signal output
rlabel metal2 s 71134 165957 71190 166757 6 io_out[25]
port 222 nsew signal output
rlabel metal2 s 73894 165957 73950 166757 6 io_out[26]
port 223 nsew signal output
rlabel metal2 s 76654 165957 76710 166757 6 io_out[27]
port 224 nsew signal output
rlabel metal2 s 79414 165957 79470 166757 6 io_out[28]
port 225 nsew signal output
rlabel metal2 s 82174 165957 82230 166757 6 io_out[29]
port 226 nsew signal output
rlabel metal2 s 7654 165957 7710 166757 6 io_out[2]
port 227 nsew signal output
rlabel metal2 s 84934 165957 84990 166757 6 io_out[30]
port 228 nsew signal output
rlabel metal2 s 87694 165957 87750 166757 6 io_out[31]
port 229 nsew signal output
rlabel metal2 s 90454 165957 90510 166757 6 io_out[32]
port 230 nsew signal output
rlabel metal2 s 93214 165957 93270 166757 6 io_out[33]
port 231 nsew signal output
rlabel metal2 s 95974 165957 96030 166757 6 io_out[34]
port 232 nsew signal output
rlabel metal2 s 98734 165957 98790 166757 6 io_out[35]
port 233 nsew signal output
rlabel metal2 s 101494 165957 101550 166757 6 io_out[36]
port 234 nsew signal output
rlabel metal2 s 104254 165957 104310 166757 6 io_out[37]
port 235 nsew signal output
rlabel metal2 s 10414 165957 10470 166757 6 io_out[3]
port 236 nsew signal output
rlabel metal2 s 13174 165957 13230 166757 6 io_out[4]
port 237 nsew signal output
rlabel metal2 s 15934 165957 15990 166757 6 io_out[5]
port 238 nsew signal output
rlabel metal2 s 18694 165957 18750 166757 6 io_out[6]
port 239 nsew signal output
rlabel metal2 s 21454 165957 21510 166757 6 io_out[7]
port 240 nsew signal output
rlabel metal2 s 24214 165957 24270 166757 6 io_out[8]
port 241 nsew signal output
rlabel metal2 s 26974 165957 27030 166757 6 io_out[9]
port 242 nsew signal output
rlabel metal2 s 109498 0 109554 800 6 irq[0]
port 243 nsew signal output
rlabel metal2 s 110510 0 110566 800 6 irq[1]
port 244 nsew signal output
rlabel metal2 s 111522 0 111578 800 6 irq[2]
port 245 nsew signal output
rlabel metal2 s 115662 0 115718 800 6 o_addr1[0]
port 246 nsew signal output
rlabel metal2 s 109774 165957 109830 166757 6 o_addr1[1]
port 247 nsew signal output
rlabel metal3 s 163813 29520 164613 29640 6 o_addr1[2]
port 248 nsew signal output
rlabel metal3 s 0 38224 800 38344 6 o_addr1[3]
port 249 nsew signal output
rlabel metal2 s 124862 0 124918 800 6 o_addr1[4]
port 250 nsew signal output
rlabel metal2 s 127990 0 128046 800 6 o_addr1[5]
port 251 nsew signal output
rlabel metal3 s 0 51552 800 51672 6 o_addr1[6]
port 252 nsew signal output
rlabel metal3 s 163813 66784 164613 66904 6 o_addr1[7]
port 253 nsew signal output
rlabel metal3 s 0 61616 800 61736 6 o_addr1[8]
port 254 nsew signal output
rlabel metal2 s 114650 0 114706 800 6 o_addr1_1[0]
port 255 nsew signal output
rlabel metal3 s 163813 14152 164613 14272 6 o_addr1_1[1]
port 256 nsew signal output
rlabel metal3 s 163813 27344 164613 27464 6 o_addr1_1[2]
port 257 nsew signal output
rlabel metal2 s 114374 165957 114430 166757 6 o_addr1_1[3]
port 258 nsew signal output
rlabel metal3 s 163813 42712 164613 42832 6 o_addr1_1[4]
port 259 nsew signal output
rlabel metal3 s 163813 49240 164613 49360 6 o_addr1_1[5]
port 260 nsew signal output
rlabel metal2 s 120814 165957 120870 166757 6 o_addr1_1[6]
port 261 nsew signal output
rlabel metal2 s 125414 165957 125470 166757 6 o_addr1_1[7]
port 262 nsew signal output
rlabel metal2 s 128174 165957 128230 166757 6 o_addr1_1[8]
port 263 nsew signal output
rlabel metal2 s 105174 165957 105230 166757 6 o_csb0
port 264 nsew signal output
rlabel metal3 s 163813 1096 164613 1216 6 o_csb0_1
port 265 nsew signal output
rlabel metal3 s 163813 3272 164613 3392 6 o_csb1
port 266 nsew signal output
rlabel metal2 s 106094 165957 106150 166757 6 o_csb1_1
port 267 nsew signal output
rlabel metal2 s 116674 0 116730 800 6 o_din0[0]
port 268 nsew signal output
rlabel metal2 s 133694 165957 133750 166757 6 o_din0[10]
port 269 nsew signal output
rlabel metal2 s 136454 165957 136510 166757 6 o_din0[11]
port 270 nsew signal output
rlabel metal3 s 163813 82152 164613 82272 6 o_din0[12]
port 271 nsew signal output
rlabel metal3 s 163813 84464 164613 84584 6 o_din0[13]
port 272 nsew signal output
rlabel metal3 s 163813 90992 164613 91112 6 o_din0[14]
port 273 nsew signal output
rlabel metal3 s 163813 97520 164613 97640 6 o_din0[15]
port 274 nsew signal output
rlabel metal2 s 147494 0 147550 800 6 o_din0[16]
port 275 nsew signal output
rlabel metal2 s 143814 165957 143870 166757 6 o_din0[17]
port 276 nsew signal output
rlabel metal3 s 163813 112888 164613 113008 6 o_din0[18]
port 277 nsew signal output
rlabel metal3 s 0 101600 800 101720 6 o_din0[19]
port 278 nsew signal output
rlabel metal2 s 110694 165957 110750 166757 6 o_din0[1]
port 279 nsew signal output
rlabel metal3 s 0 111664 800 111784 6 o_din0[20]
port 280 nsew signal output
rlabel metal2 s 148414 165957 148470 166757 6 o_din0[21]
port 281 nsew signal output
rlabel metal3 s 163813 134920 164613 135040 6 o_din0[22]
port 282 nsew signal output
rlabel metal3 s 0 128256 800 128376 6 o_din0[23]
port 283 nsew signal output
rlabel metal3 s 0 134920 800 135040 6 o_din0[24]
port 284 nsew signal output
rlabel metal3 s 163813 143624 164613 143744 6 o_din0[25]
port 285 nsew signal output
rlabel metal2 s 154854 165957 154910 166757 6 o_din0[26]
port 286 nsew signal output
rlabel metal2 s 158810 0 158866 800 6 o_din0[27]
port 287 nsew signal output
rlabel metal2 s 160926 0 160982 800 6 o_din0[28]
port 288 nsew signal output
rlabel metal3 s 163813 158992 164613 159112 6 o_din0[29]
port 289 nsew signal output
rlabel metal2 s 120814 0 120870 800 6 o_din0[2]
port 290 nsew signal output
rlabel metal2 s 162214 165957 162270 166757 6 o_din0[30]
port 291 nsew signal output
rlabel metal2 s 163962 0 164018 800 6 o_din0[31]
port 292 nsew signal output
rlabel metal2 s 121826 0 121882 800 6 o_din0[3]
port 293 nsew signal output
rlabel metal3 s 163813 44888 164613 45008 6 o_din0[4]
port 294 nsew signal output
rlabel metal3 s 163813 53728 164613 53848 6 o_din0[5]
port 295 nsew signal output
rlabel metal2 s 121734 165957 121790 166757 6 o_din0[6]
port 296 nsew signal output
rlabel metal2 s 133142 0 133198 800 6 o_din0[7]
port 297 nsew signal output
rlabel metal2 s 129094 165957 129150 166757 6 o_din0[8]
port 298 nsew signal output
rlabel metal3 s 0 64880 800 65000 6 o_din0[9]
port 299 nsew signal output
rlabel metal2 s 117686 0 117742 800 6 o_din0_1[0]
port 300 nsew signal output
rlabel metal2 s 132774 165957 132830 166757 6 o_din0_1[10]
port 301 nsew signal output
rlabel metal2 s 135534 165957 135590 166757 6 o_din0_1[11]
port 302 nsew signal output
rlabel metal2 s 140134 165957 140190 166757 6 o_din0_1[12]
port 303 nsew signal output
rlabel metal3 s 0 81608 800 81728 6 o_din0_1[13]
port 304 nsew signal output
rlabel metal3 s 163813 88816 164613 88936 6 o_din0_1[14]
port 305 nsew signal output
rlabel metal3 s 0 91672 800 91792 6 o_din0_1[15]
port 306 nsew signal output
rlabel metal2 s 142894 165957 142950 166757 6 o_din0_1[16]
port 307 nsew signal output
rlabel metal2 s 150622 0 150678 800 6 o_din0_1[17]
port 308 nsew signal output
rlabel metal3 s 163813 110712 164613 110832 6 o_din0_1[18]
port 309 nsew signal output
rlabel metal2 s 146574 165957 146630 166757 6 o_din0_1[19]
port 310 nsew signal output
rlabel metal3 s 163813 16328 164613 16448 6 o_din0_1[1]
port 311 nsew signal output
rlabel metal3 s 163813 121728 164613 121848 6 o_din0_1[20]
port 312 nsew signal output
rlabel metal2 s 152646 0 152702 800 6 o_din0_1[21]
port 313 nsew signal output
rlabel metal3 s 0 118328 800 118448 6 o_din0_1[22]
port 314 nsew signal output
rlabel metal3 s 163813 137096 164613 137216 6 o_din0_1[23]
port 315 nsew signal output
rlabel metal2 s 155774 0 155830 800 6 o_din0_1[24]
port 316 nsew signal output
rlabel metal3 s 0 144984 800 145104 6 o_din0_1[25]
port 317 nsew signal output
rlabel metal2 s 156786 0 156842 800 6 o_din0_1[26]
port 318 nsew signal output
rlabel metal2 s 157614 165957 157670 166757 6 o_din0_1[27]
port 319 nsew signal output
rlabel metal2 s 160374 165957 160430 166757 6 o_din0_1[28]
port 320 nsew signal output
rlabel metal2 s 161938 0 161994 800 6 o_din0_1[29]
port 321 nsew signal output
rlabel metal3 s 0 24896 800 25016 6 o_din0_1[2]
port 322 nsew signal output
rlabel metal3 s 163813 163344 164613 163464 6 o_din0_1[30]
port 323 nsew signal output
rlabel metal2 s 162950 0 163006 800 6 o_din0_1[31]
port 324 nsew signal output
rlabel metal3 s 163813 36184 164613 36304 6 o_din0_1[3]
port 325 nsew signal output
rlabel metal2 s 118974 165957 119030 166757 6 o_din0_1[4]
port 326 nsew signal output
rlabel metal3 s 163813 51552 164613 51672 6 o_din0_1[5]
port 327 nsew signal output
rlabel metal3 s 163813 62432 164613 62552 6 o_din0_1[6]
port 328 nsew signal output
rlabel metal2 s 132130 0 132186 800 6 o_din0_1[7]
port 329 nsew signal output
rlabel metal3 s 163813 69096 164613 69216 6 o_din0_1[8]
port 330 nsew signal output
rlabel metal3 s 163813 73448 164613 73568 6 o_din0_1[9]
port 331 nsew signal output
rlabel metal2 s 107934 165957 107990 166757 6 o_waddr0[0]
port 332 nsew signal output
rlabel metal3 s 163813 20816 164613 20936 6 o_waddr0[1]
port 333 nsew signal output
rlabel metal3 s 0 28296 800 28416 6 o_waddr0[2]
port 334 nsew signal output
rlabel metal2 s 115294 165957 115350 166757 6 o_waddr0[3]
port 335 nsew signal output
rlabel metal3 s 0 41624 800 41744 6 o_waddr0[4]
port 336 nsew signal output
rlabel metal3 s 163813 55904 164613 56024 6 o_waddr0[5]
port 337 nsew signal output
rlabel metal2 s 123574 165957 123630 166757 6 o_waddr0[6]
port 338 nsew signal output
rlabel metal3 s 0 58216 800 58336 6 o_waddr0[7]
port 339 nsew signal output
rlabel metal2 s 130014 165957 130070 166757 6 o_waddr0[8]
port 340 nsew signal output
rlabel metal2 s 118698 0 118754 800 6 o_waddr0_1[0]
port 341 nsew signal output
rlabel metal3 s 163813 18640 164613 18760 6 o_waddr0_1[1]
port 342 nsew signal output
rlabel metal3 s 163813 31696 164613 31816 6 o_waddr0_1[2]
port 343 nsew signal output
rlabel metal3 s 163813 38360 164613 38480 6 o_waddr0_1[3]
port 344 nsew signal output
rlabel metal2 s 125966 0 126022 800 6 o_waddr0_1[4]
port 345 nsew signal output
rlabel metal2 s 129002 0 129058 800 6 o_waddr0_1[5]
port 346 nsew signal output
rlabel metal2 s 122654 165957 122710 166757 6 o_waddr0_1[6]
port 347 nsew signal output
rlabel metal2 s 134154 0 134210 800 6 o_waddr0_1[7]
port 348 nsew signal output
rlabel metal2 s 137282 0 137338 800 6 o_waddr0_1[8]
port 349 nsew signal output
rlabel metal3 s 0 1640 800 1760 6 o_web0
port 350 nsew signal output
rlabel metal2 s 112534 0 112590 800 6 o_web0_1
port 351 nsew signal output
rlabel metal3 s 0 4904 800 5024 6 o_wmask0[0]
port 352 nsew signal output
rlabel metal3 s 163813 22992 164613 23112 6 o_wmask0[1]
port 353 nsew signal output
rlabel metal2 s 111614 165957 111670 166757 6 o_wmask0[2]
port 354 nsew signal output
rlabel metal3 s 163813 40536 164613 40656 6 o_wmask0[3]
port 355 nsew signal output
rlabel metal3 s 163813 9800 164613 9920 6 o_wmask0_1[0]
port 356 nsew signal output
rlabel metal3 s 0 11568 800 11688 6 o_wmask0_1[1]
port 357 nsew signal output
rlabel metal3 s 0 31560 800 31680 6 o_wmask0_1[2]
port 358 nsew signal output
rlabel metal2 s 122838 0 122894 800 6 o_wmask0_1[3]
port 359 nsew signal output
rlabel metal4 s 4208 2128 4528 164336 6 vccd1
port 360 nsew power input
rlabel metal4 s 34928 2128 35248 164336 6 vccd1
port 360 nsew power input
rlabel metal4 s 65648 2128 65968 164336 6 vccd1
port 360 nsew power input
rlabel metal4 s 96368 2128 96688 164336 6 vccd1
port 360 nsew power input
rlabel metal4 s 127088 2128 127408 164336 6 vccd1
port 360 nsew power input
rlabel metal4 s 157808 2128 158128 164336 6 vccd1
port 360 nsew power input
rlabel metal4 s 19568 2128 19888 164336 6 vssd1
port 361 nsew ground input
rlabel metal4 s 50288 2128 50608 164336 6 vssd1
port 361 nsew ground input
rlabel metal4 s 81008 2128 81328 164336 6 vssd1
port 361 nsew ground input
rlabel metal4 s 111728 2128 112048 164336 6 vssd1
port 361 nsew ground input
rlabel metal4 s 142448 2128 142768 164336 6 vssd1
port 361 nsew ground input
rlabel metal2 s 478 0 534 800 6 wb_clk_i
port 362 nsew signal input
rlabel metal2 s 1490 0 1546 800 6 wb_rst_i
port 363 nsew signal input
rlabel metal2 s 2502 0 2558 800 6 wbs_ack_o
port 364 nsew signal output
rlabel metal2 s 6642 0 6698 800 6 wbs_adr_i[0]
port 365 nsew signal input
rlabel metal2 s 41602 0 41658 800 6 wbs_adr_i[10]
port 366 nsew signal input
rlabel metal2 s 44638 0 44694 800 6 wbs_adr_i[11]
port 367 nsew signal input
rlabel metal2 s 47766 0 47822 800 6 wbs_adr_i[12]
port 368 nsew signal input
rlabel metal2 s 50802 0 50858 800 6 wbs_adr_i[13]
port 369 nsew signal input
rlabel metal2 s 53930 0 53986 800 6 wbs_adr_i[14]
port 370 nsew signal input
rlabel metal2 s 56966 0 57022 800 6 wbs_adr_i[15]
port 371 nsew signal input
rlabel metal2 s 60094 0 60150 800 6 wbs_adr_i[16]
port 372 nsew signal input
rlabel metal2 s 63222 0 63278 800 6 wbs_adr_i[17]
port 373 nsew signal input
rlabel metal2 s 66258 0 66314 800 6 wbs_adr_i[18]
port 374 nsew signal input
rlabel metal2 s 69386 0 69442 800 6 wbs_adr_i[19]
port 375 nsew signal input
rlabel metal2 s 10690 0 10746 800 6 wbs_adr_i[1]
port 376 nsew signal input
rlabel metal2 s 72422 0 72478 800 6 wbs_adr_i[20]
port 377 nsew signal input
rlabel metal2 s 75550 0 75606 800 6 wbs_adr_i[21]
port 378 nsew signal input
rlabel metal2 s 78586 0 78642 800 6 wbs_adr_i[22]
port 379 nsew signal input
rlabel metal2 s 81714 0 81770 800 6 wbs_adr_i[23]
port 380 nsew signal input
rlabel metal2 s 84750 0 84806 800 6 wbs_adr_i[24]
port 381 nsew signal input
rlabel metal2 s 87878 0 87934 800 6 wbs_adr_i[25]
port 382 nsew signal input
rlabel metal2 s 90914 0 90970 800 6 wbs_adr_i[26]
port 383 nsew signal input
rlabel metal2 s 94042 0 94098 800 6 wbs_adr_i[27]
port 384 nsew signal input
rlabel metal2 s 97170 0 97226 800 6 wbs_adr_i[28]
port 385 nsew signal input
rlabel metal2 s 100206 0 100262 800 6 wbs_adr_i[29]
port 386 nsew signal input
rlabel metal2 s 14830 0 14886 800 6 wbs_adr_i[2]
port 387 nsew signal input
rlabel metal2 s 103334 0 103390 800 6 wbs_adr_i[30]
port 388 nsew signal input
rlabel metal2 s 106370 0 106426 800 6 wbs_adr_i[31]
port 389 nsew signal input
rlabel metal2 s 18970 0 19026 800 6 wbs_adr_i[3]
port 390 nsew signal input
rlabel metal2 s 23018 0 23074 800 6 wbs_adr_i[4]
port 391 nsew signal input
rlabel metal2 s 26146 0 26202 800 6 wbs_adr_i[5]
port 392 nsew signal input
rlabel metal2 s 29274 0 29330 800 6 wbs_adr_i[6]
port 393 nsew signal input
rlabel metal2 s 32310 0 32366 800 6 wbs_adr_i[7]
port 394 nsew signal input
rlabel metal2 s 35438 0 35494 800 6 wbs_adr_i[8]
port 395 nsew signal input
rlabel metal2 s 38474 0 38530 800 6 wbs_adr_i[9]
port 396 nsew signal input
rlabel metal2 s 3514 0 3570 800 6 wbs_cyc_i
port 397 nsew signal input
rlabel metal2 s 7654 0 7710 800 6 wbs_dat_i[0]
port 398 nsew signal input
rlabel metal2 s 42614 0 42670 800 6 wbs_dat_i[10]
port 399 nsew signal input
rlabel metal2 s 45650 0 45706 800 6 wbs_dat_i[11]
port 400 nsew signal input
rlabel metal2 s 48778 0 48834 800 6 wbs_dat_i[12]
port 401 nsew signal input
rlabel metal2 s 51906 0 51962 800 6 wbs_dat_i[13]
port 402 nsew signal input
rlabel metal2 s 54942 0 54998 800 6 wbs_dat_i[14]
port 403 nsew signal input
rlabel metal2 s 58070 0 58126 800 6 wbs_dat_i[15]
port 404 nsew signal input
rlabel metal2 s 61106 0 61162 800 6 wbs_dat_i[16]
port 405 nsew signal input
rlabel metal2 s 64234 0 64290 800 6 wbs_dat_i[17]
port 406 nsew signal input
rlabel metal2 s 67270 0 67326 800 6 wbs_dat_i[18]
port 407 nsew signal input
rlabel metal2 s 70398 0 70454 800 6 wbs_dat_i[19]
port 408 nsew signal input
rlabel metal2 s 11702 0 11758 800 6 wbs_dat_i[1]
port 409 nsew signal input
rlabel metal2 s 73434 0 73490 800 6 wbs_dat_i[20]
port 410 nsew signal input
rlabel metal2 s 76562 0 76618 800 6 wbs_dat_i[21]
port 411 nsew signal input
rlabel metal2 s 79598 0 79654 800 6 wbs_dat_i[22]
port 412 nsew signal input
rlabel metal2 s 82726 0 82782 800 6 wbs_dat_i[23]
port 413 nsew signal input
rlabel metal2 s 85854 0 85910 800 6 wbs_dat_i[24]
port 414 nsew signal input
rlabel metal2 s 88890 0 88946 800 6 wbs_dat_i[25]
port 415 nsew signal input
rlabel metal2 s 92018 0 92074 800 6 wbs_dat_i[26]
port 416 nsew signal input
rlabel metal2 s 95054 0 95110 800 6 wbs_dat_i[27]
port 417 nsew signal input
rlabel metal2 s 98182 0 98238 800 6 wbs_dat_i[28]
port 418 nsew signal input
rlabel metal2 s 101218 0 101274 800 6 wbs_dat_i[29]
port 419 nsew signal input
rlabel metal2 s 15842 0 15898 800 6 wbs_dat_i[2]
port 420 nsew signal input
rlabel metal2 s 104346 0 104402 800 6 wbs_dat_i[30]
port 421 nsew signal input
rlabel metal2 s 107382 0 107438 800 6 wbs_dat_i[31]
port 422 nsew signal input
rlabel metal2 s 19982 0 20038 800 6 wbs_dat_i[3]
port 423 nsew signal input
rlabel metal2 s 24122 0 24178 800 6 wbs_dat_i[4]
port 424 nsew signal input
rlabel metal2 s 27158 0 27214 800 6 wbs_dat_i[5]
port 425 nsew signal input
rlabel metal2 s 30286 0 30342 800 6 wbs_dat_i[6]
port 426 nsew signal input
rlabel metal2 s 33322 0 33378 800 6 wbs_dat_i[7]
port 427 nsew signal input
rlabel metal2 s 36450 0 36506 800 6 wbs_dat_i[8]
port 428 nsew signal input
rlabel metal2 s 39486 0 39542 800 6 wbs_dat_i[9]
port 429 nsew signal input
rlabel metal2 s 8666 0 8722 800 6 wbs_dat_o[0]
port 430 nsew signal output
rlabel metal2 s 43626 0 43682 800 6 wbs_dat_o[10]
port 431 nsew signal output
rlabel metal2 s 46754 0 46810 800 6 wbs_dat_o[11]
port 432 nsew signal output
rlabel metal2 s 49790 0 49846 800 6 wbs_dat_o[12]
port 433 nsew signal output
rlabel metal2 s 52918 0 52974 800 6 wbs_dat_o[13]
port 434 nsew signal output
rlabel metal2 s 55954 0 56010 800 6 wbs_dat_o[14]
port 435 nsew signal output
rlabel metal2 s 59082 0 59138 800 6 wbs_dat_o[15]
port 436 nsew signal output
rlabel metal2 s 62118 0 62174 800 6 wbs_dat_o[16]
port 437 nsew signal output
rlabel metal2 s 65246 0 65302 800 6 wbs_dat_o[17]
port 438 nsew signal output
rlabel metal2 s 68282 0 68338 800 6 wbs_dat_o[18]
port 439 nsew signal output
rlabel metal2 s 71410 0 71466 800 6 wbs_dat_o[19]
port 440 nsew signal output
rlabel metal2 s 12806 0 12862 800 6 wbs_dat_o[1]
port 441 nsew signal output
rlabel metal2 s 74538 0 74594 800 6 wbs_dat_o[20]
port 442 nsew signal output
rlabel metal2 s 77574 0 77630 800 6 wbs_dat_o[21]
port 443 nsew signal output
rlabel metal2 s 80702 0 80758 800 6 wbs_dat_o[22]
port 444 nsew signal output
rlabel metal2 s 83738 0 83794 800 6 wbs_dat_o[23]
port 445 nsew signal output
rlabel metal2 s 86866 0 86922 800 6 wbs_dat_o[24]
port 446 nsew signal output
rlabel metal2 s 89902 0 89958 800 6 wbs_dat_o[25]
port 447 nsew signal output
rlabel metal2 s 93030 0 93086 800 6 wbs_dat_o[26]
port 448 nsew signal output
rlabel metal2 s 96066 0 96122 800 6 wbs_dat_o[27]
port 449 nsew signal output
rlabel metal2 s 99194 0 99250 800 6 wbs_dat_o[28]
port 450 nsew signal output
rlabel metal2 s 102230 0 102286 800 6 wbs_dat_o[29]
port 451 nsew signal output
rlabel metal2 s 16854 0 16910 800 6 wbs_dat_o[2]
port 452 nsew signal output
rlabel metal2 s 105358 0 105414 800 6 wbs_dat_o[30]
port 453 nsew signal output
rlabel metal2 s 108486 0 108542 800 6 wbs_dat_o[31]
port 454 nsew signal output
rlabel metal2 s 20994 0 21050 800 6 wbs_dat_o[3]
port 455 nsew signal output
rlabel metal2 s 25134 0 25190 800 6 wbs_dat_o[4]
port 456 nsew signal output
rlabel metal2 s 28170 0 28226 800 6 wbs_dat_o[5]
port 457 nsew signal output
rlabel metal2 s 31298 0 31354 800 6 wbs_dat_o[6]
port 458 nsew signal output
rlabel metal2 s 34334 0 34390 800 6 wbs_dat_o[7]
port 459 nsew signal output
rlabel metal2 s 37462 0 37518 800 6 wbs_dat_o[8]
port 460 nsew signal output
rlabel metal2 s 40590 0 40646 800 6 wbs_dat_o[9]
port 461 nsew signal output
rlabel metal2 s 9678 0 9734 800 6 wbs_sel_i[0]
port 462 nsew signal input
rlabel metal2 s 13818 0 13874 800 6 wbs_sel_i[1]
port 463 nsew signal input
rlabel metal2 s 17958 0 18014 800 6 wbs_sel_i[2]
port 464 nsew signal input
rlabel metal2 s 22006 0 22062 800 6 wbs_sel_i[3]
port 465 nsew signal input
rlabel metal2 s 4526 0 4582 800 6 wbs_stb_i
port 466 nsew signal input
rlabel metal2 s 5538 0 5594 800 6 wbs_we_i
port 467 nsew signal input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 164613 166757
string LEFview TRUE
string GDS_FILE /local/caravel_user_project/openlane/user_proj/runs/user_proj/results/magic/user_proj.gds
string GDS_END 79824776
string GDS_START 1360742
<< end >>

