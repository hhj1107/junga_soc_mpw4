magic
tech sky130A
magscale 1 2
timestamp 1640405866
<< obsli1 >>
rect 1104 2159 163363 164305
<< obsm1 >>
rect 106 348 163930 164336
<< metal2 >>
rect 478 165721 534 166521
rect 1398 165721 1454 166521
rect 2318 165721 2374 166521
rect 3238 165721 3294 166521
rect 4250 165721 4306 166521
rect 5170 165721 5226 166521
rect 6090 165721 6146 166521
rect 7102 165721 7158 166521
rect 8022 165721 8078 166521
rect 8942 165721 8998 166521
rect 9954 165721 10010 166521
rect 10874 165721 10930 166521
rect 11794 165721 11850 166521
rect 12806 165721 12862 166521
rect 13726 165721 13782 166521
rect 14646 165721 14702 166521
rect 15658 165721 15714 166521
rect 16578 165721 16634 166521
rect 17498 165721 17554 166521
rect 18510 165721 18566 166521
rect 19430 165721 19486 166521
rect 20350 165721 20406 166521
rect 21362 165721 21418 166521
rect 22282 165721 22338 166521
rect 23202 165721 23258 166521
rect 24214 165721 24270 166521
rect 25134 165721 25190 166521
rect 26054 165721 26110 166521
rect 27066 165721 27122 166521
rect 27986 165721 28042 166521
rect 28906 165721 28962 166521
rect 29918 165721 29974 166521
rect 30838 165721 30894 166521
rect 31758 165721 31814 166521
rect 32770 165721 32826 166521
rect 33690 165721 33746 166521
rect 34610 165721 34666 166521
rect 35622 165721 35678 166521
rect 36542 165721 36598 166521
rect 37462 165721 37518 166521
rect 38474 165721 38530 166521
rect 39394 165721 39450 166521
rect 40314 165721 40370 166521
rect 41326 165721 41382 166521
rect 42246 165721 42302 166521
rect 43166 165721 43222 166521
rect 44178 165721 44234 166521
rect 45098 165721 45154 166521
rect 46018 165721 46074 166521
rect 47030 165721 47086 166521
rect 47950 165721 48006 166521
rect 48870 165721 48926 166521
rect 49882 165721 49938 166521
rect 50802 165721 50858 166521
rect 51722 165721 51778 166521
rect 52734 165721 52790 166521
rect 53654 165721 53710 166521
rect 54574 165721 54630 166521
rect 55586 165721 55642 166521
rect 56506 165721 56562 166521
rect 57426 165721 57482 166521
rect 58438 165721 58494 166521
rect 59358 165721 59414 166521
rect 60278 165721 60334 166521
rect 61290 165721 61346 166521
rect 62210 165721 62266 166521
rect 63130 165721 63186 166521
rect 64142 165721 64198 166521
rect 65062 165721 65118 166521
rect 65982 165721 66038 166521
rect 66994 165721 67050 166521
rect 67914 165721 67970 166521
rect 68834 165721 68890 166521
rect 69846 165721 69902 166521
rect 70766 165721 70822 166521
rect 71686 165721 71742 166521
rect 72698 165721 72754 166521
rect 73618 165721 73674 166521
rect 74538 165721 74594 166521
rect 75550 165721 75606 166521
rect 76470 165721 76526 166521
rect 77390 165721 77446 166521
rect 78402 165721 78458 166521
rect 79322 165721 79378 166521
rect 80242 165721 80298 166521
rect 81254 165721 81310 166521
rect 82174 165721 82230 166521
rect 83094 165721 83150 166521
rect 84014 165721 84070 166521
rect 85026 165721 85082 166521
rect 85946 165721 86002 166521
rect 86866 165721 86922 166521
rect 87878 165721 87934 166521
rect 88798 165721 88854 166521
rect 89718 165721 89774 166521
rect 90730 165721 90786 166521
rect 91650 165721 91706 166521
rect 92570 165721 92626 166521
rect 93582 165721 93638 166521
rect 94502 165721 94558 166521
rect 95422 165721 95478 166521
rect 96434 165721 96490 166521
rect 97354 165721 97410 166521
rect 98274 165721 98330 166521
rect 99286 165721 99342 166521
rect 100206 165721 100262 166521
rect 101126 165721 101182 166521
rect 102138 165721 102194 166521
rect 103058 165721 103114 166521
rect 103978 165721 104034 166521
rect 104990 165721 105046 166521
rect 105910 165721 105966 166521
rect 106830 165721 106886 166521
rect 107842 165721 107898 166521
rect 108762 165721 108818 166521
rect 109682 165721 109738 166521
rect 110694 165721 110750 166521
rect 111614 165721 111670 166521
rect 112534 165721 112590 166521
rect 113546 165721 113602 166521
rect 114466 165721 114522 166521
rect 115386 165721 115442 166521
rect 116398 165721 116454 166521
rect 117318 165721 117374 166521
rect 118238 165721 118294 166521
rect 119250 165721 119306 166521
rect 120170 165721 120226 166521
rect 121090 165721 121146 166521
rect 122102 165721 122158 166521
rect 123022 165721 123078 166521
rect 123942 165721 123998 166521
rect 124954 165721 125010 166521
rect 125874 165721 125930 166521
rect 126794 165721 126850 166521
rect 127806 165721 127862 166521
rect 128726 165721 128782 166521
rect 129646 165721 129702 166521
rect 130658 165721 130714 166521
rect 131578 165721 131634 166521
rect 132498 165721 132554 166521
rect 133510 165721 133566 166521
rect 134430 165721 134486 166521
rect 135350 165721 135406 166521
rect 136362 165721 136418 166521
rect 137282 165721 137338 166521
rect 138202 165721 138258 166521
rect 139214 165721 139270 166521
rect 140134 165721 140190 166521
rect 141054 165721 141110 166521
rect 142066 165721 142122 166521
rect 142986 165721 143042 166521
rect 143906 165721 143962 166521
rect 144918 165721 144974 166521
rect 145838 165721 145894 166521
rect 146758 165721 146814 166521
rect 147770 165721 147826 166521
rect 148690 165721 148746 166521
rect 149610 165721 149666 166521
rect 150622 165721 150678 166521
rect 151542 165721 151598 166521
rect 152462 165721 152518 166521
rect 153474 165721 153530 166521
rect 154394 165721 154450 166521
rect 155314 165721 155370 166521
rect 156326 165721 156382 166521
rect 157246 165721 157302 166521
rect 158166 165721 158222 166521
rect 159178 165721 159234 166521
rect 160098 165721 160154 166521
rect 161018 165721 161074 166521
rect 162030 165721 162086 166521
rect 162950 165721 163006 166521
rect 163870 165721 163926 166521
rect 478 0 534 800
rect 1398 0 1454 800
rect 2410 0 2466 800
rect 3422 0 3478 800
rect 4434 0 4490 800
rect 5354 0 5410 800
rect 6366 0 6422 800
rect 7378 0 7434 800
rect 8390 0 8446 800
rect 9310 0 9366 800
rect 10322 0 10378 800
rect 11334 0 11390 800
rect 12346 0 12402 800
rect 13266 0 13322 800
rect 14278 0 14334 800
rect 15290 0 15346 800
rect 16302 0 16358 800
rect 17314 0 17370 800
rect 18234 0 18290 800
rect 19246 0 19302 800
rect 20258 0 20314 800
rect 21270 0 21326 800
rect 22190 0 22246 800
rect 23202 0 23258 800
rect 24214 0 24270 800
rect 25226 0 25282 800
rect 26146 0 26202 800
rect 27158 0 27214 800
rect 28170 0 28226 800
rect 29182 0 29238 800
rect 30102 0 30158 800
rect 31114 0 31170 800
rect 32126 0 32182 800
rect 33138 0 33194 800
rect 34150 0 34206 800
rect 35070 0 35126 800
rect 36082 0 36138 800
rect 37094 0 37150 800
rect 38106 0 38162 800
rect 39026 0 39082 800
rect 40038 0 40094 800
rect 41050 0 41106 800
rect 42062 0 42118 800
rect 42982 0 43038 800
rect 43994 0 44050 800
rect 45006 0 45062 800
rect 46018 0 46074 800
rect 46938 0 46994 800
rect 47950 0 48006 800
rect 48962 0 49018 800
rect 49974 0 50030 800
rect 50986 0 51042 800
rect 51906 0 51962 800
rect 52918 0 52974 800
rect 53930 0 53986 800
rect 54942 0 54998 800
rect 55862 0 55918 800
rect 56874 0 56930 800
rect 57886 0 57942 800
rect 58898 0 58954 800
rect 59818 0 59874 800
rect 60830 0 60886 800
rect 61842 0 61898 800
rect 62854 0 62910 800
rect 63774 0 63830 800
rect 64786 0 64842 800
rect 65798 0 65854 800
rect 66810 0 66866 800
rect 67822 0 67878 800
rect 68742 0 68798 800
rect 69754 0 69810 800
rect 70766 0 70822 800
rect 71778 0 71834 800
rect 72698 0 72754 800
rect 73710 0 73766 800
rect 74722 0 74778 800
rect 75734 0 75790 800
rect 76654 0 76710 800
rect 77666 0 77722 800
rect 78678 0 78734 800
rect 79690 0 79746 800
rect 80610 0 80666 800
rect 81622 0 81678 800
rect 82634 0 82690 800
rect 83646 0 83702 800
rect 84658 0 84714 800
rect 85578 0 85634 800
rect 86590 0 86646 800
rect 87602 0 87658 800
rect 88614 0 88670 800
rect 89534 0 89590 800
rect 90546 0 90602 800
rect 91558 0 91614 800
rect 92570 0 92626 800
rect 93490 0 93546 800
rect 94502 0 94558 800
rect 95514 0 95570 800
rect 96526 0 96582 800
rect 97446 0 97502 800
rect 98458 0 98514 800
rect 99470 0 99526 800
rect 100482 0 100538 800
rect 101494 0 101550 800
rect 102414 0 102470 800
rect 103426 0 103482 800
rect 104438 0 104494 800
rect 105450 0 105506 800
rect 106370 0 106426 800
rect 107382 0 107438 800
rect 108394 0 108450 800
rect 109406 0 109462 800
rect 110326 0 110382 800
rect 111338 0 111394 800
rect 112350 0 112406 800
rect 113362 0 113418 800
rect 114282 0 114338 800
rect 115294 0 115350 800
rect 116306 0 116362 800
rect 117318 0 117374 800
rect 118330 0 118386 800
rect 119250 0 119306 800
rect 120262 0 120318 800
rect 121274 0 121330 800
rect 122286 0 122342 800
rect 123206 0 123262 800
rect 124218 0 124274 800
rect 125230 0 125286 800
rect 126242 0 126298 800
rect 127162 0 127218 800
rect 128174 0 128230 800
rect 129186 0 129242 800
rect 130198 0 130254 800
rect 131118 0 131174 800
rect 132130 0 132186 800
rect 133142 0 133198 800
rect 134154 0 134210 800
rect 135166 0 135222 800
rect 136086 0 136142 800
rect 137098 0 137154 800
rect 138110 0 138166 800
rect 139122 0 139178 800
rect 140042 0 140098 800
rect 141054 0 141110 800
rect 142066 0 142122 800
rect 143078 0 143134 800
rect 143998 0 144054 800
rect 145010 0 145066 800
rect 146022 0 146078 800
rect 147034 0 147090 800
rect 147954 0 148010 800
rect 148966 0 149022 800
rect 149978 0 150034 800
rect 150990 0 151046 800
rect 152002 0 152058 800
rect 152922 0 152978 800
rect 153934 0 153990 800
rect 154946 0 155002 800
rect 155958 0 156014 800
rect 156878 0 156934 800
rect 157890 0 157946 800
rect 158902 0 158958 800
rect 159914 0 159970 800
rect 160834 0 160890 800
rect 161846 0 161902 800
rect 162858 0 162914 800
rect 163870 0 163926 800
<< obsm2 >>
rect 112 165665 422 165866
rect 590 165665 1342 165866
rect 1510 165665 2262 165866
rect 2430 165665 3182 165866
rect 3350 165665 4194 165866
rect 4362 165665 5114 165866
rect 5282 165665 6034 165866
rect 6202 165665 7046 165866
rect 7214 165665 7966 165866
rect 8134 165665 8886 165866
rect 9054 165665 9898 165866
rect 10066 165665 10818 165866
rect 10986 165665 11738 165866
rect 11906 165665 12750 165866
rect 12918 165665 13670 165866
rect 13838 165665 14590 165866
rect 14758 165665 15602 165866
rect 15770 165665 16522 165866
rect 16690 165665 17442 165866
rect 17610 165665 18454 165866
rect 18622 165665 19374 165866
rect 19542 165665 20294 165866
rect 20462 165665 21306 165866
rect 21474 165665 22226 165866
rect 22394 165665 23146 165866
rect 23314 165665 24158 165866
rect 24326 165665 25078 165866
rect 25246 165665 25998 165866
rect 26166 165665 27010 165866
rect 27178 165665 27930 165866
rect 28098 165665 28850 165866
rect 29018 165665 29862 165866
rect 30030 165665 30782 165866
rect 30950 165665 31702 165866
rect 31870 165665 32714 165866
rect 32882 165665 33634 165866
rect 33802 165665 34554 165866
rect 34722 165665 35566 165866
rect 35734 165665 36486 165866
rect 36654 165665 37406 165866
rect 37574 165665 38418 165866
rect 38586 165665 39338 165866
rect 39506 165665 40258 165866
rect 40426 165665 41270 165866
rect 41438 165665 42190 165866
rect 42358 165665 43110 165866
rect 43278 165665 44122 165866
rect 44290 165665 45042 165866
rect 45210 165665 45962 165866
rect 46130 165665 46974 165866
rect 47142 165665 47894 165866
rect 48062 165665 48814 165866
rect 48982 165665 49826 165866
rect 49994 165665 50746 165866
rect 50914 165665 51666 165866
rect 51834 165665 52678 165866
rect 52846 165665 53598 165866
rect 53766 165665 54518 165866
rect 54686 165665 55530 165866
rect 55698 165665 56450 165866
rect 56618 165665 57370 165866
rect 57538 165665 58382 165866
rect 58550 165665 59302 165866
rect 59470 165665 60222 165866
rect 60390 165665 61234 165866
rect 61402 165665 62154 165866
rect 62322 165665 63074 165866
rect 63242 165665 64086 165866
rect 64254 165665 65006 165866
rect 65174 165665 65926 165866
rect 66094 165665 66938 165866
rect 67106 165665 67858 165866
rect 68026 165665 68778 165866
rect 68946 165665 69790 165866
rect 69958 165665 70710 165866
rect 70878 165665 71630 165866
rect 71798 165665 72642 165866
rect 72810 165665 73562 165866
rect 73730 165665 74482 165866
rect 74650 165665 75494 165866
rect 75662 165665 76414 165866
rect 76582 165665 77334 165866
rect 77502 165665 78346 165866
rect 78514 165665 79266 165866
rect 79434 165665 80186 165866
rect 80354 165665 81198 165866
rect 81366 165665 82118 165866
rect 82286 165665 83038 165866
rect 83206 165665 83958 165866
rect 84126 165665 84970 165866
rect 85138 165665 85890 165866
rect 86058 165665 86810 165866
rect 86978 165665 87822 165866
rect 87990 165665 88742 165866
rect 88910 165665 89662 165866
rect 89830 165665 90674 165866
rect 90842 165665 91594 165866
rect 91762 165665 92514 165866
rect 92682 165665 93526 165866
rect 93694 165665 94446 165866
rect 94614 165665 95366 165866
rect 95534 165665 96378 165866
rect 96546 165665 97298 165866
rect 97466 165665 98218 165866
rect 98386 165665 99230 165866
rect 99398 165665 100150 165866
rect 100318 165665 101070 165866
rect 101238 165665 102082 165866
rect 102250 165665 103002 165866
rect 103170 165665 103922 165866
rect 104090 165665 104934 165866
rect 105102 165665 105854 165866
rect 106022 165665 106774 165866
rect 106942 165665 107786 165866
rect 107954 165665 108706 165866
rect 108874 165665 109626 165866
rect 109794 165665 110638 165866
rect 110806 165665 111558 165866
rect 111726 165665 112478 165866
rect 112646 165665 113490 165866
rect 113658 165665 114410 165866
rect 114578 165665 115330 165866
rect 115498 165665 116342 165866
rect 116510 165665 117262 165866
rect 117430 165665 118182 165866
rect 118350 165665 119194 165866
rect 119362 165665 120114 165866
rect 120282 165665 121034 165866
rect 121202 165665 122046 165866
rect 122214 165665 122966 165866
rect 123134 165665 123886 165866
rect 124054 165665 124898 165866
rect 125066 165665 125818 165866
rect 125986 165665 126738 165866
rect 126906 165665 127750 165866
rect 127918 165665 128670 165866
rect 128838 165665 129590 165866
rect 129758 165665 130602 165866
rect 130770 165665 131522 165866
rect 131690 165665 132442 165866
rect 132610 165665 133454 165866
rect 133622 165665 134374 165866
rect 134542 165665 135294 165866
rect 135462 165665 136306 165866
rect 136474 165665 137226 165866
rect 137394 165665 138146 165866
rect 138314 165665 139158 165866
rect 139326 165665 140078 165866
rect 140246 165665 140998 165866
rect 141166 165665 142010 165866
rect 142178 165665 142930 165866
rect 143098 165665 143850 165866
rect 144018 165665 144862 165866
rect 145030 165665 145782 165866
rect 145950 165665 146702 165866
rect 146870 165665 147714 165866
rect 147882 165665 148634 165866
rect 148802 165665 149554 165866
rect 149722 165665 150566 165866
rect 150734 165665 151486 165866
rect 151654 165665 152406 165866
rect 152574 165665 153418 165866
rect 153586 165665 154338 165866
rect 154506 165665 155258 165866
rect 155426 165665 156270 165866
rect 156438 165665 157190 165866
rect 157358 165665 158110 165866
rect 158278 165665 159122 165866
rect 159290 165665 160042 165866
rect 160210 165665 160962 165866
rect 161130 165665 161974 165866
rect 162142 165665 162894 165866
rect 163062 165665 163814 165866
rect 112 856 163924 165665
rect 112 342 422 856
rect 590 342 1342 856
rect 1510 342 2354 856
rect 2522 342 3366 856
rect 3534 342 4378 856
rect 4546 342 5298 856
rect 5466 342 6310 856
rect 6478 342 7322 856
rect 7490 342 8334 856
rect 8502 342 9254 856
rect 9422 342 10266 856
rect 10434 342 11278 856
rect 11446 342 12290 856
rect 12458 342 13210 856
rect 13378 342 14222 856
rect 14390 342 15234 856
rect 15402 342 16246 856
rect 16414 342 17258 856
rect 17426 342 18178 856
rect 18346 342 19190 856
rect 19358 342 20202 856
rect 20370 342 21214 856
rect 21382 342 22134 856
rect 22302 342 23146 856
rect 23314 342 24158 856
rect 24326 342 25170 856
rect 25338 342 26090 856
rect 26258 342 27102 856
rect 27270 342 28114 856
rect 28282 342 29126 856
rect 29294 342 30046 856
rect 30214 342 31058 856
rect 31226 342 32070 856
rect 32238 342 33082 856
rect 33250 342 34094 856
rect 34262 342 35014 856
rect 35182 342 36026 856
rect 36194 342 37038 856
rect 37206 342 38050 856
rect 38218 342 38970 856
rect 39138 342 39982 856
rect 40150 342 40994 856
rect 41162 342 42006 856
rect 42174 342 42926 856
rect 43094 342 43938 856
rect 44106 342 44950 856
rect 45118 342 45962 856
rect 46130 342 46882 856
rect 47050 342 47894 856
rect 48062 342 48906 856
rect 49074 342 49918 856
rect 50086 342 50930 856
rect 51098 342 51850 856
rect 52018 342 52862 856
rect 53030 342 53874 856
rect 54042 342 54886 856
rect 55054 342 55806 856
rect 55974 342 56818 856
rect 56986 342 57830 856
rect 57998 342 58842 856
rect 59010 342 59762 856
rect 59930 342 60774 856
rect 60942 342 61786 856
rect 61954 342 62798 856
rect 62966 342 63718 856
rect 63886 342 64730 856
rect 64898 342 65742 856
rect 65910 342 66754 856
rect 66922 342 67766 856
rect 67934 342 68686 856
rect 68854 342 69698 856
rect 69866 342 70710 856
rect 70878 342 71722 856
rect 71890 342 72642 856
rect 72810 342 73654 856
rect 73822 342 74666 856
rect 74834 342 75678 856
rect 75846 342 76598 856
rect 76766 342 77610 856
rect 77778 342 78622 856
rect 78790 342 79634 856
rect 79802 342 80554 856
rect 80722 342 81566 856
rect 81734 342 82578 856
rect 82746 342 83590 856
rect 83758 342 84602 856
rect 84770 342 85522 856
rect 85690 342 86534 856
rect 86702 342 87546 856
rect 87714 342 88558 856
rect 88726 342 89478 856
rect 89646 342 90490 856
rect 90658 342 91502 856
rect 91670 342 92514 856
rect 92682 342 93434 856
rect 93602 342 94446 856
rect 94614 342 95458 856
rect 95626 342 96470 856
rect 96638 342 97390 856
rect 97558 342 98402 856
rect 98570 342 99414 856
rect 99582 342 100426 856
rect 100594 342 101438 856
rect 101606 342 102358 856
rect 102526 342 103370 856
rect 103538 342 104382 856
rect 104550 342 105394 856
rect 105562 342 106314 856
rect 106482 342 107326 856
rect 107494 342 108338 856
rect 108506 342 109350 856
rect 109518 342 110270 856
rect 110438 342 111282 856
rect 111450 342 112294 856
rect 112462 342 113306 856
rect 113474 342 114226 856
rect 114394 342 115238 856
rect 115406 342 116250 856
rect 116418 342 117262 856
rect 117430 342 118274 856
rect 118442 342 119194 856
rect 119362 342 120206 856
rect 120374 342 121218 856
rect 121386 342 122230 856
rect 122398 342 123150 856
rect 123318 342 124162 856
rect 124330 342 125174 856
rect 125342 342 126186 856
rect 126354 342 127106 856
rect 127274 342 128118 856
rect 128286 342 129130 856
rect 129298 342 130142 856
rect 130310 342 131062 856
rect 131230 342 132074 856
rect 132242 342 133086 856
rect 133254 342 134098 856
rect 134266 342 135110 856
rect 135278 342 136030 856
rect 136198 342 137042 856
rect 137210 342 138054 856
rect 138222 342 139066 856
rect 139234 342 139986 856
rect 140154 342 140998 856
rect 141166 342 142010 856
rect 142178 342 143022 856
rect 143190 342 143942 856
rect 144110 342 144954 856
rect 145122 342 145966 856
rect 146134 342 146978 856
rect 147146 342 147898 856
rect 148066 342 148910 856
rect 149078 342 149922 856
rect 150090 342 150934 856
rect 151102 342 151946 856
rect 152114 342 152866 856
rect 153034 342 153878 856
rect 154046 342 154890 856
rect 155058 342 155902 856
rect 156070 342 156822 856
rect 156990 342 157834 856
rect 158002 342 158846 856
rect 159014 342 159858 856
rect 160026 342 160778 856
rect 160946 342 161790 856
rect 161958 342 162802 856
rect 162970 342 163814 856
<< metal3 >>
rect 163577 165112 164377 165232
rect 0 164840 800 164960
rect 163577 162664 164377 162784
rect 0 161984 800 162104
rect 163577 160216 164377 160336
rect 0 158992 800 159112
rect 163577 157904 164377 158024
rect 0 156136 800 156256
rect 163577 155456 164377 155576
rect 0 153144 800 153264
rect 163577 153008 164377 153128
rect 163577 150560 164377 150680
rect 0 150288 800 150408
rect 163577 148248 164377 148368
rect 0 147296 800 147416
rect 163577 145800 164377 145920
rect 0 144440 800 144560
rect 163577 143352 164377 143472
rect 0 141448 800 141568
rect 163577 140904 164377 141024
rect 0 138592 800 138712
rect 163577 138592 164377 138712
rect 163577 136144 164377 136264
rect 0 135600 800 135720
rect 163577 133696 164377 133816
rect 0 132744 800 132864
rect 163577 131248 164377 131368
rect 0 129752 800 129872
rect 163577 128936 164377 129056
rect 0 126896 800 127016
rect 163577 126488 164377 126608
rect 0 123904 800 124024
rect 163577 124040 164377 124160
rect 163577 121592 164377 121712
rect 0 121048 800 121168
rect 163577 119280 164377 119400
rect 0 118056 800 118176
rect 163577 116832 164377 116952
rect 0 115200 800 115320
rect 163577 114384 164377 114504
rect 0 112344 800 112464
rect 163577 112072 164377 112192
rect 163577 109624 164377 109744
rect 0 109352 800 109472
rect 163577 107176 164377 107296
rect 0 106496 800 106616
rect 163577 104728 164377 104848
rect 0 103504 800 103624
rect 163577 102416 164377 102536
rect 0 100648 800 100768
rect 163577 99968 164377 100088
rect 0 97656 800 97776
rect 163577 97520 164377 97640
rect 163577 95072 164377 95192
rect 0 94800 800 94920
rect 163577 92760 164377 92880
rect 0 91808 800 91928
rect 163577 90312 164377 90432
rect 0 88952 800 89072
rect 163577 87864 164377 87984
rect 0 85960 800 86080
rect 163577 85416 164377 85536
rect 0 83104 800 83224
rect 163577 83104 164377 83224
rect 163577 80656 164377 80776
rect 0 80112 800 80232
rect 163577 78208 164377 78328
rect 0 77256 800 77376
rect 163577 75760 164377 75880
rect 0 74264 800 74384
rect 163577 73448 164377 73568
rect 0 71408 800 71528
rect 163577 71000 164377 71120
rect 0 68416 800 68536
rect 163577 68552 164377 68672
rect 163577 66104 164377 66224
rect 0 65560 800 65680
rect 163577 63792 164377 63912
rect 0 62568 800 62688
rect 163577 61344 164377 61464
rect 0 59712 800 59832
rect 163577 58896 164377 59016
rect 0 56856 800 56976
rect 163577 56584 164377 56704
rect 163577 54136 164377 54256
rect 0 53864 800 53984
rect 163577 51688 164377 51808
rect 0 51008 800 51128
rect 163577 49240 164377 49360
rect 0 48016 800 48136
rect 163577 46928 164377 47048
rect 0 45160 800 45280
rect 163577 44480 164377 44600
rect 0 42168 800 42288
rect 163577 42032 164377 42152
rect 163577 39584 164377 39704
rect 0 39312 800 39432
rect 163577 37272 164377 37392
rect 0 36320 800 36440
rect 163577 34824 164377 34944
rect 0 33464 800 33584
rect 163577 32376 164377 32496
rect 0 30472 800 30592
rect 163577 29928 164377 30048
rect 0 27616 800 27736
rect 163577 27616 164377 27736
rect 163577 25168 164377 25288
rect 0 24624 800 24744
rect 163577 22720 164377 22840
rect 0 21768 800 21888
rect 163577 20272 164377 20392
rect 0 18776 800 18896
rect 163577 17960 164377 18080
rect 0 15920 800 16040
rect 163577 15512 164377 15632
rect 0 12928 800 13048
rect 163577 13064 164377 13184
rect 163577 10616 164377 10736
rect 0 10072 800 10192
rect 163577 8304 164377 8424
rect 0 7080 800 7200
rect 163577 5856 164377 5976
rect 0 4224 800 4344
rect 163577 3408 164377 3528
rect 0 1368 800 1488
rect 163577 1096 164377 1216
<< obsm3 >>
rect 197 162864 163577 164321
rect 197 162584 163497 162864
rect 197 162184 163577 162584
rect 880 161904 163577 162184
rect 197 160416 163577 161904
rect 197 160136 163497 160416
rect 197 159192 163577 160136
rect 880 158912 163577 159192
rect 197 158104 163577 158912
rect 197 157824 163497 158104
rect 197 156336 163577 157824
rect 880 156056 163577 156336
rect 197 155656 163577 156056
rect 197 155376 163497 155656
rect 197 153344 163577 155376
rect 880 153208 163577 153344
rect 880 153064 163497 153208
rect 197 152928 163497 153064
rect 197 150760 163577 152928
rect 197 150488 163497 150760
rect 880 150480 163497 150488
rect 880 150208 163577 150480
rect 197 148448 163577 150208
rect 197 148168 163497 148448
rect 197 147496 163577 148168
rect 880 147216 163577 147496
rect 197 146000 163577 147216
rect 197 145720 163497 146000
rect 197 144640 163577 145720
rect 880 144360 163577 144640
rect 197 143552 163577 144360
rect 197 143272 163497 143552
rect 197 141648 163577 143272
rect 880 141368 163577 141648
rect 197 141104 163577 141368
rect 197 140824 163497 141104
rect 197 138792 163577 140824
rect 880 138512 163497 138792
rect 197 136344 163577 138512
rect 197 136064 163497 136344
rect 197 135800 163577 136064
rect 880 135520 163577 135800
rect 197 133896 163577 135520
rect 197 133616 163497 133896
rect 197 132944 163577 133616
rect 880 132664 163577 132944
rect 197 131448 163577 132664
rect 197 131168 163497 131448
rect 197 129952 163577 131168
rect 880 129672 163577 129952
rect 197 129136 163577 129672
rect 197 128856 163497 129136
rect 197 127096 163577 128856
rect 880 126816 163577 127096
rect 197 126688 163577 126816
rect 197 126408 163497 126688
rect 197 124240 163577 126408
rect 197 124104 163497 124240
rect 880 123960 163497 124104
rect 880 123824 163577 123960
rect 197 121792 163577 123824
rect 197 121512 163497 121792
rect 197 121248 163577 121512
rect 880 120968 163577 121248
rect 197 119480 163577 120968
rect 197 119200 163497 119480
rect 197 118256 163577 119200
rect 880 117976 163577 118256
rect 197 117032 163577 117976
rect 197 116752 163497 117032
rect 197 115400 163577 116752
rect 880 115120 163577 115400
rect 197 114584 163577 115120
rect 197 114304 163497 114584
rect 197 112544 163577 114304
rect 880 112272 163577 112544
rect 880 112264 163497 112272
rect 197 111992 163497 112264
rect 197 109824 163577 111992
rect 197 109552 163497 109824
rect 880 109544 163497 109552
rect 880 109272 163577 109544
rect 197 107376 163577 109272
rect 197 107096 163497 107376
rect 197 106696 163577 107096
rect 880 106416 163577 106696
rect 197 104928 163577 106416
rect 197 104648 163497 104928
rect 197 103704 163577 104648
rect 880 103424 163577 103704
rect 197 102616 163577 103424
rect 197 102336 163497 102616
rect 197 100848 163577 102336
rect 880 100568 163577 100848
rect 197 100168 163577 100568
rect 197 99888 163497 100168
rect 197 97856 163577 99888
rect 880 97720 163577 97856
rect 880 97576 163497 97720
rect 197 97440 163497 97576
rect 197 95272 163577 97440
rect 197 95000 163497 95272
rect 880 94992 163497 95000
rect 880 94720 163577 94992
rect 197 92960 163577 94720
rect 197 92680 163497 92960
rect 197 92008 163577 92680
rect 880 91728 163577 92008
rect 197 90512 163577 91728
rect 197 90232 163497 90512
rect 197 89152 163577 90232
rect 880 88872 163577 89152
rect 197 88064 163577 88872
rect 197 87784 163497 88064
rect 197 86160 163577 87784
rect 880 85880 163577 86160
rect 197 85616 163577 85880
rect 197 85336 163497 85616
rect 197 83304 163577 85336
rect 880 83024 163497 83304
rect 197 80856 163577 83024
rect 197 80576 163497 80856
rect 197 80312 163577 80576
rect 880 80032 163577 80312
rect 197 78408 163577 80032
rect 197 78128 163497 78408
rect 197 77456 163577 78128
rect 880 77176 163577 77456
rect 197 75960 163577 77176
rect 197 75680 163497 75960
rect 197 74464 163577 75680
rect 880 74184 163577 74464
rect 197 73648 163577 74184
rect 197 73368 163497 73648
rect 197 71608 163577 73368
rect 880 71328 163577 71608
rect 197 71200 163577 71328
rect 197 70920 163497 71200
rect 197 68752 163577 70920
rect 197 68616 163497 68752
rect 880 68472 163497 68616
rect 880 68336 163577 68472
rect 197 66304 163577 68336
rect 197 66024 163497 66304
rect 197 65760 163577 66024
rect 880 65480 163577 65760
rect 197 63992 163577 65480
rect 197 63712 163497 63992
rect 197 62768 163577 63712
rect 880 62488 163577 62768
rect 197 61544 163577 62488
rect 197 61264 163497 61544
rect 197 59912 163577 61264
rect 880 59632 163577 59912
rect 197 59096 163577 59632
rect 197 58816 163497 59096
rect 197 57056 163577 58816
rect 880 56784 163577 57056
rect 880 56776 163497 56784
rect 197 56504 163497 56776
rect 197 54336 163577 56504
rect 197 54064 163497 54336
rect 880 54056 163497 54064
rect 880 53784 163577 54056
rect 197 51888 163577 53784
rect 197 51608 163497 51888
rect 197 51208 163577 51608
rect 880 50928 163577 51208
rect 197 49440 163577 50928
rect 197 49160 163497 49440
rect 197 48216 163577 49160
rect 880 47936 163577 48216
rect 197 47128 163577 47936
rect 197 46848 163497 47128
rect 197 45360 163577 46848
rect 880 45080 163577 45360
rect 197 44680 163577 45080
rect 197 44400 163497 44680
rect 197 42368 163577 44400
rect 880 42232 163577 42368
rect 880 42088 163497 42232
rect 197 41952 163497 42088
rect 197 39784 163577 41952
rect 197 39512 163497 39784
rect 880 39504 163497 39512
rect 880 39232 163577 39504
rect 197 37472 163577 39232
rect 197 37192 163497 37472
rect 197 36520 163577 37192
rect 880 36240 163577 36520
rect 197 35024 163577 36240
rect 197 34744 163497 35024
rect 197 33664 163577 34744
rect 880 33384 163577 33664
rect 197 32576 163577 33384
rect 197 32296 163497 32576
rect 197 30672 163577 32296
rect 880 30392 163577 30672
rect 197 30128 163577 30392
rect 197 29848 163497 30128
rect 197 27816 163577 29848
rect 880 27536 163497 27816
rect 197 25368 163577 27536
rect 197 25088 163497 25368
rect 197 24824 163577 25088
rect 880 24544 163577 24824
rect 197 22920 163577 24544
rect 197 22640 163497 22920
rect 197 21968 163577 22640
rect 880 21688 163577 21968
rect 197 20472 163577 21688
rect 197 20192 163497 20472
rect 197 18976 163577 20192
rect 880 18696 163577 18976
rect 197 18160 163577 18696
rect 197 17880 163497 18160
rect 197 16120 163577 17880
rect 880 15840 163577 16120
rect 197 15712 163577 15840
rect 197 15432 163497 15712
rect 197 13264 163577 15432
rect 197 13128 163497 13264
rect 880 12984 163497 13128
rect 880 12848 163577 12984
rect 197 10816 163577 12848
rect 197 10536 163497 10816
rect 197 10272 163577 10536
rect 880 9992 163577 10272
rect 197 8504 163577 9992
rect 197 8224 163497 8504
rect 197 7280 163577 8224
rect 880 7000 163577 7280
rect 197 6056 163577 7000
rect 197 5776 163497 6056
rect 197 4424 163577 5776
rect 880 4144 163577 4424
rect 197 3608 163577 4144
rect 197 3328 163497 3608
rect 197 1568 163577 3328
rect 880 1296 163577 1568
rect 880 1288 163497 1296
rect 197 1016 163497 1288
rect 197 579 163577 1016
<< metal4 >>
rect 4208 2128 4528 164336
rect 19568 2128 19888 164336
rect 34928 2128 35248 164336
rect 50288 2128 50608 164336
rect 65648 2128 65968 164336
rect 81008 2128 81328 164336
rect 96368 2128 96688 164336
rect 111728 2128 112048 164336
rect 127088 2128 127408 164336
rect 142448 2128 142768 164336
rect 157808 2128 158128 164336
<< obsm4 >>
rect 243 2048 4128 164117
rect 4608 2048 19488 164117
rect 19968 2048 34848 164117
rect 35328 2048 50208 164117
rect 50688 2048 65568 164117
rect 66048 2048 80928 164117
rect 81408 2048 96288 164117
rect 96768 2048 111648 164117
rect 112128 2048 127008 164117
rect 127488 2048 142368 164117
rect 142848 2048 157629 164117
rect 243 579 157629 2048
<< labels >>
rlabel metal2 s 110694 165721 110750 166521 6 i_dout0[0]
port 1 nsew signal input
rlabel metal3 s 163577 75760 164377 75880 6 i_dout0[10]
port 2 nsew signal input
rlabel metal3 s 163577 83104 164377 83224 6 i_dout0[11]
port 3 nsew signal input
rlabel metal2 s 137098 0 137154 800 6 i_dout0[12]
port 4 nsew signal input
rlabel metal3 s 163577 90312 164377 90432 6 i_dout0[13]
port 5 nsew signal input
rlabel metal2 s 142066 165721 142122 166521 6 i_dout0[14]
port 6 nsew signal input
rlabel metal2 s 141054 0 141110 800 6 i_dout0[15]
port 7 nsew signal input
rlabel metal3 s 163577 99968 164377 100088 6 i_dout0[16]
port 8 nsew signal input
rlabel metal2 s 145838 165721 145894 166521 6 i_dout0[17]
port 9 nsew signal input
rlabel metal3 s 163577 109624 164377 109744 6 i_dout0[18]
port 10 nsew signal input
rlabel metal2 s 147770 165721 147826 166521 6 i_dout0[19]
port 11 nsew signal input
rlabel metal3 s 163577 13064 164377 13184 6 i_dout0[1]
port 12 nsew signal input
rlabel metal2 s 149610 165721 149666 166521 6 i_dout0[20]
port 13 nsew signal input
rlabel metal2 s 149978 0 150034 800 6 i_dout0[21]
port 14 nsew signal input
rlabel metal2 s 150622 165721 150678 166521 6 i_dout0[22]
port 15 nsew signal input
rlabel metal3 s 163577 126488 164377 126608 6 i_dout0[23]
port 16 nsew signal input
rlabel metal2 s 153474 165721 153530 166521 6 i_dout0[24]
port 17 nsew signal input
rlabel metal2 s 156326 165721 156382 166521 6 i_dout0[25]
port 18 nsew signal input
rlabel metal3 s 163577 136144 164377 136264 6 i_dout0[26]
port 19 nsew signal input
rlabel metal3 s 163577 148248 164377 148368 6 i_dout0[27]
port 20 nsew signal input
rlabel metal2 s 158902 0 158958 800 6 i_dout0[28]
port 21 nsew signal input
rlabel metal3 s 163577 157904 164377 158024 6 i_dout0[29]
port 22 nsew signal input
rlabel metal3 s 163577 20272 164377 20392 6 i_dout0[2]
port 23 nsew signal input
rlabel metal2 s 161846 0 161902 800 6 i_dout0[30]
port 24 nsew signal input
rlabel metal2 s 163870 165721 163926 166521 6 i_dout0[31]
port 25 nsew signal input
rlabel metal2 s 121090 165721 121146 166521 6 i_dout0[3]
port 26 nsew signal input
rlabel metal3 s 0 27616 800 27736 6 i_dout0[4]
port 27 nsew signal input
rlabel metal2 s 125874 165721 125930 166521 6 i_dout0[5]
port 28 nsew signal input
rlabel metal2 s 125230 0 125286 800 6 i_dout0[6]
port 29 nsew signal input
rlabel metal3 s 163577 56584 164377 56704 6 i_dout0[7]
port 30 nsew signal input
rlabel metal3 s 163577 63792 164377 63912 6 i_dout0[8]
port 31 nsew signal input
rlabel metal3 s 163577 66104 164377 66224 6 i_dout0[9]
port 32 nsew signal input
rlabel metal2 s 111338 0 111394 800 6 i_dout0_1[0]
port 33 nsew signal input
rlabel metal3 s 163577 73448 164377 73568 6 i_dout0_1[10]
port 34 nsew signal input
rlabel metal3 s 163577 80656 164377 80776 6 i_dout0_1[11]
port 35 nsew signal input
rlabel metal3 s 163577 87864 164377 87984 6 i_dout0_1[12]
port 36 nsew signal input
rlabel metal2 s 138110 0 138166 800 6 i_dout0_1[13]
port 37 nsew signal input
rlabel metal3 s 163577 92760 164377 92880 6 i_dout0_1[14]
port 38 nsew signal input
rlabel metal2 s 140042 0 140098 800 6 i_dout0_1[15]
port 39 nsew signal input
rlabel metal3 s 0 91808 800 91928 6 i_dout0_1[16]
port 40 nsew signal input
rlabel metal3 s 0 100648 800 100768 6 i_dout0_1[17]
port 41 nsew signal input
rlabel metal2 s 146758 165721 146814 166521 6 i_dout0_1[18]
port 42 nsew signal input
rlabel metal3 s 0 118056 800 118176 6 i_dout0_1[19]
port 43 nsew signal input
rlabel metal3 s 163577 10616 164377 10736 6 i_dout0_1[1]
port 44 nsew signal input
rlabel metal3 s 163577 114384 164377 114504 6 i_dout0_1[20]
port 45 nsew signal input
rlabel metal2 s 148966 0 149022 800 6 i_dout0_1[21]
port 46 nsew signal input
rlabel metal3 s 163577 119280 164377 119400 6 i_dout0_1[22]
port 47 nsew signal input
rlabel metal2 s 151542 165721 151598 166521 6 i_dout0_1[23]
port 48 nsew signal input
rlabel metal3 s 0 144440 800 144560 6 i_dout0_1[24]
port 49 nsew signal input
rlabel metal2 s 154394 165721 154450 166521 6 i_dout0_1[25]
port 50 nsew signal input
rlabel metal2 s 156878 0 156934 800 6 i_dout0_1[26]
port 51 nsew signal input
rlabel metal3 s 163577 145800 164377 145920 6 i_dout0_1[27]
port 52 nsew signal input
rlabel metal3 s 163577 153008 164377 153128 6 i_dout0_1[28]
port 53 nsew signal input
rlabel metal3 s 0 156136 800 156256 6 i_dout0_1[29]
port 54 nsew signal input
rlabel metal2 s 118238 165721 118294 166521 6 i_dout0_1[2]
port 55 nsew signal input
rlabel metal3 s 163577 160216 164377 160336 6 i_dout0_1[30]
port 56 nsew signal input
rlabel metal2 s 162950 165721 163006 166521 6 i_dout0_1[31]
port 57 nsew signal input
rlabel metal3 s 0 15920 800 16040 6 i_dout0_1[3]
port 58 nsew signal input
rlabel metal2 s 122286 0 122342 800 6 i_dout0_1[4]
port 59 nsew signal input
rlabel metal3 s 0 39312 800 39432 6 i_dout0_1[5]
port 60 nsew signal input
rlabel metal3 s 0 45160 800 45280 6 i_dout0_1[6]
port 61 nsew signal input
rlabel metal2 s 127162 0 127218 800 6 i_dout0_1[7]
port 62 nsew signal input
rlabel metal3 s 0 56856 800 56976 6 i_dout0_1[8]
port 63 nsew signal input
rlabel metal3 s 0 65560 800 65680 6 i_dout0_1[9]
port 64 nsew signal input
rlabel metal2 s 111614 165721 111670 166521 6 i_dout1[0]
port 65 nsew signal input
rlabel metal3 s 163577 78208 164377 78328 6 i_dout1[10]
port 66 nsew signal input
rlabel metal2 s 138202 165721 138258 166521 6 i_dout1[11]
port 67 nsew signal input
rlabel metal3 s 0 77256 800 77376 6 i_dout1[12]
port 68 nsew signal input
rlabel metal3 s 0 85960 800 86080 6 i_dout1[13]
port 69 nsew signal input
rlabel metal3 s 163577 95072 164377 95192 6 i_dout1[14]
port 70 nsew signal input
rlabel metal2 s 142066 0 142122 800 6 i_dout1[15]
port 71 nsew signal input
rlabel metal3 s 0 94800 800 94920 6 i_dout1[16]
port 72 nsew signal input
rlabel metal3 s 163577 104728 164377 104848 6 i_dout1[17]
port 73 nsew signal input
rlabel metal3 s 0 109352 800 109472 6 i_dout1[18]
port 74 nsew signal input
rlabel metal2 s 145010 0 145066 800 6 i_dout1[19]
port 75 nsew signal input
rlabel metal3 s 163577 15512 164377 15632 6 i_dout1[1]
port 76 nsew signal input
rlabel metal3 s 0 123904 800 124024 6 i_dout1[20]
port 77 nsew signal input
rlabel metal3 s 163577 116832 164377 116952 6 i_dout1[21]
port 78 nsew signal input
rlabel metal3 s 163577 121592 164377 121712 6 i_dout1[22]
port 79 nsew signal input
rlabel metal2 s 152002 0 152058 800 6 i_dout1[23]
port 80 nsew signal input
rlabel metal3 s 163577 128936 164377 129056 6 i_dout1[24]
port 81 nsew signal input
rlabel metal2 s 154946 0 155002 800 6 i_dout1[25]
port 82 nsew signal input
rlabel metal3 s 163577 138592 164377 138712 6 i_dout1[26]
port 83 nsew signal input
rlabel metal3 s 163577 150560 164377 150680 6 i_dout1[27]
port 84 nsew signal input
rlabel metal2 s 159178 165721 159234 166521 6 i_dout1[28]
port 85 nsew signal input
rlabel metal2 s 161018 165721 161074 166521 6 i_dout1[29]
port 86 nsew signal input
rlabel metal3 s 163577 22720 164377 22840 6 i_dout1[2]
port 87 nsew signal input
rlabel metal2 s 162030 165721 162086 166521 6 i_dout1[30]
port 88 nsew signal input
rlabel metal3 s 0 164840 800 164960 6 i_dout1[31]
port 89 nsew signal input
rlabel metal3 s 0 21768 800 21888 6 i_dout1[3]
port 90 nsew signal input
rlabel metal3 s 0 30472 800 30592 6 i_dout1[4]
port 91 nsew signal input
rlabel metal3 s 163577 42032 164377 42152 6 i_dout1[5]
port 92 nsew signal input
rlabel metal2 s 126242 0 126298 800 6 i_dout1[6]
port 93 nsew signal input
rlabel metal3 s 163577 58896 164377 59016 6 i_dout1[7]
port 94 nsew signal input
rlabel metal3 s 0 59712 800 59832 6 i_dout1[8]
port 95 nsew signal input
rlabel metal3 s 163577 68552 164377 68672 6 i_dout1[9]
port 96 nsew signal input
rlabel metal3 s 163577 1096 164377 1216 6 i_dout1_1[0]
port 97 nsew signal input
rlabel metal2 s 137282 165721 137338 166521 6 i_dout1_1[10]
port 98 nsew signal input
rlabel metal3 s 0 71408 800 71528 6 i_dout1_1[11]
port 99 nsew signal input
rlabel metal2 s 136086 0 136142 800 6 i_dout1_1[12]
port 100 nsew signal input
rlabel metal3 s 0 83104 800 83224 6 i_dout1_1[13]
port 101 nsew signal input
rlabel metal2 s 141054 165721 141110 166521 6 i_dout1_1[14]
port 102 nsew signal input
rlabel metal2 s 143906 165721 143962 166521 6 i_dout1_1[15]
port 103 nsew signal input
rlabel metal2 s 144918 165721 144974 166521 6 i_dout1_1[16]
port 104 nsew signal input
rlabel metal3 s 163577 102416 164377 102536 6 i_dout1_1[17]
port 105 nsew signal input
rlabel metal3 s 0 106496 800 106616 6 i_dout1_1[18]
port 106 nsew signal input
rlabel metal3 s 163577 112072 164377 112192 6 i_dout1_1[19]
port 107 nsew signal input
rlabel metal2 s 115386 165721 115442 166521 6 i_dout1_1[1]
port 108 nsew signal input
rlabel metal3 s 0 121048 800 121168 6 i_dout1_1[20]
port 109 nsew signal input
rlabel metal3 s 0 126896 800 127016 6 i_dout1_1[21]
port 110 nsew signal input
rlabel metal2 s 150990 0 151046 800 6 i_dout1_1[22]
port 111 nsew signal input
rlabel metal2 s 152462 165721 152518 166521 6 i_dout1_1[23]
port 112 nsew signal input
rlabel metal2 s 152922 0 152978 800 6 i_dout1_1[24]
port 113 nsew signal input
rlabel metal2 s 155314 165721 155370 166521 6 i_dout1_1[25]
port 114 nsew signal input
rlabel metal2 s 157890 0 157946 800 6 i_dout1_1[26]
port 115 nsew signal input
rlabel metal2 s 157246 165721 157302 166521 6 i_dout1_1[27]
port 116 nsew signal input
rlabel metal3 s 0 150288 800 150408 6 i_dout1_1[28]
port 117 nsew signal input
rlabel metal3 s 163577 155456 164377 155576 6 i_dout1_1[29]
port 118 nsew signal input
rlabel metal2 s 118330 0 118386 800 6 i_dout1_1[2]
port 119 nsew signal input
rlabel metal2 s 160834 0 160890 800 6 i_dout1_1[30]
port 120 nsew signal input
rlabel metal3 s 163577 165112 164377 165232 6 i_dout1_1[31]
port 121 nsew signal input
rlabel metal3 s 0 18776 800 18896 6 i_dout1_1[3]
port 122 nsew signal input
rlabel metal3 s 163577 34824 164377 34944 6 i_dout1_1[4]
port 123 nsew signal input
rlabel metal2 s 124218 0 124274 800 6 i_dout1_1[5]
port 124 nsew signal input
rlabel metal2 s 130658 165721 130714 166521 6 i_dout1_1[6]
port 125 nsew signal input
rlabel metal2 s 131578 165721 131634 166521 6 i_dout1_1[7]
port 126 nsew signal input
rlabel metal2 s 134430 165721 134486 166521 6 i_dout1_1[8]
port 127 nsew signal input
rlabel metal2 s 133142 0 133198 800 6 i_dout1_1[9]
port 128 nsew signal input
rlabel metal2 s 478 165721 534 166521 6 io_in[0]
port 129 nsew signal input
rlabel metal2 s 28906 165721 28962 166521 6 io_in[10]
port 130 nsew signal input
rlabel metal2 s 31758 165721 31814 166521 6 io_in[11]
port 131 nsew signal input
rlabel metal2 s 34610 165721 34666 166521 6 io_in[12]
port 132 nsew signal input
rlabel metal2 s 37462 165721 37518 166521 6 io_in[13]
port 133 nsew signal input
rlabel metal2 s 40314 165721 40370 166521 6 io_in[14]
port 134 nsew signal input
rlabel metal2 s 43166 165721 43222 166521 6 io_in[15]
port 135 nsew signal input
rlabel metal2 s 46018 165721 46074 166521 6 io_in[16]
port 136 nsew signal input
rlabel metal2 s 48870 165721 48926 166521 6 io_in[17]
port 137 nsew signal input
rlabel metal2 s 51722 165721 51778 166521 6 io_in[18]
port 138 nsew signal input
rlabel metal2 s 54574 165721 54630 166521 6 io_in[19]
port 139 nsew signal input
rlabel metal2 s 3238 165721 3294 166521 6 io_in[1]
port 140 nsew signal input
rlabel metal2 s 57426 165721 57482 166521 6 io_in[20]
port 141 nsew signal input
rlabel metal2 s 60278 165721 60334 166521 6 io_in[21]
port 142 nsew signal input
rlabel metal2 s 63130 165721 63186 166521 6 io_in[22]
port 143 nsew signal input
rlabel metal2 s 65982 165721 66038 166521 6 io_in[23]
port 144 nsew signal input
rlabel metal2 s 68834 165721 68890 166521 6 io_in[24]
port 145 nsew signal input
rlabel metal2 s 71686 165721 71742 166521 6 io_in[25]
port 146 nsew signal input
rlabel metal2 s 74538 165721 74594 166521 6 io_in[26]
port 147 nsew signal input
rlabel metal2 s 77390 165721 77446 166521 6 io_in[27]
port 148 nsew signal input
rlabel metal2 s 80242 165721 80298 166521 6 io_in[28]
port 149 nsew signal input
rlabel metal2 s 83094 165721 83150 166521 6 io_in[29]
port 150 nsew signal input
rlabel metal2 s 6090 165721 6146 166521 6 io_in[2]
port 151 nsew signal input
rlabel metal2 s 85946 165721 86002 166521 6 io_in[30]
port 152 nsew signal input
rlabel metal2 s 88798 165721 88854 166521 6 io_in[31]
port 153 nsew signal input
rlabel metal2 s 91650 165721 91706 166521 6 io_in[32]
port 154 nsew signal input
rlabel metal2 s 94502 165721 94558 166521 6 io_in[33]
port 155 nsew signal input
rlabel metal2 s 97354 165721 97410 166521 6 io_in[34]
port 156 nsew signal input
rlabel metal2 s 100206 165721 100262 166521 6 io_in[35]
port 157 nsew signal input
rlabel metal2 s 103058 165721 103114 166521 6 io_in[36]
port 158 nsew signal input
rlabel metal2 s 105910 165721 105966 166521 6 io_in[37]
port 159 nsew signal input
rlabel metal2 s 8942 165721 8998 166521 6 io_in[3]
port 160 nsew signal input
rlabel metal2 s 11794 165721 11850 166521 6 io_in[4]
port 161 nsew signal input
rlabel metal2 s 14646 165721 14702 166521 6 io_in[5]
port 162 nsew signal input
rlabel metal2 s 17498 165721 17554 166521 6 io_in[6]
port 163 nsew signal input
rlabel metal2 s 20350 165721 20406 166521 6 io_in[7]
port 164 nsew signal input
rlabel metal2 s 23202 165721 23258 166521 6 io_in[8]
port 165 nsew signal input
rlabel metal2 s 26054 165721 26110 166521 6 io_in[9]
port 166 nsew signal input
rlabel metal2 s 1398 165721 1454 166521 6 io_oeb[0]
port 167 nsew signal output
rlabel metal2 s 29918 165721 29974 166521 6 io_oeb[10]
port 168 nsew signal output
rlabel metal2 s 32770 165721 32826 166521 6 io_oeb[11]
port 169 nsew signal output
rlabel metal2 s 35622 165721 35678 166521 6 io_oeb[12]
port 170 nsew signal output
rlabel metal2 s 38474 165721 38530 166521 6 io_oeb[13]
port 171 nsew signal output
rlabel metal2 s 41326 165721 41382 166521 6 io_oeb[14]
port 172 nsew signal output
rlabel metal2 s 44178 165721 44234 166521 6 io_oeb[15]
port 173 nsew signal output
rlabel metal2 s 47030 165721 47086 166521 6 io_oeb[16]
port 174 nsew signal output
rlabel metal2 s 49882 165721 49938 166521 6 io_oeb[17]
port 175 nsew signal output
rlabel metal2 s 52734 165721 52790 166521 6 io_oeb[18]
port 176 nsew signal output
rlabel metal2 s 55586 165721 55642 166521 6 io_oeb[19]
port 177 nsew signal output
rlabel metal2 s 4250 165721 4306 166521 6 io_oeb[1]
port 178 nsew signal output
rlabel metal2 s 58438 165721 58494 166521 6 io_oeb[20]
port 179 nsew signal output
rlabel metal2 s 61290 165721 61346 166521 6 io_oeb[21]
port 180 nsew signal output
rlabel metal2 s 64142 165721 64198 166521 6 io_oeb[22]
port 181 nsew signal output
rlabel metal2 s 66994 165721 67050 166521 6 io_oeb[23]
port 182 nsew signal output
rlabel metal2 s 69846 165721 69902 166521 6 io_oeb[24]
port 183 nsew signal output
rlabel metal2 s 72698 165721 72754 166521 6 io_oeb[25]
port 184 nsew signal output
rlabel metal2 s 75550 165721 75606 166521 6 io_oeb[26]
port 185 nsew signal output
rlabel metal2 s 78402 165721 78458 166521 6 io_oeb[27]
port 186 nsew signal output
rlabel metal2 s 81254 165721 81310 166521 6 io_oeb[28]
port 187 nsew signal output
rlabel metal2 s 84014 165721 84070 166521 6 io_oeb[29]
port 188 nsew signal output
rlabel metal2 s 7102 165721 7158 166521 6 io_oeb[2]
port 189 nsew signal output
rlabel metal2 s 86866 165721 86922 166521 6 io_oeb[30]
port 190 nsew signal output
rlabel metal2 s 89718 165721 89774 166521 6 io_oeb[31]
port 191 nsew signal output
rlabel metal2 s 92570 165721 92626 166521 6 io_oeb[32]
port 192 nsew signal output
rlabel metal2 s 95422 165721 95478 166521 6 io_oeb[33]
port 193 nsew signal output
rlabel metal2 s 98274 165721 98330 166521 6 io_oeb[34]
port 194 nsew signal output
rlabel metal2 s 101126 165721 101182 166521 6 io_oeb[35]
port 195 nsew signal output
rlabel metal2 s 103978 165721 104034 166521 6 io_oeb[36]
port 196 nsew signal output
rlabel metal2 s 106830 165721 106886 166521 6 io_oeb[37]
port 197 nsew signal output
rlabel metal2 s 9954 165721 10010 166521 6 io_oeb[3]
port 198 nsew signal output
rlabel metal2 s 12806 165721 12862 166521 6 io_oeb[4]
port 199 nsew signal output
rlabel metal2 s 15658 165721 15714 166521 6 io_oeb[5]
port 200 nsew signal output
rlabel metal2 s 18510 165721 18566 166521 6 io_oeb[6]
port 201 nsew signal output
rlabel metal2 s 21362 165721 21418 166521 6 io_oeb[7]
port 202 nsew signal output
rlabel metal2 s 24214 165721 24270 166521 6 io_oeb[8]
port 203 nsew signal output
rlabel metal2 s 27066 165721 27122 166521 6 io_oeb[9]
port 204 nsew signal output
rlabel metal2 s 2318 165721 2374 166521 6 io_out[0]
port 205 nsew signal output
rlabel metal2 s 30838 165721 30894 166521 6 io_out[10]
port 206 nsew signal output
rlabel metal2 s 33690 165721 33746 166521 6 io_out[11]
port 207 nsew signal output
rlabel metal2 s 36542 165721 36598 166521 6 io_out[12]
port 208 nsew signal output
rlabel metal2 s 39394 165721 39450 166521 6 io_out[13]
port 209 nsew signal output
rlabel metal2 s 42246 165721 42302 166521 6 io_out[14]
port 210 nsew signal output
rlabel metal2 s 45098 165721 45154 166521 6 io_out[15]
port 211 nsew signal output
rlabel metal2 s 47950 165721 48006 166521 6 io_out[16]
port 212 nsew signal output
rlabel metal2 s 50802 165721 50858 166521 6 io_out[17]
port 213 nsew signal output
rlabel metal2 s 53654 165721 53710 166521 6 io_out[18]
port 214 nsew signal output
rlabel metal2 s 56506 165721 56562 166521 6 io_out[19]
port 215 nsew signal output
rlabel metal2 s 5170 165721 5226 166521 6 io_out[1]
port 216 nsew signal output
rlabel metal2 s 59358 165721 59414 166521 6 io_out[20]
port 217 nsew signal output
rlabel metal2 s 62210 165721 62266 166521 6 io_out[21]
port 218 nsew signal output
rlabel metal2 s 65062 165721 65118 166521 6 io_out[22]
port 219 nsew signal output
rlabel metal2 s 67914 165721 67970 166521 6 io_out[23]
port 220 nsew signal output
rlabel metal2 s 70766 165721 70822 166521 6 io_out[24]
port 221 nsew signal output
rlabel metal2 s 73618 165721 73674 166521 6 io_out[25]
port 222 nsew signal output
rlabel metal2 s 76470 165721 76526 166521 6 io_out[26]
port 223 nsew signal output
rlabel metal2 s 79322 165721 79378 166521 6 io_out[27]
port 224 nsew signal output
rlabel metal2 s 82174 165721 82230 166521 6 io_out[28]
port 225 nsew signal output
rlabel metal2 s 85026 165721 85082 166521 6 io_out[29]
port 226 nsew signal output
rlabel metal2 s 8022 165721 8078 166521 6 io_out[2]
port 227 nsew signal output
rlabel metal2 s 87878 165721 87934 166521 6 io_out[30]
port 228 nsew signal output
rlabel metal2 s 90730 165721 90786 166521 6 io_out[31]
port 229 nsew signal output
rlabel metal2 s 93582 165721 93638 166521 6 io_out[32]
port 230 nsew signal output
rlabel metal2 s 96434 165721 96490 166521 6 io_out[33]
port 231 nsew signal output
rlabel metal2 s 99286 165721 99342 166521 6 io_out[34]
port 232 nsew signal output
rlabel metal2 s 102138 165721 102194 166521 6 io_out[35]
port 233 nsew signal output
rlabel metal2 s 104990 165721 105046 166521 6 io_out[36]
port 234 nsew signal output
rlabel metal2 s 107842 165721 107898 166521 6 io_out[37]
port 235 nsew signal output
rlabel metal2 s 10874 165721 10930 166521 6 io_out[3]
port 236 nsew signal output
rlabel metal2 s 13726 165721 13782 166521 6 io_out[4]
port 237 nsew signal output
rlabel metal2 s 16578 165721 16634 166521 6 io_out[5]
port 238 nsew signal output
rlabel metal2 s 19430 165721 19486 166521 6 io_out[6]
port 239 nsew signal output
rlabel metal2 s 22282 165721 22338 166521 6 io_out[7]
port 240 nsew signal output
rlabel metal2 s 25134 165721 25190 166521 6 io_out[8]
port 241 nsew signal output
rlabel metal2 s 27986 165721 28042 166521 6 io_out[9]
port 242 nsew signal output
rlabel metal2 s 105450 0 105506 800 6 irq[0]
port 243 nsew signal output
rlabel metal2 s 106370 0 106426 800 6 irq[1]
port 244 nsew signal output
rlabel metal2 s 107382 0 107438 800 6 irq[2]
port 245 nsew signal output
rlabel metal2 s 112534 165721 112590 166521 6 o_addr1[0]
port 246 nsew signal output
rlabel metal3 s 163577 17960 164377 18080 6 o_addr1[1]
port 247 nsew signal output
rlabel metal3 s 0 10072 800 10192 6 o_addr1[2]
port 248 nsew signal output
rlabel metal2 s 123022 165721 123078 166521 6 o_addr1[3]
port 249 nsew signal output
rlabel metal3 s 0 33464 800 33584 6 o_addr1[4]
port 250 nsew signal output
rlabel metal2 s 127806 165721 127862 166521 6 o_addr1[5]
port 251 nsew signal output
rlabel metal3 s 0 48016 800 48136 6 o_addr1[6]
port 252 nsew signal output
rlabel metal2 s 132498 165721 132554 166521 6 o_addr1[7]
port 253 nsew signal output
rlabel metal2 s 131118 0 131174 800 6 o_addr1[8]
port 254 nsew signal output
rlabel metal3 s 163577 3408 164377 3528 6 o_addr1_1[0]
port 255 nsew signal output
rlabel metal2 s 116398 165721 116454 166521 6 o_addr1_1[1]
port 256 nsew signal output
rlabel metal3 s 0 7080 800 7200 6 o_addr1_1[2]
port 257 nsew signal output
rlabel metal2 s 122102 165721 122158 166521 6 o_addr1_1[3]
port 258 nsew signal output
rlabel metal2 s 124954 165721 125010 166521 6 o_addr1_1[4]
port 259 nsew signal output
rlabel metal2 s 126794 165721 126850 166521 6 o_addr1_1[5]
port 260 nsew signal output
rlabel metal3 s 163577 46928 164377 47048 6 o_addr1_1[6]
port 261 nsew signal output
rlabel metal2 s 128174 0 128230 800 6 o_addr1_1[7]
port 262 nsew signal output
rlabel metal2 s 130198 0 130254 800 6 o_addr1_1[8]
port 263 nsew signal output
rlabel metal2 s 108394 0 108450 800 6 o_csb0
port 264 nsew signal output
rlabel metal2 s 108762 165721 108818 166521 6 o_csb0_1
port 265 nsew signal output
rlabel metal2 s 109682 165721 109738 166521 6 o_csb1
port 266 nsew signal output
rlabel metal2 s 109406 0 109462 800 6 o_csb1_1
port 267 nsew signal output
rlabel metal3 s 163577 5856 164377 5976 6 o_din0[0]
port 268 nsew signal output
rlabel metal2 s 135166 0 135222 800 6 o_din0[10]
port 269 nsew signal output
rlabel metal3 s 163577 85416 164377 85536 6 o_din0[11]
port 270 nsew signal output
rlabel metal3 s 0 80112 800 80232 6 o_din0[12]
port 271 nsew signal output
rlabel metal2 s 139122 0 139178 800 6 o_din0[13]
port 272 nsew signal output
rlabel metal2 s 142986 165721 143042 166521 6 o_din0[14]
port 273 nsew signal output
rlabel metal3 s 163577 97520 164377 97640 6 o_din0[15]
port 274 nsew signal output
rlabel metal2 s 143998 0 144054 800 6 o_din0[16]
port 275 nsew signal output
rlabel metal3 s 163577 107176 164377 107296 6 o_din0[17]
port 276 nsew signal output
rlabel metal3 s 0 115200 800 115320 6 o_din0[18]
port 277 nsew signal output
rlabel metal2 s 148690 165721 148746 166521 6 o_din0[19]
port 278 nsew signal output
rlabel metal2 s 115294 0 115350 800 6 o_din0[1]
port 279 nsew signal output
rlabel metal2 s 147954 0 148010 800 6 o_din0[20]
port 280 nsew signal output
rlabel metal3 s 0 132744 800 132864 6 o_din0[21]
port 281 nsew signal output
rlabel metal3 s 163577 124040 164377 124160 6 o_din0[22]
port 282 nsew signal output
rlabel metal3 s 0 141448 800 141568 6 o_din0[23]
port 283 nsew signal output
rlabel metal3 s 163577 131248 164377 131368 6 o_din0[24]
port 284 nsew signal output
rlabel metal3 s 163577 133696 164377 133816 6 o_din0[25]
port 285 nsew signal output
rlabel metal3 s 163577 143352 164377 143472 6 o_din0[26]
port 286 nsew signal output
rlabel metal3 s 0 147296 800 147416 6 o_din0[27]
port 287 nsew signal output
rlabel metal2 s 160098 165721 160154 166521 6 o_din0[28]
port 288 nsew signal output
rlabel metal3 s 0 158992 800 159112 6 o_din0[29]
port 289 nsew signal output
rlabel metal3 s 0 12928 800 13048 6 o_din0[2]
port 290 nsew signal output
rlabel metal3 s 0 161984 800 162104 6 o_din0[30]
port 291 nsew signal output
rlabel metal2 s 163870 0 163926 800 6 o_din0[31]
port 292 nsew signal output
rlabel metal3 s 163577 29928 164377 30048 6 o_din0[3]
port 293 nsew signal output
rlabel metal3 s 0 36320 800 36440 6 o_din0[4]
port 294 nsew signal output
rlabel metal2 s 129646 165721 129702 166521 6 o_din0[5]
port 295 nsew signal output
rlabel metal3 s 163577 51688 164377 51808 6 o_din0[6]
port 296 nsew signal output
rlabel metal3 s 0 53864 800 53984 6 o_din0[7]
port 297 nsew signal output
rlabel metal2 s 132130 0 132186 800 6 o_din0[8]
port 298 nsew signal output
rlabel metal3 s 163577 71000 164377 71120 6 o_din0[9]
port 299 nsew signal output
rlabel metal2 s 113546 165721 113602 166521 6 o_din0_1[0]
port 300 nsew signal output
rlabel metal2 s 134154 0 134210 800 6 o_din0_1[10]
port 301 nsew signal output
rlabel metal3 s 0 74264 800 74384 6 o_din0_1[11]
port 302 nsew signal output
rlabel metal2 s 139214 165721 139270 166521 6 o_din0_1[12]
port 303 nsew signal output
rlabel metal2 s 140134 165721 140190 166521 6 o_din0_1[13]
port 304 nsew signal output
rlabel metal3 s 0 88952 800 89072 6 o_din0_1[14]
port 305 nsew signal output
rlabel metal2 s 143078 0 143134 800 6 o_din0_1[15]
port 306 nsew signal output
rlabel metal3 s 0 97656 800 97776 6 o_din0_1[16]
port 307 nsew signal output
rlabel metal3 s 0 103504 800 103624 6 o_din0_1[17]
port 308 nsew signal output
rlabel metal3 s 0 112344 800 112464 6 o_din0_1[18]
port 309 nsew signal output
rlabel metal2 s 146022 0 146078 800 6 o_din0_1[19]
port 310 nsew signal output
rlabel metal2 s 114282 0 114338 800 6 o_din0_1[1]
port 311 nsew signal output
rlabel metal2 s 147034 0 147090 800 6 o_din0_1[20]
port 312 nsew signal output
rlabel metal3 s 0 129752 800 129872 6 o_din0_1[21]
port 313 nsew signal output
rlabel metal3 s 0 135600 800 135720 6 o_din0_1[22]
port 314 nsew signal output
rlabel metal3 s 0 138592 800 138712 6 o_din0_1[23]
port 315 nsew signal output
rlabel metal2 s 153934 0 153990 800 6 o_din0_1[24]
port 316 nsew signal output
rlabel metal2 s 155958 0 156014 800 6 o_din0_1[25]
port 317 nsew signal output
rlabel metal3 s 163577 140904 164377 141024 6 o_din0_1[26]
port 318 nsew signal output
rlabel metal2 s 158166 165721 158222 166521 6 o_din0_1[27]
port 319 nsew signal output
rlabel metal3 s 0 153144 800 153264 6 o_din0_1[28]
port 320 nsew signal output
rlabel metal2 s 159914 0 159970 800 6 o_din0_1[29]
port 321 nsew signal output
rlabel metal2 s 119250 0 119306 800 6 o_din0_1[2]
port 322 nsew signal output
rlabel metal3 s 163577 162664 164377 162784 6 o_din0_1[30]
port 323 nsew signal output
rlabel metal2 s 162858 0 162914 800 6 o_din0_1[31]
port 324 nsew signal output
rlabel metal3 s 0 24624 800 24744 6 o_din0_1[3]
port 325 nsew signal output
rlabel metal3 s 163577 37272 164377 37392 6 o_din0_1[4]
port 326 nsew signal output
rlabel metal2 s 128726 165721 128782 166521 6 o_din0_1[5]
port 327 nsew signal output
rlabel metal3 s 163577 49240 164377 49360 6 o_din0_1[6]
port 328 nsew signal output
rlabel metal2 s 129186 0 129242 800 6 o_din0_1[7]
port 329 nsew signal output
rlabel metal2 s 135350 165721 135406 166521 6 o_din0_1[8]
port 330 nsew signal output
rlabel metal3 s 0 68416 800 68536 6 o_din0_1[9]
port 331 nsew signal output
rlabel metal2 s 114466 165721 114522 166521 6 o_waddr0[0]
port 332 nsew signal output
rlabel metal2 s 117318 165721 117374 166521 6 o_waddr0[1]
port 333 nsew signal output
rlabel metal3 s 163577 25168 164377 25288 6 o_waddr0[2]
port 334 nsew signal output
rlabel metal2 s 120262 0 120318 800 6 o_waddr0[3]
port 335 nsew signal output
rlabel metal2 s 123206 0 123262 800 6 o_waddr0[4]
port 336 nsew signal output
rlabel metal3 s 163577 44480 164377 44600 6 o_waddr0[5]
port 337 nsew signal output
rlabel metal3 s 0 51008 800 51128 6 o_waddr0[6]
port 338 nsew signal output
rlabel metal3 s 163577 61344 164377 61464 6 o_waddr0[7]
port 339 nsew signal output
rlabel metal3 s 0 62568 800 62688 6 o_waddr0[8]
port 340 nsew signal output
rlabel metal3 s 163577 8304 164377 8424 6 o_waddr0_1[0]
port 341 nsew signal output
rlabel metal3 s 0 4224 800 4344 6 o_waddr0_1[1]
port 342 nsew signal output
rlabel metal2 s 119250 165721 119306 166521 6 o_waddr0_1[2]
port 343 nsew signal output
rlabel metal3 s 163577 32376 164377 32496 6 o_waddr0_1[3]
port 344 nsew signal output
rlabel metal3 s 163577 39584 164377 39704 6 o_waddr0_1[4]
port 345 nsew signal output
rlabel metal3 s 0 42168 800 42288 6 o_waddr0_1[5]
port 346 nsew signal output
rlabel metal3 s 163577 54136 164377 54256 6 o_waddr0_1[6]
port 347 nsew signal output
rlabel metal2 s 133510 165721 133566 166521 6 o_waddr0_1[7]
port 348 nsew signal output
rlabel metal2 s 136362 165721 136418 166521 6 o_waddr0_1[8]
port 349 nsew signal output
rlabel metal2 s 110326 0 110382 800 6 o_web0
port 350 nsew signal output
rlabel metal3 s 0 1368 800 1488 6 o_web0_1
port 351 nsew signal output
rlabel metal2 s 112350 0 112406 800 6 o_wmask0[0]
port 352 nsew signal output
rlabel metal2 s 117318 0 117374 800 6 o_wmask0[1]
port 353 nsew signal output
rlabel metal2 s 120170 165721 120226 166521 6 o_wmask0[2]
port 354 nsew signal output
rlabel metal2 s 121274 0 121330 800 6 o_wmask0[3]
port 355 nsew signal output
rlabel metal2 s 113362 0 113418 800 6 o_wmask0_1[0]
port 356 nsew signal output
rlabel metal2 s 116306 0 116362 800 6 o_wmask0_1[1]
port 357 nsew signal output
rlabel metal3 s 163577 27616 164377 27736 6 o_wmask0_1[2]
port 358 nsew signal output
rlabel metal2 s 123942 165721 123998 166521 6 o_wmask0_1[3]
port 359 nsew signal output
rlabel metal4 s 4208 2128 4528 164336 6 vccd1
port 360 nsew power input
rlabel metal4 s 34928 2128 35248 164336 6 vccd1
port 360 nsew power input
rlabel metal4 s 65648 2128 65968 164336 6 vccd1
port 360 nsew power input
rlabel metal4 s 96368 2128 96688 164336 6 vccd1
port 360 nsew power input
rlabel metal4 s 127088 2128 127408 164336 6 vccd1
port 360 nsew power input
rlabel metal4 s 157808 2128 158128 164336 6 vccd1
port 360 nsew power input
rlabel metal4 s 19568 2128 19888 164336 6 vssd1
port 361 nsew ground input
rlabel metal4 s 50288 2128 50608 164336 6 vssd1
port 361 nsew ground input
rlabel metal4 s 81008 2128 81328 164336 6 vssd1
port 361 nsew ground input
rlabel metal4 s 111728 2128 112048 164336 6 vssd1
port 361 nsew ground input
rlabel metal4 s 142448 2128 142768 164336 6 vssd1
port 361 nsew ground input
rlabel metal2 s 478 0 534 800 6 wb_clk_i
port 362 nsew signal input
rlabel metal2 s 1398 0 1454 800 6 wb_rst_i
port 363 nsew signal input
rlabel metal2 s 2410 0 2466 800 6 wbs_ack_o
port 364 nsew signal output
rlabel metal2 s 6366 0 6422 800 6 wbs_adr_i[0]
port 365 nsew signal input
rlabel metal2 s 40038 0 40094 800 6 wbs_adr_i[10]
port 366 nsew signal input
rlabel metal2 s 42982 0 43038 800 6 wbs_adr_i[11]
port 367 nsew signal input
rlabel metal2 s 46018 0 46074 800 6 wbs_adr_i[12]
port 368 nsew signal input
rlabel metal2 s 48962 0 49018 800 6 wbs_adr_i[13]
port 369 nsew signal input
rlabel metal2 s 51906 0 51962 800 6 wbs_adr_i[14]
port 370 nsew signal input
rlabel metal2 s 54942 0 54998 800 6 wbs_adr_i[15]
port 371 nsew signal input
rlabel metal2 s 57886 0 57942 800 6 wbs_adr_i[16]
port 372 nsew signal input
rlabel metal2 s 60830 0 60886 800 6 wbs_adr_i[17]
port 373 nsew signal input
rlabel metal2 s 63774 0 63830 800 6 wbs_adr_i[18]
port 374 nsew signal input
rlabel metal2 s 66810 0 66866 800 6 wbs_adr_i[19]
port 375 nsew signal input
rlabel metal2 s 10322 0 10378 800 6 wbs_adr_i[1]
port 376 nsew signal input
rlabel metal2 s 69754 0 69810 800 6 wbs_adr_i[20]
port 377 nsew signal input
rlabel metal2 s 72698 0 72754 800 6 wbs_adr_i[21]
port 378 nsew signal input
rlabel metal2 s 75734 0 75790 800 6 wbs_adr_i[22]
port 379 nsew signal input
rlabel metal2 s 78678 0 78734 800 6 wbs_adr_i[23]
port 380 nsew signal input
rlabel metal2 s 81622 0 81678 800 6 wbs_adr_i[24]
port 381 nsew signal input
rlabel metal2 s 84658 0 84714 800 6 wbs_adr_i[25]
port 382 nsew signal input
rlabel metal2 s 87602 0 87658 800 6 wbs_adr_i[26]
port 383 nsew signal input
rlabel metal2 s 90546 0 90602 800 6 wbs_adr_i[27]
port 384 nsew signal input
rlabel metal2 s 93490 0 93546 800 6 wbs_adr_i[28]
port 385 nsew signal input
rlabel metal2 s 96526 0 96582 800 6 wbs_adr_i[29]
port 386 nsew signal input
rlabel metal2 s 14278 0 14334 800 6 wbs_adr_i[2]
port 387 nsew signal input
rlabel metal2 s 99470 0 99526 800 6 wbs_adr_i[30]
port 388 nsew signal input
rlabel metal2 s 102414 0 102470 800 6 wbs_adr_i[31]
port 389 nsew signal input
rlabel metal2 s 18234 0 18290 800 6 wbs_adr_i[3]
port 390 nsew signal input
rlabel metal2 s 22190 0 22246 800 6 wbs_adr_i[4]
port 391 nsew signal input
rlabel metal2 s 25226 0 25282 800 6 wbs_adr_i[5]
port 392 nsew signal input
rlabel metal2 s 28170 0 28226 800 6 wbs_adr_i[6]
port 393 nsew signal input
rlabel metal2 s 31114 0 31170 800 6 wbs_adr_i[7]
port 394 nsew signal input
rlabel metal2 s 34150 0 34206 800 6 wbs_adr_i[8]
port 395 nsew signal input
rlabel metal2 s 37094 0 37150 800 6 wbs_adr_i[9]
port 396 nsew signal input
rlabel metal2 s 3422 0 3478 800 6 wbs_cyc_i
port 397 nsew signal input
rlabel metal2 s 7378 0 7434 800 6 wbs_dat_i[0]
port 398 nsew signal input
rlabel metal2 s 41050 0 41106 800 6 wbs_dat_i[10]
port 399 nsew signal input
rlabel metal2 s 43994 0 44050 800 6 wbs_dat_i[11]
port 400 nsew signal input
rlabel metal2 s 46938 0 46994 800 6 wbs_dat_i[12]
port 401 nsew signal input
rlabel metal2 s 49974 0 50030 800 6 wbs_dat_i[13]
port 402 nsew signal input
rlabel metal2 s 52918 0 52974 800 6 wbs_dat_i[14]
port 403 nsew signal input
rlabel metal2 s 55862 0 55918 800 6 wbs_dat_i[15]
port 404 nsew signal input
rlabel metal2 s 58898 0 58954 800 6 wbs_dat_i[16]
port 405 nsew signal input
rlabel metal2 s 61842 0 61898 800 6 wbs_dat_i[17]
port 406 nsew signal input
rlabel metal2 s 64786 0 64842 800 6 wbs_dat_i[18]
port 407 nsew signal input
rlabel metal2 s 67822 0 67878 800 6 wbs_dat_i[19]
port 408 nsew signal input
rlabel metal2 s 11334 0 11390 800 6 wbs_dat_i[1]
port 409 nsew signal input
rlabel metal2 s 70766 0 70822 800 6 wbs_dat_i[20]
port 410 nsew signal input
rlabel metal2 s 73710 0 73766 800 6 wbs_dat_i[21]
port 411 nsew signal input
rlabel metal2 s 76654 0 76710 800 6 wbs_dat_i[22]
port 412 nsew signal input
rlabel metal2 s 79690 0 79746 800 6 wbs_dat_i[23]
port 413 nsew signal input
rlabel metal2 s 82634 0 82690 800 6 wbs_dat_i[24]
port 414 nsew signal input
rlabel metal2 s 85578 0 85634 800 6 wbs_dat_i[25]
port 415 nsew signal input
rlabel metal2 s 88614 0 88670 800 6 wbs_dat_i[26]
port 416 nsew signal input
rlabel metal2 s 91558 0 91614 800 6 wbs_dat_i[27]
port 417 nsew signal input
rlabel metal2 s 94502 0 94558 800 6 wbs_dat_i[28]
port 418 nsew signal input
rlabel metal2 s 97446 0 97502 800 6 wbs_dat_i[29]
port 419 nsew signal input
rlabel metal2 s 15290 0 15346 800 6 wbs_dat_i[2]
port 420 nsew signal input
rlabel metal2 s 100482 0 100538 800 6 wbs_dat_i[30]
port 421 nsew signal input
rlabel metal2 s 103426 0 103482 800 6 wbs_dat_i[31]
port 422 nsew signal input
rlabel metal2 s 19246 0 19302 800 6 wbs_dat_i[3]
port 423 nsew signal input
rlabel metal2 s 23202 0 23258 800 6 wbs_dat_i[4]
port 424 nsew signal input
rlabel metal2 s 26146 0 26202 800 6 wbs_dat_i[5]
port 425 nsew signal input
rlabel metal2 s 29182 0 29238 800 6 wbs_dat_i[6]
port 426 nsew signal input
rlabel metal2 s 32126 0 32182 800 6 wbs_dat_i[7]
port 427 nsew signal input
rlabel metal2 s 35070 0 35126 800 6 wbs_dat_i[8]
port 428 nsew signal input
rlabel metal2 s 38106 0 38162 800 6 wbs_dat_i[9]
port 429 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 wbs_dat_o[0]
port 430 nsew signal output
rlabel metal2 s 42062 0 42118 800 6 wbs_dat_o[10]
port 431 nsew signal output
rlabel metal2 s 45006 0 45062 800 6 wbs_dat_o[11]
port 432 nsew signal output
rlabel metal2 s 47950 0 48006 800 6 wbs_dat_o[12]
port 433 nsew signal output
rlabel metal2 s 50986 0 51042 800 6 wbs_dat_o[13]
port 434 nsew signal output
rlabel metal2 s 53930 0 53986 800 6 wbs_dat_o[14]
port 435 nsew signal output
rlabel metal2 s 56874 0 56930 800 6 wbs_dat_o[15]
port 436 nsew signal output
rlabel metal2 s 59818 0 59874 800 6 wbs_dat_o[16]
port 437 nsew signal output
rlabel metal2 s 62854 0 62910 800 6 wbs_dat_o[17]
port 438 nsew signal output
rlabel metal2 s 65798 0 65854 800 6 wbs_dat_o[18]
port 439 nsew signal output
rlabel metal2 s 68742 0 68798 800 6 wbs_dat_o[19]
port 440 nsew signal output
rlabel metal2 s 12346 0 12402 800 6 wbs_dat_o[1]
port 441 nsew signal output
rlabel metal2 s 71778 0 71834 800 6 wbs_dat_o[20]
port 442 nsew signal output
rlabel metal2 s 74722 0 74778 800 6 wbs_dat_o[21]
port 443 nsew signal output
rlabel metal2 s 77666 0 77722 800 6 wbs_dat_o[22]
port 444 nsew signal output
rlabel metal2 s 80610 0 80666 800 6 wbs_dat_o[23]
port 445 nsew signal output
rlabel metal2 s 83646 0 83702 800 6 wbs_dat_o[24]
port 446 nsew signal output
rlabel metal2 s 86590 0 86646 800 6 wbs_dat_o[25]
port 447 nsew signal output
rlabel metal2 s 89534 0 89590 800 6 wbs_dat_o[26]
port 448 nsew signal output
rlabel metal2 s 92570 0 92626 800 6 wbs_dat_o[27]
port 449 nsew signal output
rlabel metal2 s 95514 0 95570 800 6 wbs_dat_o[28]
port 450 nsew signal output
rlabel metal2 s 98458 0 98514 800 6 wbs_dat_o[29]
port 451 nsew signal output
rlabel metal2 s 16302 0 16358 800 6 wbs_dat_o[2]
port 452 nsew signal output
rlabel metal2 s 101494 0 101550 800 6 wbs_dat_o[30]
port 453 nsew signal output
rlabel metal2 s 104438 0 104494 800 6 wbs_dat_o[31]
port 454 nsew signal output
rlabel metal2 s 20258 0 20314 800 6 wbs_dat_o[3]
port 455 nsew signal output
rlabel metal2 s 24214 0 24270 800 6 wbs_dat_o[4]
port 456 nsew signal output
rlabel metal2 s 27158 0 27214 800 6 wbs_dat_o[5]
port 457 nsew signal output
rlabel metal2 s 30102 0 30158 800 6 wbs_dat_o[6]
port 458 nsew signal output
rlabel metal2 s 33138 0 33194 800 6 wbs_dat_o[7]
port 459 nsew signal output
rlabel metal2 s 36082 0 36138 800 6 wbs_dat_o[8]
port 460 nsew signal output
rlabel metal2 s 39026 0 39082 800 6 wbs_dat_o[9]
port 461 nsew signal output
rlabel metal2 s 9310 0 9366 800 6 wbs_sel_i[0]
port 462 nsew signal input
rlabel metal2 s 13266 0 13322 800 6 wbs_sel_i[1]
port 463 nsew signal input
rlabel metal2 s 17314 0 17370 800 6 wbs_sel_i[2]
port 464 nsew signal input
rlabel metal2 s 21270 0 21326 800 6 wbs_sel_i[3]
port 465 nsew signal input
rlabel metal2 s 4434 0 4490 800 6 wbs_stb_i
port 466 nsew signal input
rlabel metal2 s 5354 0 5410 800 6 wbs_we_i
port 467 nsew signal input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 164377 166521
string LEFview TRUE
string GDS_FILE /local/caravel_user_project/openlane/user_proj/runs/user_proj/results/magic/user_proj.gds
string GDS_END 81744398
string GDS_START 1419336
<< end >>

