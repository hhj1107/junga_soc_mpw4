magic
tech sky130A
magscale 1 2
timestamp 1640633896
<< obsli1 >>
rect 1104 2159 164191 164305
<< obsm1 >>
rect 106 8 164298 164336
<< metal2 >>
rect 478 165864 534 166664
rect 1398 165864 1454 166664
rect 2318 165864 2374 166664
rect 3238 165864 3294 166664
rect 4158 165864 4214 166664
rect 5170 165864 5226 166664
rect 6090 165864 6146 166664
rect 7010 165864 7066 166664
rect 7930 165864 7986 166664
rect 8850 165864 8906 166664
rect 9862 165864 9918 166664
rect 10782 165864 10838 166664
rect 11702 165864 11758 166664
rect 12622 165864 12678 166664
rect 13634 165864 13690 166664
rect 14554 165864 14610 166664
rect 15474 165864 15530 166664
rect 16394 165864 16450 166664
rect 17314 165864 17370 166664
rect 18326 165864 18382 166664
rect 19246 165864 19302 166664
rect 20166 165864 20222 166664
rect 21086 165864 21142 166664
rect 22006 165864 22062 166664
rect 23018 165864 23074 166664
rect 23938 165864 23994 166664
rect 24858 165864 24914 166664
rect 25778 165864 25834 166664
rect 26790 165864 26846 166664
rect 27710 165864 27766 166664
rect 28630 165864 28686 166664
rect 29550 165864 29606 166664
rect 30470 165864 30526 166664
rect 31482 165864 31538 166664
rect 32402 165864 32458 166664
rect 33322 165864 33378 166664
rect 34242 165864 34298 166664
rect 35254 165864 35310 166664
rect 36174 165864 36230 166664
rect 37094 165864 37150 166664
rect 38014 165864 38070 166664
rect 38934 165864 38990 166664
rect 39946 165864 40002 166664
rect 40866 165864 40922 166664
rect 41786 165864 41842 166664
rect 42706 165864 42762 166664
rect 43626 165864 43682 166664
rect 44638 165864 44694 166664
rect 45558 165864 45614 166664
rect 46478 165864 46534 166664
rect 47398 165864 47454 166664
rect 48410 165864 48466 166664
rect 49330 165864 49386 166664
rect 50250 165864 50306 166664
rect 51170 165864 51226 166664
rect 52090 165864 52146 166664
rect 53102 165864 53158 166664
rect 54022 165864 54078 166664
rect 54942 165864 54998 166664
rect 55862 165864 55918 166664
rect 56874 165864 56930 166664
rect 57794 165864 57850 166664
rect 58714 165864 58770 166664
rect 59634 165864 59690 166664
rect 60554 165864 60610 166664
rect 61566 165864 61622 166664
rect 62486 165864 62542 166664
rect 63406 165864 63462 166664
rect 64326 165864 64382 166664
rect 65246 165864 65302 166664
rect 66258 165864 66314 166664
rect 67178 165864 67234 166664
rect 68098 165864 68154 166664
rect 69018 165864 69074 166664
rect 70030 165864 70086 166664
rect 70950 165864 71006 166664
rect 71870 165864 71926 166664
rect 72790 165864 72846 166664
rect 73710 165864 73766 166664
rect 74722 165864 74778 166664
rect 75642 165864 75698 166664
rect 76562 165864 76618 166664
rect 77482 165864 77538 166664
rect 78494 165864 78550 166664
rect 79414 165864 79470 166664
rect 80334 165864 80390 166664
rect 81254 165864 81310 166664
rect 82174 165864 82230 166664
rect 83186 165864 83242 166664
rect 84106 165864 84162 166664
rect 85026 165864 85082 166664
rect 85946 165864 86002 166664
rect 86866 165864 86922 166664
rect 87878 165864 87934 166664
rect 88798 165864 88854 166664
rect 89718 165864 89774 166664
rect 90638 165864 90694 166664
rect 91650 165864 91706 166664
rect 92570 165864 92626 166664
rect 93490 165864 93546 166664
rect 94410 165864 94466 166664
rect 95330 165864 95386 166664
rect 96342 165864 96398 166664
rect 97262 165864 97318 166664
rect 98182 165864 98238 166664
rect 99102 165864 99158 166664
rect 100114 165864 100170 166664
rect 101034 165864 101090 166664
rect 101954 165864 102010 166664
rect 102874 165864 102930 166664
rect 103794 165864 103850 166664
rect 104806 165864 104862 166664
rect 105726 165864 105782 166664
rect 106646 165864 106702 166664
rect 107566 165864 107622 166664
rect 108486 165864 108542 166664
rect 109498 165864 109554 166664
rect 110418 165864 110474 166664
rect 111338 165864 111394 166664
rect 112258 165864 112314 166664
rect 113270 165864 113326 166664
rect 114190 165864 114246 166664
rect 115110 165864 115166 166664
rect 116030 165864 116086 166664
rect 116950 165864 117006 166664
rect 117962 165864 118018 166664
rect 118882 165864 118938 166664
rect 119802 165864 119858 166664
rect 120722 165864 120778 166664
rect 121734 165864 121790 166664
rect 122654 165864 122710 166664
rect 123574 165864 123630 166664
rect 124494 165864 124550 166664
rect 125414 165864 125470 166664
rect 126426 165864 126482 166664
rect 127346 165864 127402 166664
rect 128266 165864 128322 166664
rect 129186 165864 129242 166664
rect 130106 165864 130162 166664
rect 131118 165864 131174 166664
rect 132038 165864 132094 166664
rect 132958 165864 133014 166664
rect 133878 165864 133934 166664
rect 134890 165864 134946 166664
rect 135810 165864 135866 166664
rect 136730 165864 136786 166664
rect 137650 165864 137706 166664
rect 138570 165864 138626 166664
rect 139582 165864 139638 166664
rect 140502 165864 140558 166664
rect 141422 165864 141478 166664
rect 142342 165864 142398 166664
rect 143354 165864 143410 166664
rect 144274 165864 144330 166664
rect 145194 165864 145250 166664
rect 146114 165864 146170 166664
rect 147034 165864 147090 166664
rect 148046 165864 148102 166664
rect 148966 165864 149022 166664
rect 149886 165864 149942 166664
rect 150806 165864 150862 166664
rect 151726 165864 151782 166664
rect 152738 165864 152794 166664
rect 153658 165864 153714 166664
rect 154578 165864 154634 166664
rect 155498 165864 155554 166664
rect 156510 165864 156566 166664
rect 157430 165864 157486 166664
rect 158350 165864 158406 166664
rect 159270 165864 159326 166664
rect 160190 165864 160246 166664
rect 161202 165864 161258 166664
rect 162122 165864 162178 166664
rect 163042 165864 163098 166664
rect 163962 165864 164018 166664
rect 478 0 534 800
rect 1398 0 1454 800
rect 2318 0 2374 800
rect 3330 0 3386 800
rect 4250 0 4306 800
rect 5262 0 5318 800
rect 6182 0 6238 800
rect 7194 0 7250 800
rect 8114 0 8170 800
rect 9126 0 9182 800
rect 10046 0 10102 800
rect 11058 0 11114 800
rect 11978 0 12034 800
rect 12898 0 12954 800
rect 13910 0 13966 800
rect 14830 0 14886 800
rect 15842 0 15898 800
rect 16762 0 16818 800
rect 17774 0 17830 800
rect 18694 0 18750 800
rect 19706 0 19762 800
rect 20626 0 20682 800
rect 21638 0 21694 800
rect 22558 0 22614 800
rect 23478 0 23534 800
rect 24490 0 24546 800
rect 25410 0 25466 800
rect 26422 0 26478 800
rect 27342 0 27398 800
rect 28354 0 28410 800
rect 29274 0 29330 800
rect 30286 0 30342 800
rect 31206 0 31262 800
rect 32218 0 32274 800
rect 33138 0 33194 800
rect 34058 0 34114 800
rect 35070 0 35126 800
rect 35990 0 36046 800
rect 37002 0 37058 800
rect 37922 0 37978 800
rect 38934 0 38990 800
rect 39854 0 39910 800
rect 40866 0 40922 800
rect 41786 0 41842 800
rect 42798 0 42854 800
rect 43718 0 43774 800
rect 44638 0 44694 800
rect 45650 0 45706 800
rect 46570 0 46626 800
rect 47582 0 47638 800
rect 48502 0 48558 800
rect 49514 0 49570 800
rect 50434 0 50490 800
rect 51446 0 51502 800
rect 52366 0 52422 800
rect 53378 0 53434 800
rect 54298 0 54354 800
rect 55310 0 55366 800
rect 56230 0 56286 800
rect 57150 0 57206 800
rect 58162 0 58218 800
rect 59082 0 59138 800
rect 60094 0 60150 800
rect 61014 0 61070 800
rect 62026 0 62082 800
rect 62946 0 63002 800
rect 63958 0 64014 800
rect 64878 0 64934 800
rect 65890 0 65946 800
rect 66810 0 66866 800
rect 67730 0 67786 800
rect 68742 0 68798 800
rect 69662 0 69718 800
rect 70674 0 70730 800
rect 71594 0 71650 800
rect 72606 0 72662 800
rect 73526 0 73582 800
rect 74538 0 74594 800
rect 75458 0 75514 800
rect 76470 0 76526 800
rect 77390 0 77446 800
rect 78310 0 78366 800
rect 79322 0 79378 800
rect 80242 0 80298 800
rect 81254 0 81310 800
rect 82174 0 82230 800
rect 83186 0 83242 800
rect 84106 0 84162 800
rect 85118 0 85174 800
rect 86038 0 86094 800
rect 87050 0 87106 800
rect 87970 0 88026 800
rect 88890 0 88946 800
rect 89902 0 89958 800
rect 90822 0 90878 800
rect 91834 0 91890 800
rect 92754 0 92810 800
rect 93766 0 93822 800
rect 94686 0 94742 800
rect 95698 0 95754 800
rect 96618 0 96674 800
rect 97630 0 97686 800
rect 98550 0 98606 800
rect 99470 0 99526 800
rect 100482 0 100538 800
rect 101402 0 101458 800
rect 102414 0 102470 800
rect 103334 0 103390 800
rect 104346 0 104402 800
rect 105266 0 105322 800
rect 106278 0 106334 800
rect 107198 0 107254 800
rect 108210 0 108266 800
rect 109130 0 109186 800
rect 110142 0 110198 800
rect 111062 0 111118 800
rect 111982 0 112038 800
rect 112994 0 113050 800
rect 113914 0 113970 800
rect 114926 0 114982 800
rect 115846 0 115902 800
rect 116858 0 116914 800
rect 117778 0 117834 800
rect 118790 0 118846 800
rect 119710 0 119766 800
rect 120722 0 120778 800
rect 121642 0 121698 800
rect 122562 0 122618 800
rect 123574 0 123630 800
rect 124494 0 124550 800
rect 125506 0 125562 800
rect 126426 0 126482 800
rect 127438 0 127494 800
rect 128358 0 128414 800
rect 129370 0 129426 800
rect 130290 0 130346 800
rect 131302 0 131358 800
rect 132222 0 132278 800
rect 133142 0 133198 800
rect 134154 0 134210 800
rect 135074 0 135130 800
rect 136086 0 136142 800
rect 137006 0 137062 800
rect 138018 0 138074 800
rect 138938 0 138994 800
rect 139950 0 140006 800
rect 140870 0 140926 800
rect 141882 0 141938 800
rect 142802 0 142858 800
rect 143722 0 143778 800
rect 144734 0 144790 800
rect 145654 0 145710 800
rect 146666 0 146722 800
rect 147586 0 147642 800
rect 148598 0 148654 800
rect 149518 0 149574 800
rect 150530 0 150586 800
rect 151450 0 151506 800
rect 152462 0 152518 800
rect 153382 0 153438 800
rect 154302 0 154358 800
rect 155314 0 155370 800
rect 156234 0 156290 800
rect 157246 0 157302 800
rect 158166 0 158222 800
rect 159178 0 159234 800
rect 160098 0 160154 800
rect 161110 0 161166 800
rect 162030 0 162086 800
rect 163042 0 163098 800
rect 163962 0 164018 800
<< obsm2 >>
rect 18 165808 422 166002
rect 590 165808 1342 166002
rect 1510 165808 2262 166002
rect 2430 165808 3182 166002
rect 3350 165808 4102 166002
rect 4270 165808 5114 166002
rect 5282 165808 6034 166002
rect 6202 165808 6954 166002
rect 7122 165808 7874 166002
rect 8042 165808 8794 166002
rect 8962 165808 9806 166002
rect 9974 165808 10726 166002
rect 10894 165808 11646 166002
rect 11814 165808 12566 166002
rect 12734 165808 13578 166002
rect 13746 165808 14498 166002
rect 14666 165808 15418 166002
rect 15586 165808 16338 166002
rect 16506 165808 17258 166002
rect 17426 165808 18270 166002
rect 18438 165808 19190 166002
rect 19358 165808 20110 166002
rect 20278 165808 21030 166002
rect 21198 165808 21950 166002
rect 22118 165808 22962 166002
rect 23130 165808 23882 166002
rect 24050 165808 24802 166002
rect 24970 165808 25722 166002
rect 25890 165808 26734 166002
rect 26902 165808 27654 166002
rect 27822 165808 28574 166002
rect 28742 165808 29494 166002
rect 29662 165808 30414 166002
rect 30582 165808 31426 166002
rect 31594 165808 32346 166002
rect 32514 165808 33266 166002
rect 33434 165808 34186 166002
rect 34354 165808 35198 166002
rect 35366 165808 36118 166002
rect 36286 165808 37038 166002
rect 37206 165808 37958 166002
rect 38126 165808 38878 166002
rect 39046 165808 39890 166002
rect 40058 165808 40810 166002
rect 40978 165808 41730 166002
rect 41898 165808 42650 166002
rect 42818 165808 43570 166002
rect 43738 165808 44582 166002
rect 44750 165808 45502 166002
rect 45670 165808 46422 166002
rect 46590 165808 47342 166002
rect 47510 165808 48354 166002
rect 48522 165808 49274 166002
rect 49442 165808 50194 166002
rect 50362 165808 51114 166002
rect 51282 165808 52034 166002
rect 52202 165808 53046 166002
rect 53214 165808 53966 166002
rect 54134 165808 54886 166002
rect 55054 165808 55806 166002
rect 55974 165808 56818 166002
rect 56986 165808 57738 166002
rect 57906 165808 58658 166002
rect 58826 165808 59578 166002
rect 59746 165808 60498 166002
rect 60666 165808 61510 166002
rect 61678 165808 62430 166002
rect 62598 165808 63350 166002
rect 63518 165808 64270 166002
rect 64438 165808 65190 166002
rect 65358 165808 66202 166002
rect 66370 165808 67122 166002
rect 67290 165808 68042 166002
rect 68210 165808 68962 166002
rect 69130 165808 69974 166002
rect 70142 165808 70894 166002
rect 71062 165808 71814 166002
rect 71982 165808 72734 166002
rect 72902 165808 73654 166002
rect 73822 165808 74666 166002
rect 74834 165808 75586 166002
rect 75754 165808 76506 166002
rect 76674 165808 77426 166002
rect 77594 165808 78438 166002
rect 78606 165808 79358 166002
rect 79526 165808 80278 166002
rect 80446 165808 81198 166002
rect 81366 165808 82118 166002
rect 82286 165808 83130 166002
rect 83298 165808 84050 166002
rect 84218 165808 84970 166002
rect 85138 165808 85890 166002
rect 86058 165808 86810 166002
rect 86978 165808 87822 166002
rect 87990 165808 88742 166002
rect 88910 165808 89662 166002
rect 89830 165808 90582 166002
rect 90750 165808 91594 166002
rect 91762 165808 92514 166002
rect 92682 165808 93434 166002
rect 93602 165808 94354 166002
rect 94522 165808 95274 166002
rect 95442 165808 96286 166002
rect 96454 165808 97206 166002
rect 97374 165808 98126 166002
rect 98294 165808 99046 166002
rect 99214 165808 100058 166002
rect 100226 165808 100978 166002
rect 101146 165808 101898 166002
rect 102066 165808 102818 166002
rect 102986 165808 103738 166002
rect 103906 165808 104750 166002
rect 104918 165808 105670 166002
rect 105838 165808 106590 166002
rect 106758 165808 107510 166002
rect 107678 165808 108430 166002
rect 108598 165808 109442 166002
rect 109610 165808 110362 166002
rect 110530 165808 111282 166002
rect 111450 165808 112202 166002
rect 112370 165808 113214 166002
rect 113382 165808 114134 166002
rect 114302 165808 115054 166002
rect 115222 165808 115974 166002
rect 116142 165808 116894 166002
rect 117062 165808 117906 166002
rect 118074 165808 118826 166002
rect 118994 165808 119746 166002
rect 119914 165808 120666 166002
rect 120834 165808 121678 166002
rect 121846 165808 122598 166002
rect 122766 165808 123518 166002
rect 123686 165808 124438 166002
rect 124606 165808 125358 166002
rect 125526 165808 126370 166002
rect 126538 165808 127290 166002
rect 127458 165808 128210 166002
rect 128378 165808 129130 166002
rect 129298 165808 130050 166002
rect 130218 165808 131062 166002
rect 131230 165808 131982 166002
rect 132150 165808 132902 166002
rect 133070 165808 133822 166002
rect 133990 165808 134834 166002
rect 135002 165808 135754 166002
rect 135922 165808 136674 166002
rect 136842 165808 137594 166002
rect 137762 165808 138514 166002
rect 138682 165808 139526 166002
rect 139694 165808 140446 166002
rect 140614 165808 141366 166002
rect 141534 165808 142286 166002
rect 142454 165808 143298 166002
rect 143466 165808 144218 166002
rect 144386 165808 145138 166002
rect 145306 165808 146058 166002
rect 146226 165808 146978 166002
rect 147146 165808 147990 166002
rect 148158 165808 148910 166002
rect 149078 165808 149830 166002
rect 149998 165808 150750 166002
rect 150918 165808 151670 166002
rect 151838 165808 152682 166002
rect 152850 165808 153602 166002
rect 153770 165808 154522 166002
rect 154690 165808 155442 166002
rect 155610 165808 156454 166002
rect 156622 165808 157374 166002
rect 157542 165808 158294 166002
rect 158462 165808 159214 166002
rect 159382 165808 160134 166002
rect 160302 165808 161146 166002
rect 161314 165808 162066 166002
rect 162234 165808 162986 166002
rect 163154 165808 163906 166002
rect 164074 165808 164294 166002
rect 18 856 164294 165808
rect 18 2 422 856
rect 590 2 1342 856
rect 1510 2 2262 856
rect 2430 2 3274 856
rect 3442 2 4194 856
rect 4362 2 5206 856
rect 5374 2 6126 856
rect 6294 2 7138 856
rect 7306 2 8058 856
rect 8226 2 9070 856
rect 9238 2 9990 856
rect 10158 2 11002 856
rect 11170 2 11922 856
rect 12090 2 12842 856
rect 13010 2 13854 856
rect 14022 2 14774 856
rect 14942 2 15786 856
rect 15954 2 16706 856
rect 16874 2 17718 856
rect 17886 2 18638 856
rect 18806 2 19650 856
rect 19818 2 20570 856
rect 20738 2 21582 856
rect 21750 2 22502 856
rect 22670 2 23422 856
rect 23590 2 24434 856
rect 24602 2 25354 856
rect 25522 2 26366 856
rect 26534 2 27286 856
rect 27454 2 28298 856
rect 28466 2 29218 856
rect 29386 2 30230 856
rect 30398 2 31150 856
rect 31318 2 32162 856
rect 32330 2 33082 856
rect 33250 2 34002 856
rect 34170 2 35014 856
rect 35182 2 35934 856
rect 36102 2 36946 856
rect 37114 2 37866 856
rect 38034 2 38878 856
rect 39046 2 39798 856
rect 39966 2 40810 856
rect 40978 2 41730 856
rect 41898 2 42742 856
rect 42910 2 43662 856
rect 43830 2 44582 856
rect 44750 2 45594 856
rect 45762 2 46514 856
rect 46682 2 47526 856
rect 47694 2 48446 856
rect 48614 2 49458 856
rect 49626 2 50378 856
rect 50546 2 51390 856
rect 51558 2 52310 856
rect 52478 2 53322 856
rect 53490 2 54242 856
rect 54410 2 55254 856
rect 55422 2 56174 856
rect 56342 2 57094 856
rect 57262 2 58106 856
rect 58274 2 59026 856
rect 59194 2 60038 856
rect 60206 2 60958 856
rect 61126 2 61970 856
rect 62138 2 62890 856
rect 63058 2 63902 856
rect 64070 2 64822 856
rect 64990 2 65834 856
rect 66002 2 66754 856
rect 66922 2 67674 856
rect 67842 2 68686 856
rect 68854 2 69606 856
rect 69774 2 70618 856
rect 70786 2 71538 856
rect 71706 2 72550 856
rect 72718 2 73470 856
rect 73638 2 74482 856
rect 74650 2 75402 856
rect 75570 2 76414 856
rect 76582 2 77334 856
rect 77502 2 78254 856
rect 78422 2 79266 856
rect 79434 2 80186 856
rect 80354 2 81198 856
rect 81366 2 82118 856
rect 82286 2 83130 856
rect 83298 2 84050 856
rect 84218 2 85062 856
rect 85230 2 85982 856
rect 86150 2 86994 856
rect 87162 2 87914 856
rect 88082 2 88834 856
rect 89002 2 89846 856
rect 90014 2 90766 856
rect 90934 2 91778 856
rect 91946 2 92698 856
rect 92866 2 93710 856
rect 93878 2 94630 856
rect 94798 2 95642 856
rect 95810 2 96562 856
rect 96730 2 97574 856
rect 97742 2 98494 856
rect 98662 2 99414 856
rect 99582 2 100426 856
rect 100594 2 101346 856
rect 101514 2 102358 856
rect 102526 2 103278 856
rect 103446 2 104290 856
rect 104458 2 105210 856
rect 105378 2 106222 856
rect 106390 2 107142 856
rect 107310 2 108154 856
rect 108322 2 109074 856
rect 109242 2 110086 856
rect 110254 2 111006 856
rect 111174 2 111926 856
rect 112094 2 112938 856
rect 113106 2 113858 856
rect 114026 2 114870 856
rect 115038 2 115790 856
rect 115958 2 116802 856
rect 116970 2 117722 856
rect 117890 2 118734 856
rect 118902 2 119654 856
rect 119822 2 120666 856
rect 120834 2 121586 856
rect 121754 2 122506 856
rect 122674 2 123518 856
rect 123686 2 124438 856
rect 124606 2 125450 856
rect 125618 2 126370 856
rect 126538 2 127382 856
rect 127550 2 128302 856
rect 128470 2 129314 856
rect 129482 2 130234 856
rect 130402 2 131246 856
rect 131414 2 132166 856
rect 132334 2 133086 856
rect 133254 2 134098 856
rect 134266 2 135018 856
rect 135186 2 136030 856
rect 136198 2 136950 856
rect 137118 2 137962 856
rect 138130 2 138882 856
rect 139050 2 139894 856
rect 140062 2 140814 856
rect 140982 2 141826 856
rect 141994 2 142746 856
rect 142914 2 143666 856
rect 143834 2 144678 856
rect 144846 2 145598 856
rect 145766 2 146610 856
rect 146778 2 147530 856
rect 147698 2 148542 856
rect 148710 2 149462 856
rect 149630 2 150474 856
rect 150642 2 151394 856
rect 151562 2 152406 856
rect 152574 2 153326 856
rect 153494 2 154246 856
rect 154414 2 155258 856
rect 155426 2 156178 856
rect 156346 2 157190 856
rect 157358 2 158110 856
rect 158278 2 159122 856
rect 159290 2 160042 856
rect 160210 2 161054 856
rect 161222 2 161974 856
rect 162142 2 162986 856
rect 163154 2 163906 856
rect 164074 2 164294 856
<< metal3 >>
rect 0 165112 800 165232
rect 163720 165112 164520 165232
rect 0 162392 800 162512
rect 163720 162256 164520 162376
rect 0 159536 800 159656
rect 163720 159400 164520 159520
rect 0 156816 800 156936
rect 163720 156544 164520 156664
rect 0 153960 800 154080
rect 163720 153824 164520 153944
rect 0 151240 800 151360
rect 163720 150968 164520 151088
rect 0 148520 800 148640
rect 163720 148112 164520 148232
rect 0 145664 800 145784
rect 163720 145256 164520 145376
rect 0 142944 800 143064
rect 163720 142536 164520 142656
rect 0 140088 800 140208
rect 163720 139680 164520 139800
rect 0 137368 800 137488
rect 163720 136824 164520 136944
rect 0 134648 800 134768
rect 163720 133968 164520 134088
rect 0 131792 800 131912
rect 163720 131248 164520 131368
rect 0 129072 800 129192
rect 163720 128392 164520 128512
rect 0 126216 800 126336
rect 163720 125536 164520 125656
rect 0 123496 800 123616
rect 163720 122680 164520 122800
rect 0 120640 800 120760
rect 163720 119960 164520 120080
rect 0 117920 800 118040
rect 163720 117104 164520 117224
rect 0 115200 800 115320
rect 163720 114248 164520 114368
rect 0 112344 800 112464
rect 163720 111392 164520 111512
rect 0 109624 800 109744
rect 163720 108536 164520 108656
rect 0 106768 800 106888
rect 163720 105816 164520 105936
rect 0 104048 800 104168
rect 163720 102960 164520 103080
rect 0 101328 800 101448
rect 163720 100104 164520 100224
rect 0 98472 800 98592
rect 163720 97248 164520 97368
rect 0 95752 800 95872
rect 163720 94528 164520 94648
rect 0 92896 800 93016
rect 163720 91672 164520 91792
rect 0 90176 800 90296
rect 163720 88816 164520 88936
rect 0 87320 800 87440
rect 163720 85960 164520 86080
rect 0 84600 800 84720
rect 163720 83240 164520 83360
rect 0 81880 800 82000
rect 163720 80384 164520 80504
rect 0 79024 800 79144
rect 163720 77528 164520 77648
rect 0 76304 800 76424
rect 163720 74672 164520 74792
rect 0 73448 800 73568
rect 163720 71952 164520 72072
rect 0 70728 800 70848
rect 163720 69096 164520 69216
rect 0 68008 800 68128
rect 163720 66240 164520 66360
rect 0 65152 800 65272
rect 163720 63384 164520 63504
rect 0 62432 800 62552
rect 163720 60664 164520 60784
rect 0 59576 800 59696
rect 163720 57808 164520 57928
rect 0 56856 800 56976
rect 163720 54952 164520 55072
rect 0 54000 800 54120
rect 163720 52096 164520 52216
rect 0 51280 800 51400
rect 163720 49240 164520 49360
rect 0 48560 800 48680
rect 163720 46520 164520 46640
rect 0 45704 800 45824
rect 163720 43664 164520 43784
rect 0 42984 800 43104
rect 163720 40808 164520 40928
rect 0 40128 800 40248
rect 163720 37952 164520 38072
rect 0 37408 800 37528
rect 163720 35232 164520 35352
rect 0 34688 800 34808
rect 163720 32376 164520 32496
rect 0 31832 800 31952
rect 163720 29520 164520 29640
rect 0 29112 800 29232
rect 163720 26664 164520 26784
rect 0 26256 800 26376
rect 163720 23944 164520 24064
rect 0 23536 800 23656
rect 163720 21088 164520 21208
rect 0 20680 800 20800
rect 163720 18232 164520 18352
rect 0 17960 800 18080
rect 0 15240 800 15360
rect 163720 15376 164520 15496
rect 163720 12656 164520 12776
rect 0 12384 800 12504
rect 0 9664 800 9784
rect 163720 9800 164520 9920
rect 0 6808 800 6928
rect 163720 6944 164520 7064
rect 0 4088 800 4208
rect 163720 4088 164520 4208
rect 0 1368 800 1488
rect 163720 1368 164520 1488
<< obsm3 >>
rect 13 162592 164299 164321
rect 880 162456 164299 162592
rect 880 162312 163640 162456
rect 13 162176 163640 162312
rect 13 159736 164299 162176
rect 880 159600 164299 159736
rect 880 159456 163640 159600
rect 13 159320 163640 159456
rect 13 157016 164299 159320
rect 880 156744 164299 157016
rect 880 156736 163640 156744
rect 13 156464 163640 156736
rect 13 154160 164299 156464
rect 880 154024 164299 154160
rect 880 153880 163640 154024
rect 13 153744 163640 153880
rect 13 151440 164299 153744
rect 880 151168 164299 151440
rect 880 151160 163640 151168
rect 13 150888 163640 151160
rect 13 148720 164299 150888
rect 880 148440 164299 148720
rect 13 148312 164299 148440
rect 13 148032 163640 148312
rect 13 145864 164299 148032
rect 880 145584 164299 145864
rect 13 145456 164299 145584
rect 13 145176 163640 145456
rect 13 143144 164299 145176
rect 880 142864 164299 143144
rect 13 142736 164299 142864
rect 13 142456 163640 142736
rect 13 140288 164299 142456
rect 880 140008 164299 140288
rect 13 139880 164299 140008
rect 13 139600 163640 139880
rect 13 137568 164299 139600
rect 880 137288 164299 137568
rect 13 137024 164299 137288
rect 13 136744 163640 137024
rect 13 134848 164299 136744
rect 880 134568 164299 134848
rect 13 134168 164299 134568
rect 13 133888 163640 134168
rect 13 131992 164299 133888
rect 880 131712 164299 131992
rect 13 131448 164299 131712
rect 13 131168 163640 131448
rect 13 129272 164299 131168
rect 880 128992 164299 129272
rect 13 128592 164299 128992
rect 13 128312 163640 128592
rect 13 126416 164299 128312
rect 880 126136 164299 126416
rect 13 125736 164299 126136
rect 13 125456 163640 125736
rect 13 123696 164299 125456
rect 880 123416 164299 123696
rect 13 122880 164299 123416
rect 13 122600 163640 122880
rect 13 120840 164299 122600
rect 880 120560 164299 120840
rect 13 120160 164299 120560
rect 13 119880 163640 120160
rect 13 118120 164299 119880
rect 880 117840 164299 118120
rect 13 117304 164299 117840
rect 13 117024 163640 117304
rect 13 115400 164299 117024
rect 880 115120 164299 115400
rect 13 114448 164299 115120
rect 13 114168 163640 114448
rect 13 112544 164299 114168
rect 880 112264 164299 112544
rect 13 111592 164299 112264
rect 13 111312 163640 111592
rect 13 109824 164299 111312
rect 880 109544 164299 109824
rect 13 108736 164299 109544
rect 13 108456 163640 108736
rect 13 106968 164299 108456
rect 880 106688 164299 106968
rect 13 106016 164299 106688
rect 13 105736 163640 106016
rect 13 104248 164299 105736
rect 880 103968 164299 104248
rect 13 103160 164299 103968
rect 13 102880 163640 103160
rect 13 101528 164299 102880
rect 880 101248 164299 101528
rect 13 100304 164299 101248
rect 13 100024 163640 100304
rect 13 98672 164299 100024
rect 880 98392 164299 98672
rect 13 97448 164299 98392
rect 13 97168 163640 97448
rect 13 95952 164299 97168
rect 880 95672 164299 95952
rect 13 94728 164299 95672
rect 13 94448 163640 94728
rect 13 93096 164299 94448
rect 880 92816 164299 93096
rect 13 91872 164299 92816
rect 13 91592 163640 91872
rect 13 90376 164299 91592
rect 880 90096 164299 90376
rect 13 89016 164299 90096
rect 13 88736 163640 89016
rect 13 87520 164299 88736
rect 880 87240 164299 87520
rect 13 86160 164299 87240
rect 13 85880 163640 86160
rect 13 84800 164299 85880
rect 880 84520 164299 84800
rect 13 83440 164299 84520
rect 13 83160 163640 83440
rect 13 82080 164299 83160
rect 880 81800 164299 82080
rect 13 80584 164299 81800
rect 13 80304 163640 80584
rect 13 79224 164299 80304
rect 880 78944 164299 79224
rect 13 77728 164299 78944
rect 13 77448 163640 77728
rect 13 76504 164299 77448
rect 880 76224 164299 76504
rect 13 74872 164299 76224
rect 13 74592 163640 74872
rect 13 73648 164299 74592
rect 880 73368 164299 73648
rect 13 72152 164299 73368
rect 13 71872 163640 72152
rect 13 70928 164299 71872
rect 880 70648 164299 70928
rect 13 69296 164299 70648
rect 13 69016 163640 69296
rect 13 68208 164299 69016
rect 880 67928 164299 68208
rect 13 66440 164299 67928
rect 13 66160 163640 66440
rect 13 65352 164299 66160
rect 880 65072 164299 65352
rect 13 63584 164299 65072
rect 13 63304 163640 63584
rect 13 62632 164299 63304
rect 880 62352 164299 62632
rect 13 60864 164299 62352
rect 13 60584 163640 60864
rect 13 59776 164299 60584
rect 880 59496 164299 59776
rect 13 58008 164299 59496
rect 13 57728 163640 58008
rect 13 57056 164299 57728
rect 880 56776 164299 57056
rect 13 55152 164299 56776
rect 13 54872 163640 55152
rect 13 54200 164299 54872
rect 880 53920 164299 54200
rect 13 52296 164299 53920
rect 13 52016 163640 52296
rect 13 51480 164299 52016
rect 880 51200 164299 51480
rect 13 49440 164299 51200
rect 13 49160 163640 49440
rect 13 48760 164299 49160
rect 880 48480 164299 48760
rect 13 46720 164299 48480
rect 13 46440 163640 46720
rect 13 45904 164299 46440
rect 880 45624 164299 45904
rect 13 43864 164299 45624
rect 13 43584 163640 43864
rect 13 43184 164299 43584
rect 880 42904 164299 43184
rect 13 41008 164299 42904
rect 13 40728 163640 41008
rect 13 40328 164299 40728
rect 880 40048 164299 40328
rect 13 38152 164299 40048
rect 13 37872 163640 38152
rect 13 37608 164299 37872
rect 880 37328 164299 37608
rect 13 35432 164299 37328
rect 13 35152 163640 35432
rect 13 34888 164299 35152
rect 880 34608 164299 34888
rect 13 32576 164299 34608
rect 13 32296 163640 32576
rect 13 32032 164299 32296
rect 880 31752 164299 32032
rect 13 29720 164299 31752
rect 13 29440 163640 29720
rect 13 29312 164299 29440
rect 880 29032 164299 29312
rect 13 26864 164299 29032
rect 13 26584 163640 26864
rect 13 26456 164299 26584
rect 880 26176 164299 26456
rect 13 24144 164299 26176
rect 13 23864 163640 24144
rect 13 23736 164299 23864
rect 880 23456 164299 23736
rect 13 21288 164299 23456
rect 13 21008 163640 21288
rect 13 20880 164299 21008
rect 880 20600 164299 20880
rect 13 18432 164299 20600
rect 13 18160 163640 18432
rect 880 18152 163640 18160
rect 880 17880 164299 18152
rect 13 15576 164299 17880
rect 13 15440 163640 15576
rect 880 15296 163640 15440
rect 880 15160 164299 15296
rect 13 12856 164299 15160
rect 13 12584 163640 12856
rect 880 12576 163640 12584
rect 880 12304 164299 12576
rect 13 10000 164299 12304
rect 13 9864 163640 10000
rect 880 9720 163640 9864
rect 880 9584 164299 9720
rect 13 7144 164299 9584
rect 13 7008 163640 7144
rect 880 6864 163640 7008
rect 880 6728 164299 6864
rect 13 4288 164299 6728
rect 880 4008 163640 4288
rect 13 1568 164299 4008
rect 880 1288 163640 1568
rect 13 35 164299 1288
<< metal4 >>
rect 4208 2128 4528 164336
rect 19568 2128 19888 164336
rect 34928 2128 35248 164336
rect 50288 2128 50608 164336
rect 65648 2128 65968 164336
rect 81008 2128 81328 164336
rect 96368 2128 96688 164336
rect 111728 2128 112048 164336
rect 127088 2128 127408 164336
rect 142448 2128 142768 164336
rect 157808 2128 158128 164336
<< obsm4 >>
rect 427 2048 4128 164117
rect 4608 2048 19488 164117
rect 19968 2048 34848 164117
rect 35328 2048 50208 164117
rect 50688 2048 65568 164117
rect 66048 2048 80928 164117
rect 81408 2048 96288 164117
rect 96768 2048 111648 164117
rect 112128 2048 127008 164117
rect 127488 2048 142368 164117
rect 142848 2048 147509 164117
rect 427 1259 147509 2048
<< labels >>
rlabel metal2 s 109130 0 109186 800 6 i_dout0[0]
port 1 nsew signal input
rlabel metal3 s 163720 83240 164520 83360 6 i_dout0[10]
port 2 nsew signal input
rlabel metal2 s 134154 0 134210 800 6 i_dout0[11]
port 3 nsew signal input
rlabel metal3 s 0 84600 800 84720 6 i_dout0[12]
port 4 nsew signal input
rlabel metal3 s 163720 97248 164520 97368 6 i_dout0[13]
port 5 nsew signal input
rlabel metal2 s 133878 165864 133934 166664 6 i_dout0[14]
port 6 nsew signal input
rlabel metal2 s 143722 0 143778 800 6 i_dout0[15]
port 7 nsew signal input
rlabel metal2 s 137650 165864 137706 166664 6 i_dout0[16]
port 8 nsew signal input
rlabel metal2 s 147586 0 147642 800 6 i_dout0[17]
port 9 nsew signal input
rlabel metal2 s 138570 165864 138626 166664 6 i_dout0[18]
port 10 nsew signal input
rlabel metal3 s 163720 125536 164520 125656 6 i_dout0[19]
port 11 nsew signal input
rlabel metal3 s 163720 15376 164520 15496 6 i_dout0[1]
port 12 nsew signal input
rlabel metal3 s 163720 128392 164520 128512 6 i_dout0[20]
port 13 nsew signal input
rlabel metal3 s 163720 133968 164520 134088 6 i_dout0[21]
port 14 nsew signal input
rlabel metal2 s 146114 165864 146170 166664 6 i_dout0[22]
port 15 nsew signal input
rlabel metal3 s 163720 139680 164520 139800 6 i_dout0[23]
port 16 nsew signal input
rlabel metal2 s 150806 165864 150862 166664 6 i_dout0[24]
port 17 nsew signal input
rlabel metal2 s 157246 0 157302 800 6 i_dout0[25]
port 18 nsew signal input
rlabel metal3 s 0 134648 800 134768 6 i_dout0[26]
port 19 nsew signal input
rlabel metal2 s 156510 165864 156566 166664 6 i_dout0[27]
port 20 nsew signal input
rlabel metal3 s 0 148520 800 148640 6 i_dout0[28]
port 21 nsew signal input
rlabel metal3 s 163720 159400 164520 159520 6 i_dout0[29]
port 22 nsew signal input
rlabel metal2 s 116858 0 116914 800 6 i_dout0[2]
port 23 nsew signal input
rlabel metal2 s 161202 165864 161258 166664 6 i_dout0[30]
port 24 nsew signal input
rlabel metal3 s 0 165112 800 165232 6 i_dout0[31]
port 25 nsew signal input
rlabel metal3 s 163720 37952 164520 38072 6 i_dout0[3]
port 26 nsew signal input
rlabel metal3 s 0 40128 800 40248 6 i_dout0[4]
port 27 nsew signal input
rlabel metal3 s 0 51280 800 51400 6 i_dout0[5]
port 28 nsew signal input
rlabel metal2 s 118882 165864 118938 166664 6 i_dout0[6]
port 29 nsew signal input
rlabel metal3 s 163720 63384 164520 63504 6 i_dout0[7]
port 30 nsew signal input
rlabel metal3 s 0 76304 800 76424 6 i_dout0[8]
port 31 nsew signal input
rlabel metal2 s 131302 0 131358 800 6 i_dout0[9]
port 32 nsew signal input
rlabel metal3 s 163720 4088 164520 4208 6 i_dout0_1[0]
port 33 nsew signal input
rlabel metal2 s 129186 165864 129242 166664 6 i_dout0_1[10]
port 34 nsew signal input
rlabel metal2 s 133142 0 133198 800 6 i_dout0_1[11]
port 35 nsew signal input
rlabel metal3 s 163720 91672 164520 91792 6 i_dout0_1[12]
port 36 nsew signal input
rlabel metal2 s 132958 165864 133014 166664 6 i_dout0_1[13]
port 37 nsew signal input
rlabel metal2 s 141882 0 141938 800 6 i_dout0_1[14]
port 38 nsew signal input
rlabel metal3 s 0 90176 800 90296 6 i_dout0_1[15]
port 39 nsew signal input
rlabel metal3 s 0 95752 800 95872 6 i_dout0_1[16]
port 40 nsew signal input
rlabel metal3 s 163720 114248 164520 114368 6 i_dout0_1[17]
port 41 nsew signal input
rlabel metal3 s 163720 117104 164520 117224 6 i_dout0_1[18]
port 42 nsew signal input
rlabel metal2 s 139582 165864 139638 166664 6 i_dout0_1[19]
port 43 nsew signal input
rlabel metal3 s 163720 12656 164520 12776 6 i_dout0_1[1]
port 44 nsew signal input
rlabel metal2 s 142342 165864 142398 166664 6 i_dout0_1[20]
port 45 nsew signal input
rlabel metal3 s 0 115200 800 115320 6 i_dout0_1[21]
port 46 nsew signal input
rlabel metal3 s 163720 136824 164520 136944 6 i_dout0_1[22]
port 47 nsew signal input
rlabel metal2 s 153382 0 153438 800 6 i_dout0_1[23]
port 48 nsew signal input
rlabel metal2 s 149886 165864 149942 166664 6 i_dout0_1[24]
port 49 nsew signal input
rlabel metal2 s 151726 165864 151782 166664 6 i_dout0_1[25]
port 50 nsew signal input
rlabel metal2 s 158166 0 158222 800 6 i_dout0_1[26]
port 51 nsew signal input
rlabel metal3 s 0 140088 800 140208 6 i_dout0_1[27]
port 52 nsew signal input
rlabel metal2 s 159270 165864 159326 166664 6 i_dout0_1[28]
port 53 nsew signal input
rlabel metal2 s 161110 0 161166 800 6 i_dout0_1[29]
port 54 nsew signal input
rlabel metal2 s 115846 0 115902 800 6 i_dout0_1[2]
port 55 nsew signal input
rlabel metal2 s 160190 165864 160246 166664 6 i_dout0_1[30]
port 56 nsew signal input
rlabel metal3 s 0 162392 800 162512 6 i_dout0_1[31]
port 57 nsew signal input
rlabel metal3 s 163720 35232 164520 35352 6 i_dout0_1[3]
port 58 nsew signal input
rlabel metal3 s 0 37408 800 37528 6 i_dout0_1[4]
port 59 nsew signal input
rlabel metal3 s 163720 49240 164520 49360 6 i_dout0_1[5]
port 60 nsew signal input
rlabel metal3 s 0 56856 800 56976 6 i_dout0_1[6]
port 61 nsew signal input
rlabel metal2 s 123574 165864 123630 166664 6 i_dout0_1[7]
port 62 nsew signal input
rlabel metal3 s 0 70728 800 70848 6 i_dout0_1[8]
port 63 nsew signal input
rlabel metal3 s 163720 77528 164520 77648 6 i_dout0_1[9]
port 64 nsew signal input
rlabel metal3 s 163720 9800 164520 9920 6 i_dout1[0]
port 65 nsew signal input
rlabel metal3 s 163720 85960 164520 86080 6 i_dout1[10]
port 66 nsew signal input
rlabel metal2 s 135074 0 135130 800 6 i_dout1[11]
port 67 nsew signal input
rlabel metal3 s 163720 94528 164520 94648 6 i_dout1[12]
port 68 nsew signal input
rlabel metal3 s 163720 100104 164520 100224 6 i_dout1[13]
port 69 nsew signal input
rlabel metal3 s 163720 102960 164520 103080 6 i_dout1[14]
port 70 nsew signal input
rlabel metal2 s 144734 0 144790 800 6 i_dout1[15]
port 71 nsew signal input
rlabel metal3 s 163720 111392 164520 111512 6 i_dout1[16]
port 72 nsew signal input
rlabel metal2 s 148598 0 148654 800 6 i_dout1[17]
port 73 nsew signal input
rlabel metal3 s 0 104048 800 104168 6 i_dout1[18]
port 74 nsew signal input
rlabel metal2 s 150530 0 150586 800 6 i_dout1[19]
port 75 nsew signal input
rlabel metal2 s 108486 165864 108542 166664 6 i_dout1[1]
port 76 nsew signal input
rlabel metal3 s 0 112344 800 112464 6 i_dout1[20]
port 77 nsew signal input
rlabel metal3 s 0 120640 800 120760 6 i_dout1[21]
port 78 nsew signal input
rlabel metal2 s 147034 165864 147090 166664 6 i_dout1[22]
port 79 nsew signal input
rlabel metal2 s 154302 0 154358 800 6 i_dout1[23]
port 80 nsew signal input
rlabel metal3 s 163720 142536 164520 142656 6 i_dout1[24]
port 81 nsew signal input
rlabel metal3 s 0 131792 800 131912 6 i_dout1[25]
port 82 nsew signal input
rlabel metal3 s 0 137368 800 137488 6 i_dout1[26]
port 83 nsew signal input
rlabel metal3 s 0 142944 800 143064 6 i_dout1[27]
port 84 nsew signal input
rlabel metal3 s 163720 156544 164520 156664 6 i_dout1[28]
port 85 nsew signal input
rlabel metal3 s 0 151240 800 151360 6 i_dout1[29]
port 86 nsew signal input
rlabel metal3 s 163720 29520 164520 29640 6 i_dout1[2]
port 87 nsew signal input
rlabel metal2 s 162122 165864 162178 166664 6 i_dout1[30]
port 88 nsew signal input
rlabel metal3 s 163720 165112 164520 165232 6 i_dout1[31]
port 89 nsew signal input
rlabel metal3 s 0 29112 800 29232 6 i_dout1[3]
port 90 nsew signal input
rlabel metal3 s 0 42984 800 43104 6 i_dout1[4]
port 91 nsew signal input
rlabel metal3 s 163720 54952 164520 55072 6 i_dout1[5]
port 92 nsew signal input
rlabel metal3 s 163720 60664 164520 60784 6 i_dout1[6]
port 93 nsew signal input
rlabel metal2 s 127438 0 127494 800 6 i_dout1[7]
port 94 nsew signal input
rlabel metal2 s 126426 165864 126482 166664 6 i_dout1[8]
port 95 nsew signal input
rlabel metal2 s 132222 0 132278 800 6 i_dout1[9]
port 96 nsew signal input
rlabel metal3 s 163720 6944 164520 7064 6 i_dout1_1[0]
port 97 nsew signal input
rlabel metal2 s 130106 165864 130162 166664 6 i_dout1_1[10]
port 98 nsew signal input
rlabel metal3 s 0 81880 800 82000 6 i_dout1_1[11]
port 99 nsew signal input
rlabel metal2 s 137006 0 137062 800 6 i_dout1_1[12]
port 100 nsew signal input
rlabel metal2 s 139950 0 140006 800 6 i_dout1_1[13]
port 101 nsew signal input
rlabel metal2 s 142802 0 142858 800 6 i_dout1_1[14]
port 102 nsew signal input
rlabel metal2 s 134890 165864 134946 166664 6 i_dout1_1[15]
port 103 nsew signal input
rlabel metal2 s 136730 165864 136786 166664 6 i_dout1_1[16]
port 104 nsew signal input
rlabel metal3 s 0 98472 800 98592 6 i_dout1_1[17]
port 105 nsew signal input
rlabel metal3 s 163720 119960 164520 120080 6 i_dout1_1[18]
port 106 nsew signal input
rlabel metal2 s 140502 165864 140558 166664 6 i_dout1_1[19]
port 107 nsew signal input
rlabel metal2 s 112994 0 113050 800 6 i_dout1_1[1]
port 108 nsew signal input
rlabel metal2 s 143354 165864 143410 166664 6 i_dout1_1[20]
port 109 nsew signal input
rlabel metal3 s 0 117920 800 118040 6 i_dout1_1[21]
port 110 nsew signal input
rlabel metal2 s 151450 0 151506 800 6 i_dout1_1[22]
port 111 nsew signal input
rlabel metal2 s 148966 165864 149022 166664 6 i_dout1_1[23]
port 112 nsew signal input
rlabel metal3 s 0 129072 800 129192 6 i_dout1_1[24]
port 113 nsew signal input
rlabel metal2 s 152738 165864 152794 166664 6 i_dout1_1[25]
port 114 nsew signal input
rlabel metal3 s 163720 150968 164520 151088 6 i_dout1_1[26]
port 115 nsew signal input
rlabel metal2 s 155498 165864 155554 166664 6 i_dout1_1[27]
port 116 nsew signal input
rlabel metal3 s 0 145664 800 145784 6 i_dout1_1[28]
port 117 nsew signal input
rlabel metal2 s 162030 0 162086 800 6 i_dout1_1[29]
port 118 nsew signal input
rlabel metal3 s 163720 26664 164520 26784 6 i_dout1_1[2]
port 119 nsew signal input
rlabel metal3 s 163720 162256 164520 162376 6 i_dout1_1[30]
port 120 nsew signal input
rlabel metal2 s 163962 165864 164018 166664 6 i_dout1_1[31]
port 121 nsew signal input
rlabel metal3 s 0 26256 800 26376 6 i_dout1_1[3]
port 122 nsew signal input
rlabel metal2 s 115110 165864 115166 166664 6 i_dout1_1[4]
port 123 nsew signal input
rlabel metal3 s 163720 52096 164520 52216 6 i_dout1_1[5]
port 124 nsew signal input
rlabel metal3 s 0 59576 800 59696 6 i_dout1_1[6]
port 125 nsew signal input
rlabel metal3 s 0 62432 800 62552 6 i_dout1_1[7]
port 126 nsew signal input
rlabel metal3 s 0 73448 800 73568 6 i_dout1_1[8]
port 127 nsew signal input
rlabel metal2 s 128266 165864 128322 166664 6 i_dout1_1[9]
port 128 nsew signal input
rlabel metal2 s 478 165864 534 166664 6 io_in[0]
port 129 nsew signal input
rlabel metal2 s 28630 165864 28686 166664 6 io_in[10]
port 130 nsew signal input
rlabel metal2 s 31482 165864 31538 166664 6 io_in[11]
port 131 nsew signal input
rlabel metal2 s 34242 165864 34298 166664 6 io_in[12]
port 132 nsew signal input
rlabel metal2 s 37094 165864 37150 166664 6 io_in[13]
port 133 nsew signal input
rlabel metal2 s 39946 165864 40002 166664 6 io_in[14]
port 134 nsew signal input
rlabel metal2 s 42706 165864 42762 166664 6 io_in[15]
port 135 nsew signal input
rlabel metal2 s 45558 165864 45614 166664 6 io_in[16]
port 136 nsew signal input
rlabel metal2 s 48410 165864 48466 166664 6 io_in[17]
port 137 nsew signal input
rlabel metal2 s 51170 165864 51226 166664 6 io_in[18]
port 138 nsew signal input
rlabel metal2 s 54022 165864 54078 166664 6 io_in[19]
port 139 nsew signal input
rlabel metal2 s 3238 165864 3294 166664 6 io_in[1]
port 140 nsew signal input
rlabel metal2 s 56874 165864 56930 166664 6 io_in[20]
port 141 nsew signal input
rlabel metal2 s 59634 165864 59690 166664 6 io_in[21]
port 142 nsew signal input
rlabel metal2 s 62486 165864 62542 166664 6 io_in[22]
port 143 nsew signal input
rlabel metal2 s 65246 165864 65302 166664 6 io_in[23]
port 144 nsew signal input
rlabel metal2 s 68098 165864 68154 166664 6 io_in[24]
port 145 nsew signal input
rlabel metal2 s 70950 165864 71006 166664 6 io_in[25]
port 146 nsew signal input
rlabel metal2 s 73710 165864 73766 166664 6 io_in[26]
port 147 nsew signal input
rlabel metal2 s 76562 165864 76618 166664 6 io_in[27]
port 148 nsew signal input
rlabel metal2 s 79414 165864 79470 166664 6 io_in[28]
port 149 nsew signal input
rlabel metal2 s 82174 165864 82230 166664 6 io_in[29]
port 150 nsew signal input
rlabel metal2 s 6090 165864 6146 166664 6 io_in[2]
port 151 nsew signal input
rlabel metal2 s 85026 165864 85082 166664 6 io_in[30]
port 152 nsew signal input
rlabel metal2 s 87878 165864 87934 166664 6 io_in[31]
port 153 nsew signal input
rlabel metal2 s 90638 165864 90694 166664 6 io_in[32]
port 154 nsew signal input
rlabel metal2 s 93490 165864 93546 166664 6 io_in[33]
port 155 nsew signal input
rlabel metal2 s 96342 165864 96398 166664 6 io_in[34]
port 156 nsew signal input
rlabel metal2 s 99102 165864 99158 166664 6 io_in[35]
port 157 nsew signal input
rlabel metal2 s 101954 165864 102010 166664 6 io_in[36]
port 158 nsew signal input
rlabel metal2 s 104806 165864 104862 166664 6 io_in[37]
port 159 nsew signal input
rlabel metal2 s 8850 165864 8906 166664 6 io_in[3]
port 160 nsew signal input
rlabel metal2 s 11702 165864 11758 166664 6 io_in[4]
port 161 nsew signal input
rlabel metal2 s 14554 165864 14610 166664 6 io_in[5]
port 162 nsew signal input
rlabel metal2 s 17314 165864 17370 166664 6 io_in[6]
port 163 nsew signal input
rlabel metal2 s 20166 165864 20222 166664 6 io_in[7]
port 164 nsew signal input
rlabel metal2 s 23018 165864 23074 166664 6 io_in[8]
port 165 nsew signal input
rlabel metal2 s 25778 165864 25834 166664 6 io_in[9]
port 166 nsew signal input
rlabel metal2 s 1398 165864 1454 166664 6 io_oeb[0]
port 167 nsew signal output
rlabel metal2 s 29550 165864 29606 166664 6 io_oeb[10]
port 168 nsew signal output
rlabel metal2 s 32402 165864 32458 166664 6 io_oeb[11]
port 169 nsew signal output
rlabel metal2 s 35254 165864 35310 166664 6 io_oeb[12]
port 170 nsew signal output
rlabel metal2 s 38014 165864 38070 166664 6 io_oeb[13]
port 171 nsew signal output
rlabel metal2 s 40866 165864 40922 166664 6 io_oeb[14]
port 172 nsew signal output
rlabel metal2 s 43626 165864 43682 166664 6 io_oeb[15]
port 173 nsew signal output
rlabel metal2 s 46478 165864 46534 166664 6 io_oeb[16]
port 174 nsew signal output
rlabel metal2 s 49330 165864 49386 166664 6 io_oeb[17]
port 175 nsew signal output
rlabel metal2 s 52090 165864 52146 166664 6 io_oeb[18]
port 176 nsew signal output
rlabel metal2 s 54942 165864 54998 166664 6 io_oeb[19]
port 177 nsew signal output
rlabel metal2 s 4158 165864 4214 166664 6 io_oeb[1]
port 178 nsew signal output
rlabel metal2 s 57794 165864 57850 166664 6 io_oeb[20]
port 179 nsew signal output
rlabel metal2 s 60554 165864 60610 166664 6 io_oeb[21]
port 180 nsew signal output
rlabel metal2 s 63406 165864 63462 166664 6 io_oeb[22]
port 181 nsew signal output
rlabel metal2 s 66258 165864 66314 166664 6 io_oeb[23]
port 182 nsew signal output
rlabel metal2 s 69018 165864 69074 166664 6 io_oeb[24]
port 183 nsew signal output
rlabel metal2 s 71870 165864 71926 166664 6 io_oeb[25]
port 184 nsew signal output
rlabel metal2 s 74722 165864 74778 166664 6 io_oeb[26]
port 185 nsew signal output
rlabel metal2 s 77482 165864 77538 166664 6 io_oeb[27]
port 186 nsew signal output
rlabel metal2 s 80334 165864 80390 166664 6 io_oeb[28]
port 187 nsew signal output
rlabel metal2 s 83186 165864 83242 166664 6 io_oeb[29]
port 188 nsew signal output
rlabel metal2 s 7010 165864 7066 166664 6 io_oeb[2]
port 189 nsew signal output
rlabel metal2 s 85946 165864 86002 166664 6 io_oeb[30]
port 190 nsew signal output
rlabel metal2 s 88798 165864 88854 166664 6 io_oeb[31]
port 191 nsew signal output
rlabel metal2 s 91650 165864 91706 166664 6 io_oeb[32]
port 192 nsew signal output
rlabel metal2 s 94410 165864 94466 166664 6 io_oeb[33]
port 193 nsew signal output
rlabel metal2 s 97262 165864 97318 166664 6 io_oeb[34]
port 194 nsew signal output
rlabel metal2 s 100114 165864 100170 166664 6 io_oeb[35]
port 195 nsew signal output
rlabel metal2 s 102874 165864 102930 166664 6 io_oeb[36]
port 196 nsew signal output
rlabel metal2 s 105726 165864 105782 166664 6 io_oeb[37]
port 197 nsew signal output
rlabel metal2 s 9862 165864 9918 166664 6 io_oeb[3]
port 198 nsew signal output
rlabel metal2 s 12622 165864 12678 166664 6 io_oeb[4]
port 199 nsew signal output
rlabel metal2 s 15474 165864 15530 166664 6 io_oeb[5]
port 200 nsew signal output
rlabel metal2 s 18326 165864 18382 166664 6 io_oeb[6]
port 201 nsew signal output
rlabel metal2 s 21086 165864 21142 166664 6 io_oeb[7]
port 202 nsew signal output
rlabel metal2 s 23938 165864 23994 166664 6 io_oeb[8]
port 203 nsew signal output
rlabel metal2 s 26790 165864 26846 166664 6 io_oeb[9]
port 204 nsew signal output
rlabel metal2 s 2318 165864 2374 166664 6 io_out[0]
port 205 nsew signal output
rlabel metal2 s 30470 165864 30526 166664 6 io_out[10]
port 206 nsew signal output
rlabel metal2 s 33322 165864 33378 166664 6 io_out[11]
port 207 nsew signal output
rlabel metal2 s 36174 165864 36230 166664 6 io_out[12]
port 208 nsew signal output
rlabel metal2 s 38934 165864 38990 166664 6 io_out[13]
port 209 nsew signal output
rlabel metal2 s 41786 165864 41842 166664 6 io_out[14]
port 210 nsew signal output
rlabel metal2 s 44638 165864 44694 166664 6 io_out[15]
port 211 nsew signal output
rlabel metal2 s 47398 165864 47454 166664 6 io_out[16]
port 212 nsew signal output
rlabel metal2 s 50250 165864 50306 166664 6 io_out[17]
port 213 nsew signal output
rlabel metal2 s 53102 165864 53158 166664 6 io_out[18]
port 214 nsew signal output
rlabel metal2 s 55862 165864 55918 166664 6 io_out[19]
port 215 nsew signal output
rlabel metal2 s 5170 165864 5226 166664 6 io_out[1]
port 216 nsew signal output
rlabel metal2 s 58714 165864 58770 166664 6 io_out[20]
port 217 nsew signal output
rlabel metal2 s 61566 165864 61622 166664 6 io_out[21]
port 218 nsew signal output
rlabel metal2 s 64326 165864 64382 166664 6 io_out[22]
port 219 nsew signal output
rlabel metal2 s 67178 165864 67234 166664 6 io_out[23]
port 220 nsew signal output
rlabel metal2 s 70030 165864 70086 166664 6 io_out[24]
port 221 nsew signal output
rlabel metal2 s 72790 165864 72846 166664 6 io_out[25]
port 222 nsew signal output
rlabel metal2 s 75642 165864 75698 166664 6 io_out[26]
port 223 nsew signal output
rlabel metal2 s 78494 165864 78550 166664 6 io_out[27]
port 224 nsew signal output
rlabel metal2 s 81254 165864 81310 166664 6 io_out[28]
port 225 nsew signal output
rlabel metal2 s 84106 165864 84162 166664 6 io_out[29]
port 226 nsew signal output
rlabel metal2 s 7930 165864 7986 166664 6 io_out[2]
port 227 nsew signal output
rlabel metal2 s 86866 165864 86922 166664 6 io_out[30]
port 228 nsew signal output
rlabel metal2 s 89718 165864 89774 166664 6 io_out[31]
port 229 nsew signal output
rlabel metal2 s 92570 165864 92626 166664 6 io_out[32]
port 230 nsew signal output
rlabel metal2 s 95330 165864 95386 166664 6 io_out[33]
port 231 nsew signal output
rlabel metal2 s 98182 165864 98238 166664 6 io_out[34]
port 232 nsew signal output
rlabel metal2 s 101034 165864 101090 166664 6 io_out[35]
port 233 nsew signal output
rlabel metal2 s 103794 165864 103850 166664 6 io_out[36]
port 234 nsew signal output
rlabel metal2 s 106646 165864 106702 166664 6 io_out[37]
port 235 nsew signal output
rlabel metal2 s 10782 165864 10838 166664 6 io_out[3]
port 236 nsew signal output
rlabel metal2 s 13634 165864 13690 166664 6 io_out[4]
port 237 nsew signal output
rlabel metal2 s 16394 165864 16450 166664 6 io_out[5]
port 238 nsew signal output
rlabel metal2 s 19246 165864 19302 166664 6 io_out[6]
port 239 nsew signal output
rlabel metal2 s 22006 165864 22062 166664 6 io_out[7]
port 240 nsew signal output
rlabel metal2 s 24858 165864 24914 166664 6 io_out[8]
port 241 nsew signal output
rlabel metal2 s 27710 165864 27766 166664 6 io_out[9]
port 242 nsew signal output
rlabel metal2 s 102414 0 102470 800 6 irq[0]
port 243 nsew signal output
rlabel metal2 s 103334 0 103390 800 6 irq[1]
port 244 nsew signal output
rlabel metal2 s 104346 0 104402 800 6 irq[2]
port 245 nsew signal output
rlabel metal3 s 0 4088 800 4208 6 o_addr1[0]
port 246 nsew signal output
rlabel metal2 s 113914 0 113970 800 6 o_addr1[1]
port 247 nsew signal output
rlabel metal3 s 0 17960 800 18080 6 o_addr1[2]
port 248 nsew signal output
rlabel metal2 s 120722 0 120778 800 6 o_addr1[3]
port 249 nsew signal output
rlabel metal3 s 163720 43664 164520 43784 6 o_addr1[4]
port 250 nsew signal output
rlabel metal3 s 0 54000 800 54120 6 o_addr1[5]
port 251 nsew signal output
rlabel metal2 s 125506 0 125562 800 6 o_addr1[6]
port 252 nsew signal output
rlabel metal2 s 124494 165864 124550 166664 6 o_addr1[7]
port 253 nsew signal output
rlabel metal3 s 163720 69096 164520 69216 6 o_addr1[8]
port 254 nsew signal output
rlabel metal2 s 110142 0 110198 800 6 o_addr1_1[0]
port 255 nsew signal output
rlabel metal3 s 0 15240 800 15360 6 o_addr1_1[1]
port 256 nsew signal output
rlabel metal3 s 163720 32376 164520 32496 6 o_addr1_1[2]
port 257 nsew signal output
rlabel metal2 s 119710 0 119766 800 6 o_addr1_1[3]
port 258 nsew signal output
rlabel metal2 s 116030 165864 116086 166664 6 o_addr1_1[4]
port 259 nsew signal output
rlabel metal2 s 117962 165864 118018 166664 6 o_addr1_1[5]
port 260 nsew signal output
rlabel metal2 s 119802 165864 119858 166664 6 o_addr1_1[6]
port 261 nsew signal output
rlabel metal3 s 0 65152 800 65272 6 o_addr1_1[7]
port 262 nsew signal output
rlabel metal2 s 127346 165864 127402 166664 6 o_addr1_1[8]
port 263 nsew signal output
rlabel metal3 s 163720 1368 164520 1488 6 o_csb0
port 264 nsew signal output
rlabel metal3 s 0 1368 800 1488 6 o_csb0_1
port 265 nsew signal output
rlabel metal2 s 105266 0 105322 800 6 o_csb1
port 266 nsew signal output
rlabel metal2 s 106278 0 106334 800 6 o_csb1_1
port 267 nsew signal output
rlabel metal3 s 0 6808 800 6928 6 o_din0[0]
port 268 nsew signal output
rlabel metal2 s 131118 165864 131174 166664 6 o_din0[10]
port 269 nsew signal output
rlabel metal2 s 136086 0 136142 800 6 o_din0[11]
port 270 nsew signal output
rlabel metal2 s 138938 0 138994 800 6 o_din0[12]
port 271 nsew signal output
rlabel metal3 s 0 87320 800 87440 6 o_din0[13]
port 272 nsew signal output
rlabel metal3 s 163720 108536 164520 108656 6 o_din0[14]
port 273 nsew signal output
rlabel metal2 s 135810 165864 135866 166664 6 o_din0[15]
port 274 nsew signal output
rlabel metal2 s 146666 0 146722 800 6 o_din0[16]
port 275 nsew signal output
rlabel metal2 s 149518 0 149574 800 6 o_din0[17]
port 276 nsew signal output
rlabel metal3 s 0 106768 800 106888 6 o_din0[18]
port 277 nsew signal output
rlabel metal2 s 141422 165864 141478 166664 6 o_din0[19]
port 278 nsew signal output
rlabel metal3 s 163720 21088 164520 21208 6 o_din0[1]
port 279 nsew signal output
rlabel metal2 s 144274 165864 144330 166664 6 o_din0[20]
port 280 nsew signal output
rlabel metal2 s 145194 165864 145250 166664 6 o_din0[21]
port 281 nsew signal output
rlabel metal2 s 148046 165864 148102 166664 6 o_din0[22]
port 282 nsew signal output
rlabel metal2 s 155314 0 155370 800 6 o_din0[23]
port 283 nsew signal output
rlabel metal2 s 156234 0 156290 800 6 o_din0[24]
port 284 nsew signal output
rlabel metal2 s 153658 165864 153714 166664 6 o_din0[25]
port 285 nsew signal output
rlabel metal3 s 163720 153824 164520 153944 6 o_din0[26]
port 286 nsew signal output
rlabel metal2 s 158350 165864 158406 166664 6 o_din0[27]
port 287 nsew signal output
rlabel metal2 s 160098 0 160154 800 6 o_din0[28]
port 288 nsew signal output
rlabel metal3 s 0 156816 800 156936 6 o_din0[29]
port 289 nsew signal output
rlabel metal2 s 111338 165864 111394 166664 6 o_din0[2]
port 290 nsew signal output
rlabel metal2 s 163042 165864 163098 166664 6 o_din0[30]
port 291 nsew signal output
rlabel metal2 s 163962 0 164018 800 6 o_din0[31]
port 292 nsew signal output
rlabel metal2 s 113270 165864 113326 166664 6 o_din0[3]
port 293 nsew signal output
rlabel metal3 s 163720 46520 164520 46640 6 o_din0[4]
port 294 nsew signal output
rlabel metal2 s 123574 0 123630 800 6 o_din0[5]
port 295 nsew signal output
rlabel metal2 s 121734 165864 121790 166664 6 o_din0[6]
port 296 nsew signal output
rlabel metal2 s 128358 0 128414 800 6 o_din0[7]
port 297 nsew signal output
rlabel metal3 s 163720 74672 164520 74792 6 o_din0[8]
port 298 nsew signal output
rlabel metal3 s 163720 80384 164520 80504 6 o_din0[9]
port 299 nsew signal output
rlabel metal2 s 111062 0 111118 800 6 o_din0_1[0]
port 300 nsew signal output
rlabel metal3 s 163720 88816 164520 88936 6 o_din0_1[10]
port 301 nsew signal output
rlabel metal2 s 132038 165864 132094 166664 6 o_din0_1[11]
port 302 nsew signal output
rlabel metal2 s 138018 0 138074 800 6 o_din0_1[12]
port 303 nsew signal output
rlabel metal2 s 140870 0 140926 800 6 o_din0_1[13]
port 304 nsew signal output
rlabel metal3 s 163720 105816 164520 105936 6 o_din0_1[14]
port 305 nsew signal output
rlabel metal3 s 0 92896 800 93016 6 o_din0_1[15]
port 306 nsew signal output
rlabel metal2 s 145654 0 145710 800 6 o_din0_1[16]
port 307 nsew signal output
rlabel metal3 s 0 101328 800 101448 6 o_din0_1[17]
port 308 nsew signal output
rlabel metal3 s 163720 122680 164520 122800 6 o_din0_1[18]
port 309 nsew signal output
rlabel metal3 s 0 109624 800 109744 6 o_din0_1[19]
port 310 nsew signal output
rlabel metal3 s 163720 18232 164520 18352 6 o_din0_1[1]
port 311 nsew signal output
rlabel metal3 s 163720 131248 164520 131368 6 o_din0_1[20]
port 312 nsew signal output
rlabel metal3 s 0 123496 800 123616 6 o_din0_1[21]
port 313 nsew signal output
rlabel metal2 s 152462 0 152518 800 6 o_din0_1[22]
port 314 nsew signal output
rlabel metal3 s 0 126216 800 126336 6 o_din0_1[23]
port 315 nsew signal output
rlabel metal3 s 163720 145256 164520 145376 6 o_din0_1[24]
port 316 nsew signal output
rlabel metal3 s 163720 148112 164520 148232 6 o_din0_1[25]
port 317 nsew signal output
rlabel metal2 s 154578 165864 154634 166664 6 o_din0_1[26]
port 318 nsew signal output
rlabel metal2 s 157430 165864 157486 166664 6 o_din0_1[27]
port 319 nsew signal output
rlabel metal2 s 159178 0 159234 800 6 o_din0_1[28]
port 320 nsew signal output
rlabel metal3 s 0 153960 800 154080 6 o_din0_1[29]
port 321 nsew signal output
rlabel metal3 s 0 20680 800 20800 6 o_din0_1[2]
port 322 nsew signal output
rlabel metal3 s 0 159536 800 159656 6 o_din0_1[30]
port 323 nsew signal output
rlabel metal2 s 163042 0 163098 800 6 o_din0_1[31]
port 324 nsew signal output
rlabel metal3 s 163720 40808 164520 40928 6 o_din0_1[3]
port 325 nsew signal output
rlabel metal3 s 0 45704 800 45824 6 o_din0_1[4]
port 326 nsew signal output
rlabel metal2 s 122562 0 122618 800 6 o_din0_1[5]
port 327 nsew signal output
rlabel metal2 s 120722 165864 120778 166664 6 o_din0_1[6]
port 328 nsew signal output
rlabel metal3 s 0 68008 800 68128 6 o_din0_1[7]
port 329 nsew signal output
rlabel metal3 s 163720 71952 164520 72072 6 o_din0_1[8]
port 330 nsew signal output
rlabel metal3 s 0 79024 800 79144 6 o_din0_1[9]
port 331 nsew signal output
rlabel metal3 s 0 9664 800 9784 6 o_waddr0[0]
port 332 nsew signal output
rlabel metal3 s 163720 23944 164520 24064 6 o_waddr0[1]
port 333 nsew signal output
rlabel metal2 s 117778 0 117834 800 6 o_waddr0[2]
port 334 nsew signal output
rlabel metal3 s 0 31832 800 31952 6 o_waddr0[3]
port 335 nsew signal output
rlabel metal2 s 116950 165864 117006 166664 6 o_waddr0[4]
port 336 nsew signal output
rlabel metal2 s 124494 0 124550 800 6 o_waddr0[5]
port 337 nsew signal output
rlabel metal2 s 126426 0 126482 800 6 o_waddr0[6]
port 338 nsew signal output
rlabel metal2 s 125414 165864 125470 166664 6 o_waddr0[7]
port 339 nsew signal output
rlabel metal2 s 130290 0 130346 800 6 o_waddr0[8]
port 340 nsew signal output
rlabel metal2 s 107566 165864 107622 166664 6 o_waddr0_1[0]
port 341 nsew signal output
rlabel metal2 s 114926 0 114982 800 6 o_waddr0_1[1]
port 342 nsew signal output
rlabel metal3 s 0 23536 800 23656 6 o_waddr0_1[2]
port 343 nsew signal output
rlabel metal2 s 121642 0 121698 800 6 o_waddr0_1[3]
port 344 nsew signal output
rlabel metal3 s 0 48560 800 48680 6 o_waddr0_1[4]
port 345 nsew signal output
rlabel metal3 s 163720 57808 164520 57928 6 o_waddr0_1[5]
port 346 nsew signal output
rlabel metal2 s 122654 165864 122710 166664 6 o_waddr0_1[6]
port 347 nsew signal output
rlabel metal3 s 163720 66240 164520 66360 6 o_waddr0_1[7]
port 348 nsew signal output
rlabel metal2 s 129370 0 129426 800 6 o_waddr0_1[8]
port 349 nsew signal output
rlabel metal2 s 107198 0 107254 800 6 o_web0
port 350 nsew signal output
rlabel metal2 s 108210 0 108266 800 6 o_web0_1
port 351 nsew signal output
rlabel metal2 s 111982 0 112038 800 6 o_wmask0[0]
port 352 nsew signal output
rlabel metal2 s 110418 165864 110474 166664 6 o_wmask0[1]
port 353 nsew signal output
rlabel metal2 s 112258 165864 112314 166664 6 o_wmask0[2]
port 354 nsew signal output
rlabel metal3 s 0 34688 800 34808 6 o_wmask0[3]
port 355 nsew signal output
rlabel metal3 s 0 12384 800 12504 6 o_wmask0_1[0]
port 356 nsew signal output
rlabel metal2 s 109498 165864 109554 166664 6 o_wmask0_1[1]
port 357 nsew signal output
rlabel metal2 s 118790 0 118846 800 6 o_wmask0_1[2]
port 358 nsew signal output
rlabel metal2 s 114190 165864 114246 166664 6 o_wmask0_1[3]
port 359 nsew signal output
rlabel metal4 s 4208 2128 4528 164336 6 vccd1
port 360 nsew power input
rlabel metal4 s 34928 2128 35248 164336 6 vccd1
port 360 nsew power input
rlabel metal4 s 65648 2128 65968 164336 6 vccd1
port 360 nsew power input
rlabel metal4 s 96368 2128 96688 164336 6 vccd1
port 360 nsew power input
rlabel metal4 s 127088 2128 127408 164336 6 vccd1
port 360 nsew power input
rlabel metal4 s 157808 2128 158128 164336 6 vccd1
port 360 nsew power input
rlabel metal4 s 19568 2128 19888 164336 6 vssd1
port 361 nsew ground input
rlabel metal4 s 50288 2128 50608 164336 6 vssd1
port 361 nsew ground input
rlabel metal4 s 81008 2128 81328 164336 6 vssd1
port 361 nsew ground input
rlabel metal4 s 111728 2128 112048 164336 6 vssd1
port 361 nsew ground input
rlabel metal4 s 142448 2128 142768 164336 6 vssd1
port 361 nsew ground input
rlabel metal2 s 478 0 534 800 6 wb_clk_i
port 362 nsew signal input
rlabel metal2 s 1398 0 1454 800 6 wb_rst_i
port 363 nsew signal input
rlabel metal2 s 2318 0 2374 800 6 wbs_ack_o
port 364 nsew signal output
rlabel metal2 s 6182 0 6238 800 6 wbs_adr_i[0]
port 365 nsew signal input
rlabel metal2 s 38934 0 38990 800 6 wbs_adr_i[10]
port 366 nsew signal input
rlabel metal2 s 41786 0 41842 800 6 wbs_adr_i[11]
port 367 nsew signal input
rlabel metal2 s 44638 0 44694 800 6 wbs_adr_i[12]
port 368 nsew signal input
rlabel metal2 s 47582 0 47638 800 6 wbs_adr_i[13]
port 369 nsew signal input
rlabel metal2 s 50434 0 50490 800 6 wbs_adr_i[14]
port 370 nsew signal input
rlabel metal2 s 53378 0 53434 800 6 wbs_adr_i[15]
port 371 nsew signal input
rlabel metal2 s 56230 0 56286 800 6 wbs_adr_i[16]
port 372 nsew signal input
rlabel metal2 s 59082 0 59138 800 6 wbs_adr_i[17]
port 373 nsew signal input
rlabel metal2 s 62026 0 62082 800 6 wbs_adr_i[18]
port 374 nsew signal input
rlabel metal2 s 64878 0 64934 800 6 wbs_adr_i[19]
port 375 nsew signal input
rlabel metal2 s 10046 0 10102 800 6 wbs_adr_i[1]
port 376 nsew signal input
rlabel metal2 s 67730 0 67786 800 6 wbs_adr_i[20]
port 377 nsew signal input
rlabel metal2 s 70674 0 70730 800 6 wbs_adr_i[21]
port 378 nsew signal input
rlabel metal2 s 73526 0 73582 800 6 wbs_adr_i[22]
port 379 nsew signal input
rlabel metal2 s 76470 0 76526 800 6 wbs_adr_i[23]
port 380 nsew signal input
rlabel metal2 s 79322 0 79378 800 6 wbs_adr_i[24]
port 381 nsew signal input
rlabel metal2 s 82174 0 82230 800 6 wbs_adr_i[25]
port 382 nsew signal input
rlabel metal2 s 85118 0 85174 800 6 wbs_adr_i[26]
port 383 nsew signal input
rlabel metal2 s 87970 0 88026 800 6 wbs_adr_i[27]
port 384 nsew signal input
rlabel metal2 s 90822 0 90878 800 6 wbs_adr_i[28]
port 385 nsew signal input
rlabel metal2 s 93766 0 93822 800 6 wbs_adr_i[29]
port 386 nsew signal input
rlabel metal2 s 13910 0 13966 800 6 wbs_adr_i[2]
port 387 nsew signal input
rlabel metal2 s 96618 0 96674 800 6 wbs_adr_i[30]
port 388 nsew signal input
rlabel metal2 s 99470 0 99526 800 6 wbs_adr_i[31]
port 389 nsew signal input
rlabel metal2 s 17774 0 17830 800 6 wbs_adr_i[3]
port 390 nsew signal input
rlabel metal2 s 21638 0 21694 800 6 wbs_adr_i[4]
port 391 nsew signal input
rlabel metal2 s 24490 0 24546 800 6 wbs_adr_i[5]
port 392 nsew signal input
rlabel metal2 s 27342 0 27398 800 6 wbs_adr_i[6]
port 393 nsew signal input
rlabel metal2 s 30286 0 30342 800 6 wbs_adr_i[7]
port 394 nsew signal input
rlabel metal2 s 33138 0 33194 800 6 wbs_adr_i[8]
port 395 nsew signal input
rlabel metal2 s 35990 0 36046 800 6 wbs_adr_i[9]
port 396 nsew signal input
rlabel metal2 s 3330 0 3386 800 6 wbs_cyc_i
port 397 nsew signal input
rlabel metal2 s 7194 0 7250 800 6 wbs_dat_i[0]
port 398 nsew signal input
rlabel metal2 s 39854 0 39910 800 6 wbs_dat_i[10]
port 399 nsew signal input
rlabel metal2 s 42798 0 42854 800 6 wbs_dat_i[11]
port 400 nsew signal input
rlabel metal2 s 45650 0 45706 800 6 wbs_dat_i[12]
port 401 nsew signal input
rlabel metal2 s 48502 0 48558 800 6 wbs_dat_i[13]
port 402 nsew signal input
rlabel metal2 s 51446 0 51502 800 6 wbs_dat_i[14]
port 403 nsew signal input
rlabel metal2 s 54298 0 54354 800 6 wbs_dat_i[15]
port 404 nsew signal input
rlabel metal2 s 57150 0 57206 800 6 wbs_dat_i[16]
port 405 nsew signal input
rlabel metal2 s 60094 0 60150 800 6 wbs_dat_i[17]
port 406 nsew signal input
rlabel metal2 s 62946 0 63002 800 6 wbs_dat_i[18]
port 407 nsew signal input
rlabel metal2 s 65890 0 65946 800 6 wbs_dat_i[19]
port 408 nsew signal input
rlabel metal2 s 11058 0 11114 800 6 wbs_dat_i[1]
port 409 nsew signal input
rlabel metal2 s 68742 0 68798 800 6 wbs_dat_i[20]
port 410 nsew signal input
rlabel metal2 s 71594 0 71650 800 6 wbs_dat_i[21]
port 411 nsew signal input
rlabel metal2 s 74538 0 74594 800 6 wbs_dat_i[22]
port 412 nsew signal input
rlabel metal2 s 77390 0 77446 800 6 wbs_dat_i[23]
port 413 nsew signal input
rlabel metal2 s 80242 0 80298 800 6 wbs_dat_i[24]
port 414 nsew signal input
rlabel metal2 s 83186 0 83242 800 6 wbs_dat_i[25]
port 415 nsew signal input
rlabel metal2 s 86038 0 86094 800 6 wbs_dat_i[26]
port 416 nsew signal input
rlabel metal2 s 88890 0 88946 800 6 wbs_dat_i[27]
port 417 nsew signal input
rlabel metal2 s 91834 0 91890 800 6 wbs_dat_i[28]
port 418 nsew signal input
rlabel metal2 s 94686 0 94742 800 6 wbs_dat_i[29]
port 419 nsew signal input
rlabel metal2 s 14830 0 14886 800 6 wbs_dat_i[2]
port 420 nsew signal input
rlabel metal2 s 97630 0 97686 800 6 wbs_dat_i[30]
port 421 nsew signal input
rlabel metal2 s 100482 0 100538 800 6 wbs_dat_i[31]
port 422 nsew signal input
rlabel metal2 s 18694 0 18750 800 6 wbs_dat_i[3]
port 423 nsew signal input
rlabel metal2 s 22558 0 22614 800 6 wbs_dat_i[4]
port 424 nsew signal input
rlabel metal2 s 25410 0 25466 800 6 wbs_dat_i[5]
port 425 nsew signal input
rlabel metal2 s 28354 0 28410 800 6 wbs_dat_i[6]
port 426 nsew signal input
rlabel metal2 s 31206 0 31262 800 6 wbs_dat_i[7]
port 427 nsew signal input
rlabel metal2 s 34058 0 34114 800 6 wbs_dat_i[8]
port 428 nsew signal input
rlabel metal2 s 37002 0 37058 800 6 wbs_dat_i[9]
port 429 nsew signal input
rlabel metal2 s 8114 0 8170 800 6 wbs_dat_o[0]
port 430 nsew signal output
rlabel metal2 s 40866 0 40922 800 6 wbs_dat_o[10]
port 431 nsew signal output
rlabel metal2 s 43718 0 43774 800 6 wbs_dat_o[11]
port 432 nsew signal output
rlabel metal2 s 46570 0 46626 800 6 wbs_dat_o[12]
port 433 nsew signal output
rlabel metal2 s 49514 0 49570 800 6 wbs_dat_o[13]
port 434 nsew signal output
rlabel metal2 s 52366 0 52422 800 6 wbs_dat_o[14]
port 435 nsew signal output
rlabel metal2 s 55310 0 55366 800 6 wbs_dat_o[15]
port 436 nsew signal output
rlabel metal2 s 58162 0 58218 800 6 wbs_dat_o[16]
port 437 nsew signal output
rlabel metal2 s 61014 0 61070 800 6 wbs_dat_o[17]
port 438 nsew signal output
rlabel metal2 s 63958 0 64014 800 6 wbs_dat_o[18]
port 439 nsew signal output
rlabel metal2 s 66810 0 66866 800 6 wbs_dat_o[19]
port 440 nsew signal output
rlabel metal2 s 11978 0 12034 800 6 wbs_dat_o[1]
port 441 nsew signal output
rlabel metal2 s 69662 0 69718 800 6 wbs_dat_o[20]
port 442 nsew signal output
rlabel metal2 s 72606 0 72662 800 6 wbs_dat_o[21]
port 443 nsew signal output
rlabel metal2 s 75458 0 75514 800 6 wbs_dat_o[22]
port 444 nsew signal output
rlabel metal2 s 78310 0 78366 800 6 wbs_dat_o[23]
port 445 nsew signal output
rlabel metal2 s 81254 0 81310 800 6 wbs_dat_o[24]
port 446 nsew signal output
rlabel metal2 s 84106 0 84162 800 6 wbs_dat_o[25]
port 447 nsew signal output
rlabel metal2 s 87050 0 87106 800 6 wbs_dat_o[26]
port 448 nsew signal output
rlabel metal2 s 89902 0 89958 800 6 wbs_dat_o[27]
port 449 nsew signal output
rlabel metal2 s 92754 0 92810 800 6 wbs_dat_o[28]
port 450 nsew signal output
rlabel metal2 s 95698 0 95754 800 6 wbs_dat_o[29]
port 451 nsew signal output
rlabel metal2 s 15842 0 15898 800 6 wbs_dat_o[2]
port 452 nsew signal output
rlabel metal2 s 98550 0 98606 800 6 wbs_dat_o[30]
port 453 nsew signal output
rlabel metal2 s 101402 0 101458 800 6 wbs_dat_o[31]
port 454 nsew signal output
rlabel metal2 s 19706 0 19762 800 6 wbs_dat_o[3]
port 455 nsew signal output
rlabel metal2 s 23478 0 23534 800 6 wbs_dat_o[4]
port 456 nsew signal output
rlabel metal2 s 26422 0 26478 800 6 wbs_dat_o[5]
port 457 nsew signal output
rlabel metal2 s 29274 0 29330 800 6 wbs_dat_o[6]
port 458 nsew signal output
rlabel metal2 s 32218 0 32274 800 6 wbs_dat_o[7]
port 459 nsew signal output
rlabel metal2 s 35070 0 35126 800 6 wbs_dat_o[8]
port 460 nsew signal output
rlabel metal2 s 37922 0 37978 800 6 wbs_dat_o[9]
port 461 nsew signal output
rlabel metal2 s 9126 0 9182 800 6 wbs_sel_i[0]
port 462 nsew signal input
rlabel metal2 s 12898 0 12954 800 6 wbs_sel_i[1]
port 463 nsew signal input
rlabel metal2 s 16762 0 16818 800 6 wbs_sel_i[2]
port 464 nsew signal input
rlabel metal2 s 20626 0 20682 800 6 wbs_sel_i[3]
port 465 nsew signal input
rlabel metal2 s 4250 0 4306 800 6 wbs_stb_i
port 466 nsew signal input
rlabel metal2 s 5262 0 5318 800 6 wbs_we_i
port 467 nsew signal input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 164520 166664
string LEFview TRUE
string GDS_FILE /local/caravel_user_project/openlane/user_proj/runs/user_proj/results/magic/user_proj.gds
string GDS_END 79988650
string GDS_START 1329456
<< end >>

