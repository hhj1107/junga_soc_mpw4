magic
tech sky130A
magscale 1 2
timestamp 1640602795
<< obsli1 >>
rect 1104 1445 164467 164305
<< obsm1 >>
rect 14 8 164482 164336
<< metal2 >>
rect 478 165864 534 166664
rect 1398 165864 1454 166664
rect 2410 165864 2466 166664
rect 3330 165864 3386 166664
rect 4342 165864 4398 166664
rect 5354 165864 5410 166664
rect 6274 165864 6330 166664
rect 7286 165864 7342 166664
rect 8298 165864 8354 166664
rect 9218 165864 9274 166664
rect 10230 165864 10286 166664
rect 11242 165864 11298 166664
rect 12162 165864 12218 166664
rect 13174 165864 13230 166664
rect 14186 165864 14242 166664
rect 15106 165864 15162 166664
rect 16118 165864 16174 166664
rect 17038 165864 17094 166664
rect 18050 165864 18106 166664
rect 19062 165864 19118 166664
rect 19982 165864 20038 166664
rect 20994 165864 21050 166664
rect 22006 165864 22062 166664
rect 22926 165864 22982 166664
rect 23938 165864 23994 166664
rect 24950 165864 25006 166664
rect 25870 165864 25926 166664
rect 26882 165864 26938 166664
rect 27894 165864 27950 166664
rect 28814 165864 28870 166664
rect 29826 165864 29882 166664
rect 30746 165864 30802 166664
rect 31758 165864 31814 166664
rect 32770 165864 32826 166664
rect 33690 165864 33746 166664
rect 34702 165864 34758 166664
rect 35714 165864 35770 166664
rect 36634 165864 36690 166664
rect 37646 165864 37702 166664
rect 38658 165864 38714 166664
rect 39578 165864 39634 166664
rect 40590 165864 40646 166664
rect 41602 165864 41658 166664
rect 42522 165864 42578 166664
rect 43534 165864 43590 166664
rect 44454 165864 44510 166664
rect 45466 165864 45522 166664
rect 46478 165864 46534 166664
rect 47398 165864 47454 166664
rect 48410 165864 48466 166664
rect 49422 165864 49478 166664
rect 50342 165864 50398 166664
rect 51354 165864 51410 166664
rect 52366 165864 52422 166664
rect 53286 165864 53342 166664
rect 54298 165864 54354 166664
rect 55310 165864 55366 166664
rect 56230 165864 56286 166664
rect 57242 165864 57298 166664
rect 58162 165864 58218 166664
rect 59174 165864 59230 166664
rect 60186 165864 60242 166664
rect 61106 165864 61162 166664
rect 62118 165864 62174 166664
rect 63130 165864 63186 166664
rect 64050 165864 64106 166664
rect 65062 165864 65118 166664
rect 66074 165864 66130 166664
rect 66994 165864 67050 166664
rect 68006 165864 68062 166664
rect 69018 165864 69074 166664
rect 69938 165864 69994 166664
rect 70950 165864 71006 166664
rect 71870 165864 71926 166664
rect 72882 165864 72938 166664
rect 73894 165864 73950 166664
rect 74814 165864 74870 166664
rect 75826 165864 75882 166664
rect 76838 165864 76894 166664
rect 77758 165864 77814 166664
rect 78770 165864 78826 166664
rect 79782 165864 79838 166664
rect 80702 165864 80758 166664
rect 81714 165864 81770 166664
rect 82726 165864 82782 166664
rect 83646 165864 83702 166664
rect 84658 165864 84714 166664
rect 85578 165864 85634 166664
rect 86590 165864 86646 166664
rect 87602 165864 87658 166664
rect 88522 165864 88578 166664
rect 89534 165864 89590 166664
rect 90546 165864 90602 166664
rect 91466 165864 91522 166664
rect 92478 165864 92534 166664
rect 93490 165864 93546 166664
rect 94410 165864 94466 166664
rect 95422 165864 95478 166664
rect 96434 165864 96490 166664
rect 97354 165864 97410 166664
rect 98366 165864 98422 166664
rect 99286 165864 99342 166664
rect 100298 165864 100354 166664
rect 101310 165864 101366 166664
rect 102230 165864 102286 166664
rect 103242 165864 103298 166664
rect 104254 165864 104310 166664
rect 105174 165864 105230 166664
rect 106186 165864 106242 166664
rect 107198 165864 107254 166664
rect 108118 165864 108174 166664
rect 109130 165864 109186 166664
rect 110142 165864 110198 166664
rect 111062 165864 111118 166664
rect 112074 165864 112130 166664
rect 112994 165864 113050 166664
rect 114006 165864 114062 166664
rect 115018 165864 115074 166664
rect 115938 165864 115994 166664
rect 116950 165864 117006 166664
rect 117962 165864 118018 166664
rect 118882 165864 118938 166664
rect 119894 165864 119950 166664
rect 120906 165864 120962 166664
rect 121826 165864 121882 166664
rect 122838 165864 122894 166664
rect 123850 165864 123906 166664
rect 124770 165864 124826 166664
rect 125782 165864 125838 166664
rect 126702 165864 126758 166664
rect 127714 165864 127770 166664
rect 128726 165864 128782 166664
rect 129646 165864 129702 166664
rect 130658 165864 130714 166664
rect 131670 165864 131726 166664
rect 132590 165864 132646 166664
rect 133602 165864 133658 166664
rect 134614 165864 134670 166664
rect 135534 165864 135590 166664
rect 136546 165864 136602 166664
rect 137558 165864 137614 166664
rect 138478 165864 138534 166664
rect 139490 165864 139546 166664
rect 140410 165864 140466 166664
rect 141422 165864 141478 166664
rect 142434 165864 142490 166664
rect 143354 165864 143410 166664
rect 144366 165864 144422 166664
rect 145378 165864 145434 166664
rect 146298 165864 146354 166664
rect 147310 165864 147366 166664
rect 148322 165864 148378 166664
rect 149242 165864 149298 166664
rect 150254 165864 150310 166664
rect 151266 165864 151322 166664
rect 152186 165864 152242 166664
rect 153198 165864 153254 166664
rect 154118 165864 154174 166664
rect 155130 165864 155186 166664
rect 156142 165864 156198 166664
rect 157062 165864 157118 166664
rect 158074 165864 158130 166664
rect 159086 165864 159142 166664
rect 160006 165864 160062 166664
rect 161018 165864 161074 166664
rect 162030 165864 162086 166664
rect 162950 165864 163006 166664
rect 163962 165864 164018 166664
rect 478 0 534 800
rect 1398 0 1454 800
rect 2318 0 2374 800
rect 3330 0 3386 800
rect 4250 0 4306 800
rect 5170 0 5226 800
rect 6182 0 6238 800
rect 7102 0 7158 800
rect 8114 0 8170 800
rect 9034 0 9090 800
rect 9954 0 10010 800
rect 10966 0 11022 800
rect 11886 0 11942 800
rect 12898 0 12954 800
rect 13818 0 13874 800
rect 14738 0 14794 800
rect 15750 0 15806 800
rect 16670 0 16726 800
rect 17682 0 17738 800
rect 18602 0 18658 800
rect 19522 0 19578 800
rect 20534 0 20590 800
rect 21454 0 21510 800
rect 22466 0 22522 800
rect 23386 0 23442 800
rect 24306 0 24362 800
rect 25318 0 25374 800
rect 26238 0 26294 800
rect 27250 0 27306 800
rect 28170 0 28226 800
rect 29090 0 29146 800
rect 30102 0 30158 800
rect 31022 0 31078 800
rect 32034 0 32090 800
rect 32954 0 33010 800
rect 33874 0 33930 800
rect 34886 0 34942 800
rect 35806 0 35862 800
rect 36818 0 36874 800
rect 37738 0 37794 800
rect 38658 0 38714 800
rect 39670 0 39726 800
rect 40590 0 40646 800
rect 41602 0 41658 800
rect 42522 0 42578 800
rect 43442 0 43498 800
rect 44454 0 44510 800
rect 45374 0 45430 800
rect 46294 0 46350 800
rect 47306 0 47362 800
rect 48226 0 48282 800
rect 49238 0 49294 800
rect 50158 0 50214 800
rect 51078 0 51134 800
rect 52090 0 52146 800
rect 53010 0 53066 800
rect 54022 0 54078 800
rect 54942 0 54998 800
rect 55862 0 55918 800
rect 56874 0 56930 800
rect 57794 0 57850 800
rect 58806 0 58862 800
rect 59726 0 59782 800
rect 60646 0 60702 800
rect 61658 0 61714 800
rect 62578 0 62634 800
rect 63590 0 63646 800
rect 64510 0 64566 800
rect 65430 0 65486 800
rect 66442 0 66498 800
rect 67362 0 67418 800
rect 68374 0 68430 800
rect 69294 0 69350 800
rect 70214 0 70270 800
rect 71226 0 71282 800
rect 72146 0 72202 800
rect 73158 0 73214 800
rect 74078 0 74134 800
rect 74998 0 75054 800
rect 76010 0 76066 800
rect 76930 0 76986 800
rect 77942 0 77998 800
rect 78862 0 78918 800
rect 79782 0 79838 800
rect 80794 0 80850 800
rect 81714 0 81770 800
rect 82726 0 82782 800
rect 83646 0 83702 800
rect 84566 0 84622 800
rect 85578 0 85634 800
rect 86498 0 86554 800
rect 87418 0 87474 800
rect 88430 0 88486 800
rect 89350 0 89406 800
rect 90362 0 90418 800
rect 91282 0 91338 800
rect 92202 0 92258 800
rect 93214 0 93270 800
rect 94134 0 94190 800
rect 95146 0 95202 800
rect 96066 0 96122 800
rect 96986 0 97042 800
rect 97998 0 98054 800
rect 98918 0 98974 800
rect 99930 0 99986 800
rect 100850 0 100906 800
rect 101770 0 101826 800
rect 102782 0 102838 800
rect 103702 0 103758 800
rect 104714 0 104770 800
rect 105634 0 105690 800
rect 106554 0 106610 800
rect 107566 0 107622 800
rect 108486 0 108542 800
rect 109498 0 109554 800
rect 110418 0 110474 800
rect 111338 0 111394 800
rect 112350 0 112406 800
rect 113270 0 113326 800
rect 114282 0 114338 800
rect 115202 0 115258 800
rect 116122 0 116178 800
rect 117134 0 117190 800
rect 118054 0 118110 800
rect 119066 0 119122 800
rect 119986 0 120042 800
rect 120906 0 120962 800
rect 121918 0 121974 800
rect 122838 0 122894 800
rect 123850 0 123906 800
rect 124770 0 124826 800
rect 125690 0 125746 800
rect 126702 0 126758 800
rect 127622 0 127678 800
rect 128542 0 128598 800
rect 129554 0 129610 800
rect 130474 0 130530 800
rect 131486 0 131542 800
rect 132406 0 132462 800
rect 133326 0 133382 800
rect 134338 0 134394 800
rect 135258 0 135314 800
rect 136270 0 136326 800
rect 137190 0 137246 800
rect 138110 0 138166 800
rect 139122 0 139178 800
rect 140042 0 140098 800
rect 141054 0 141110 800
rect 141974 0 142030 800
rect 142894 0 142950 800
rect 143906 0 143962 800
rect 144826 0 144882 800
rect 145838 0 145894 800
rect 146758 0 146814 800
rect 147678 0 147734 800
rect 148690 0 148746 800
rect 149610 0 149666 800
rect 150622 0 150678 800
rect 151542 0 151598 800
rect 152462 0 152518 800
rect 153474 0 153530 800
rect 154394 0 154450 800
rect 155406 0 155462 800
rect 156326 0 156382 800
rect 157246 0 157302 800
rect 158258 0 158314 800
rect 159178 0 159234 800
rect 160190 0 160246 800
rect 161110 0 161166 800
rect 162030 0 162086 800
rect 163042 0 163098 800
rect 163962 0 164018 800
<< obsm2 >>
rect 20 165808 422 166002
rect 590 165808 1342 166002
rect 1510 165808 2354 166002
rect 2522 165808 3274 166002
rect 3442 165808 4286 166002
rect 4454 165808 5298 166002
rect 5466 165808 6218 166002
rect 6386 165808 7230 166002
rect 7398 165808 8242 166002
rect 8410 165808 9162 166002
rect 9330 165808 10174 166002
rect 10342 165808 11186 166002
rect 11354 165808 12106 166002
rect 12274 165808 13118 166002
rect 13286 165808 14130 166002
rect 14298 165808 15050 166002
rect 15218 165808 16062 166002
rect 16230 165808 16982 166002
rect 17150 165808 17994 166002
rect 18162 165808 19006 166002
rect 19174 165808 19926 166002
rect 20094 165808 20938 166002
rect 21106 165808 21950 166002
rect 22118 165808 22870 166002
rect 23038 165808 23882 166002
rect 24050 165808 24894 166002
rect 25062 165808 25814 166002
rect 25982 165808 26826 166002
rect 26994 165808 27838 166002
rect 28006 165808 28758 166002
rect 28926 165808 29770 166002
rect 29938 165808 30690 166002
rect 30858 165808 31702 166002
rect 31870 165808 32714 166002
rect 32882 165808 33634 166002
rect 33802 165808 34646 166002
rect 34814 165808 35658 166002
rect 35826 165808 36578 166002
rect 36746 165808 37590 166002
rect 37758 165808 38602 166002
rect 38770 165808 39522 166002
rect 39690 165808 40534 166002
rect 40702 165808 41546 166002
rect 41714 165808 42466 166002
rect 42634 165808 43478 166002
rect 43646 165808 44398 166002
rect 44566 165808 45410 166002
rect 45578 165808 46422 166002
rect 46590 165808 47342 166002
rect 47510 165808 48354 166002
rect 48522 165808 49366 166002
rect 49534 165808 50286 166002
rect 50454 165808 51298 166002
rect 51466 165808 52310 166002
rect 52478 165808 53230 166002
rect 53398 165808 54242 166002
rect 54410 165808 55254 166002
rect 55422 165808 56174 166002
rect 56342 165808 57186 166002
rect 57354 165808 58106 166002
rect 58274 165808 59118 166002
rect 59286 165808 60130 166002
rect 60298 165808 61050 166002
rect 61218 165808 62062 166002
rect 62230 165808 63074 166002
rect 63242 165808 63994 166002
rect 64162 165808 65006 166002
rect 65174 165808 66018 166002
rect 66186 165808 66938 166002
rect 67106 165808 67950 166002
rect 68118 165808 68962 166002
rect 69130 165808 69882 166002
rect 70050 165808 70894 166002
rect 71062 165808 71814 166002
rect 71982 165808 72826 166002
rect 72994 165808 73838 166002
rect 74006 165808 74758 166002
rect 74926 165808 75770 166002
rect 75938 165808 76782 166002
rect 76950 165808 77702 166002
rect 77870 165808 78714 166002
rect 78882 165808 79726 166002
rect 79894 165808 80646 166002
rect 80814 165808 81658 166002
rect 81826 165808 82670 166002
rect 82838 165808 83590 166002
rect 83758 165808 84602 166002
rect 84770 165808 85522 166002
rect 85690 165808 86534 166002
rect 86702 165808 87546 166002
rect 87714 165808 88466 166002
rect 88634 165808 89478 166002
rect 89646 165808 90490 166002
rect 90658 165808 91410 166002
rect 91578 165808 92422 166002
rect 92590 165808 93434 166002
rect 93602 165808 94354 166002
rect 94522 165808 95366 166002
rect 95534 165808 96378 166002
rect 96546 165808 97298 166002
rect 97466 165808 98310 166002
rect 98478 165808 99230 166002
rect 99398 165808 100242 166002
rect 100410 165808 101254 166002
rect 101422 165808 102174 166002
rect 102342 165808 103186 166002
rect 103354 165808 104198 166002
rect 104366 165808 105118 166002
rect 105286 165808 106130 166002
rect 106298 165808 107142 166002
rect 107310 165808 108062 166002
rect 108230 165808 109074 166002
rect 109242 165808 110086 166002
rect 110254 165808 111006 166002
rect 111174 165808 112018 166002
rect 112186 165808 112938 166002
rect 113106 165808 113950 166002
rect 114118 165808 114962 166002
rect 115130 165808 115882 166002
rect 116050 165808 116894 166002
rect 117062 165808 117906 166002
rect 118074 165808 118826 166002
rect 118994 165808 119838 166002
rect 120006 165808 120850 166002
rect 121018 165808 121770 166002
rect 121938 165808 122782 166002
rect 122950 165808 123794 166002
rect 123962 165808 124714 166002
rect 124882 165808 125726 166002
rect 125894 165808 126646 166002
rect 126814 165808 127658 166002
rect 127826 165808 128670 166002
rect 128838 165808 129590 166002
rect 129758 165808 130602 166002
rect 130770 165808 131614 166002
rect 131782 165808 132534 166002
rect 132702 165808 133546 166002
rect 133714 165808 134558 166002
rect 134726 165808 135478 166002
rect 135646 165808 136490 166002
rect 136658 165808 137502 166002
rect 137670 165808 138422 166002
rect 138590 165808 139434 166002
rect 139602 165808 140354 166002
rect 140522 165808 141366 166002
rect 141534 165808 142378 166002
rect 142546 165808 143298 166002
rect 143466 165808 144310 166002
rect 144478 165808 145322 166002
rect 145490 165808 146242 166002
rect 146410 165808 147254 166002
rect 147422 165808 148266 166002
rect 148434 165808 149186 166002
rect 149354 165808 150198 166002
rect 150366 165808 151210 166002
rect 151378 165808 152130 166002
rect 152298 165808 153142 166002
rect 153310 165808 154062 166002
rect 154230 165808 155074 166002
rect 155242 165808 156086 166002
rect 156254 165808 157006 166002
rect 157174 165808 158018 166002
rect 158186 165808 159030 166002
rect 159198 165808 159950 166002
rect 160118 165808 160962 166002
rect 161130 165808 161974 166002
rect 162142 165808 162894 166002
rect 163062 165808 163906 166002
rect 164074 165808 164478 166002
rect 20 856 164478 165808
rect 20 2 422 856
rect 590 2 1342 856
rect 1510 2 2262 856
rect 2430 2 3274 856
rect 3442 2 4194 856
rect 4362 2 5114 856
rect 5282 2 6126 856
rect 6294 2 7046 856
rect 7214 2 8058 856
rect 8226 2 8978 856
rect 9146 2 9898 856
rect 10066 2 10910 856
rect 11078 2 11830 856
rect 11998 2 12842 856
rect 13010 2 13762 856
rect 13930 2 14682 856
rect 14850 2 15694 856
rect 15862 2 16614 856
rect 16782 2 17626 856
rect 17794 2 18546 856
rect 18714 2 19466 856
rect 19634 2 20478 856
rect 20646 2 21398 856
rect 21566 2 22410 856
rect 22578 2 23330 856
rect 23498 2 24250 856
rect 24418 2 25262 856
rect 25430 2 26182 856
rect 26350 2 27194 856
rect 27362 2 28114 856
rect 28282 2 29034 856
rect 29202 2 30046 856
rect 30214 2 30966 856
rect 31134 2 31978 856
rect 32146 2 32898 856
rect 33066 2 33818 856
rect 33986 2 34830 856
rect 34998 2 35750 856
rect 35918 2 36762 856
rect 36930 2 37682 856
rect 37850 2 38602 856
rect 38770 2 39614 856
rect 39782 2 40534 856
rect 40702 2 41546 856
rect 41714 2 42466 856
rect 42634 2 43386 856
rect 43554 2 44398 856
rect 44566 2 45318 856
rect 45486 2 46238 856
rect 46406 2 47250 856
rect 47418 2 48170 856
rect 48338 2 49182 856
rect 49350 2 50102 856
rect 50270 2 51022 856
rect 51190 2 52034 856
rect 52202 2 52954 856
rect 53122 2 53966 856
rect 54134 2 54886 856
rect 55054 2 55806 856
rect 55974 2 56818 856
rect 56986 2 57738 856
rect 57906 2 58750 856
rect 58918 2 59670 856
rect 59838 2 60590 856
rect 60758 2 61602 856
rect 61770 2 62522 856
rect 62690 2 63534 856
rect 63702 2 64454 856
rect 64622 2 65374 856
rect 65542 2 66386 856
rect 66554 2 67306 856
rect 67474 2 68318 856
rect 68486 2 69238 856
rect 69406 2 70158 856
rect 70326 2 71170 856
rect 71338 2 72090 856
rect 72258 2 73102 856
rect 73270 2 74022 856
rect 74190 2 74942 856
rect 75110 2 75954 856
rect 76122 2 76874 856
rect 77042 2 77886 856
rect 78054 2 78806 856
rect 78974 2 79726 856
rect 79894 2 80738 856
rect 80906 2 81658 856
rect 81826 2 82670 856
rect 82838 2 83590 856
rect 83758 2 84510 856
rect 84678 2 85522 856
rect 85690 2 86442 856
rect 86610 2 87362 856
rect 87530 2 88374 856
rect 88542 2 89294 856
rect 89462 2 90306 856
rect 90474 2 91226 856
rect 91394 2 92146 856
rect 92314 2 93158 856
rect 93326 2 94078 856
rect 94246 2 95090 856
rect 95258 2 96010 856
rect 96178 2 96930 856
rect 97098 2 97942 856
rect 98110 2 98862 856
rect 99030 2 99874 856
rect 100042 2 100794 856
rect 100962 2 101714 856
rect 101882 2 102726 856
rect 102894 2 103646 856
rect 103814 2 104658 856
rect 104826 2 105578 856
rect 105746 2 106498 856
rect 106666 2 107510 856
rect 107678 2 108430 856
rect 108598 2 109442 856
rect 109610 2 110362 856
rect 110530 2 111282 856
rect 111450 2 112294 856
rect 112462 2 113214 856
rect 113382 2 114226 856
rect 114394 2 115146 856
rect 115314 2 116066 856
rect 116234 2 117078 856
rect 117246 2 117998 856
rect 118166 2 119010 856
rect 119178 2 119930 856
rect 120098 2 120850 856
rect 121018 2 121862 856
rect 122030 2 122782 856
rect 122950 2 123794 856
rect 123962 2 124714 856
rect 124882 2 125634 856
rect 125802 2 126646 856
rect 126814 2 127566 856
rect 127734 2 128486 856
rect 128654 2 129498 856
rect 129666 2 130418 856
rect 130586 2 131430 856
rect 131598 2 132350 856
rect 132518 2 133270 856
rect 133438 2 134282 856
rect 134450 2 135202 856
rect 135370 2 136214 856
rect 136382 2 137134 856
rect 137302 2 138054 856
rect 138222 2 139066 856
rect 139234 2 139986 856
rect 140154 2 140998 856
rect 141166 2 141918 856
rect 142086 2 142838 856
rect 143006 2 143850 856
rect 144018 2 144770 856
rect 144938 2 145782 856
rect 145950 2 146702 856
rect 146870 2 147622 856
rect 147790 2 148634 856
rect 148802 2 149554 856
rect 149722 2 150566 856
rect 150734 2 151486 856
rect 151654 2 152406 856
rect 152574 2 153418 856
rect 153586 2 154338 856
rect 154506 2 155350 856
rect 155518 2 156270 856
rect 156438 2 157190 856
rect 157358 2 158202 856
rect 158370 2 159122 856
rect 159290 2 160134 856
rect 160302 2 161054 856
rect 161222 2 161974 856
rect 162142 2 162986 856
rect 163154 2 163906 856
rect 164074 2 164478 856
<< metal3 >>
rect 0 165248 800 165368
rect 163720 165112 164520 165232
rect 0 162664 800 162784
rect 163720 162392 164520 162512
rect 0 160080 800 160200
rect 163720 159536 164520 159656
rect 0 157496 800 157616
rect 163720 156816 164520 156936
rect 0 154912 800 155032
rect 163720 153960 164520 154080
rect 0 152328 800 152448
rect 163720 151240 164520 151360
rect 0 149880 800 150000
rect 163720 148520 164520 148640
rect 0 147296 800 147416
rect 163720 145664 164520 145784
rect 0 144712 800 144832
rect 163720 142944 164520 143064
rect 0 142128 800 142248
rect 163720 140088 164520 140208
rect 0 139544 800 139664
rect 163720 137368 164520 137488
rect 0 136960 800 137080
rect 0 134512 800 134632
rect 163720 134648 164520 134768
rect 0 131928 800 132048
rect 163720 131792 164520 131912
rect 0 129344 800 129464
rect 163720 129072 164520 129192
rect 0 126760 800 126880
rect 163720 126216 164520 126336
rect 0 124176 800 124296
rect 163720 123496 164520 123616
rect 0 121592 800 121712
rect 163720 120640 164520 120760
rect 0 119008 800 119128
rect 163720 117920 164520 118040
rect 0 116560 800 116680
rect 163720 115200 164520 115320
rect 0 113976 800 114096
rect 163720 112344 164520 112464
rect 0 111392 800 111512
rect 163720 109624 164520 109744
rect 0 108808 800 108928
rect 163720 106768 164520 106888
rect 0 106224 800 106344
rect 163720 104048 164520 104168
rect 0 103640 800 103760
rect 0 101192 800 101312
rect 163720 101328 164520 101448
rect 0 98608 800 98728
rect 163720 98472 164520 98592
rect 0 96024 800 96144
rect 163720 95752 164520 95872
rect 0 93440 800 93560
rect 163720 92896 164520 93016
rect 0 90856 800 90976
rect 163720 90176 164520 90296
rect 0 88272 800 88392
rect 163720 87320 164520 87440
rect 0 85688 800 85808
rect 163720 84600 164520 84720
rect 0 83240 800 83360
rect 163720 81880 164520 82000
rect 0 80656 800 80776
rect 163720 79024 164520 79144
rect 0 78072 800 78192
rect 163720 76304 164520 76424
rect 0 75488 800 75608
rect 163720 73448 164520 73568
rect 0 72904 800 73024
rect 163720 70728 164520 70848
rect 0 70320 800 70440
rect 0 67872 800 67992
rect 163720 68008 164520 68128
rect 0 65288 800 65408
rect 163720 65152 164520 65272
rect 0 62704 800 62824
rect 163720 62432 164520 62552
rect 0 60120 800 60240
rect 163720 59576 164520 59696
rect 0 57536 800 57656
rect 163720 56856 164520 56976
rect 0 54952 800 55072
rect 163720 54000 164520 54120
rect 0 52368 800 52488
rect 163720 51280 164520 51400
rect 0 49920 800 50040
rect 163720 48560 164520 48680
rect 0 47336 800 47456
rect 163720 45704 164520 45824
rect 0 44752 800 44872
rect 163720 42984 164520 43104
rect 0 42168 800 42288
rect 163720 40128 164520 40248
rect 0 39584 800 39704
rect 163720 37408 164520 37528
rect 0 37000 800 37120
rect 0 34552 800 34672
rect 163720 34688 164520 34808
rect 0 31968 800 32088
rect 163720 31832 164520 31952
rect 0 29384 800 29504
rect 163720 29112 164520 29232
rect 0 26800 800 26920
rect 163720 26256 164520 26376
rect 0 24216 800 24336
rect 163720 23536 164520 23656
rect 0 21632 800 21752
rect 163720 20680 164520 20800
rect 0 19048 800 19168
rect 163720 17960 164520 18080
rect 0 16600 800 16720
rect 163720 15240 164520 15360
rect 0 14016 800 14136
rect 163720 12384 164520 12504
rect 0 11432 800 11552
rect 163720 9664 164520 9784
rect 0 8848 800 8968
rect 163720 6808 164520 6928
rect 0 6264 800 6384
rect 163720 4088 164520 4208
rect 0 3680 800 3800
rect 0 1232 800 1352
rect 163720 1368 164520 1488
<< obsm3 >>
rect 800 162864 164483 164321
rect 880 162592 164483 162864
rect 880 162584 163640 162592
rect 800 162312 163640 162584
rect 800 160280 164483 162312
rect 880 160000 164483 160280
rect 800 159736 164483 160000
rect 800 159456 163640 159736
rect 800 157696 164483 159456
rect 880 157416 164483 157696
rect 800 157016 164483 157416
rect 800 156736 163640 157016
rect 800 155112 164483 156736
rect 880 154832 164483 155112
rect 800 154160 164483 154832
rect 800 153880 163640 154160
rect 800 152528 164483 153880
rect 880 152248 164483 152528
rect 800 151440 164483 152248
rect 800 151160 163640 151440
rect 800 150080 164483 151160
rect 880 149800 164483 150080
rect 800 148720 164483 149800
rect 800 148440 163640 148720
rect 800 147496 164483 148440
rect 880 147216 164483 147496
rect 800 145864 164483 147216
rect 800 145584 163640 145864
rect 800 144912 164483 145584
rect 880 144632 164483 144912
rect 800 143144 164483 144632
rect 800 142864 163640 143144
rect 800 142328 164483 142864
rect 880 142048 164483 142328
rect 800 140288 164483 142048
rect 800 140008 163640 140288
rect 800 139744 164483 140008
rect 880 139464 164483 139744
rect 800 137568 164483 139464
rect 800 137288 163640 137568
rect 800 137160 164483 137288
rect 880 136880 164483 137160
rect 800 134848 164483 136880
rect 800 134712 163640 134848
rect 880 134568 163640 134712
rect 880 134432 164483 134568
rect 800 132128 164483 134432
rect 880 131992 164483 132128
rect 880 131848 163640 131992
rect 800 131712 163640 131848
rect 800 129544 164483 131712
rect 880 129272 164483 129544
rect 880 129264 163640 129272
rect 800 128992 163640 129264
rect 800 126960 164483 128992
rect 880 126680 164483 126960
rect 800 126416 164483 126680
rect 800 126136 163640 126416
rect 800 124376 164483 126136
rect 880 124096 164483 124376
rect 800 123696 164483 124096
rect 800 123416 163640 123696
rect 800 121792 164483 123416
rect 880 121512 164483 121792
rect 800 120840 164483 121512
rect 800 120560 163640 120840
rect 800 119208 164483 120560
rect 880 118928 164483 119208
rect 800 118120 164483 118928
rect 800 117840 163640 118120
rect 800 116760 164483 117840
rect 880 116480 164483 116760
rect 800 115400 164483 116480
rect 800 115120 163640 115400
rect 800 114176 164483 115120
rect 880 113896 164483 114176
rect 800 112544 164483 113896
rect 800 112264 163640 112544
rect 800 111592 164483 112264
rect 880 111312 164483 111592
rect 800 109824 164483 111312
rect 800 109544 163640 109824
rect 800 109008 164483 109544
rect 880 108728 164483 109008
rect 800 106968 164483 108728
rect 800 106688 163640 106968
rect 800 106424 164483 106688
rect 880 106144 164483 106424
rect 800 104248 164483 106144
rect 800 103968 163640 104248
rect 800 103840 164483 103968
rect 880 103560 164483 103840
rect 800 101528 164483 103560
rect 800 101392 163640 101528
rect 880 101248 163640 101392
rect 880 101112 164483 101248
rect 800 98808 164483 101112
rect 880 98672 164483 98808
rect 880 98528 163640 98672
rect 800 98392 163640 98528
rect 800 96224 164483 98392
rect 880 95952 164483 96224
rect 880 95944 163640 95952
rect 800 95672 163640 95944
rect 800 93640 164483 95672
rect 880 93360 164483 93640
rect 800 93096 164483 93360
rect 800 92816 163640 93096
rect 800 91056 164483 92816
rect 880 90776 164483 91056
rect 800 90376 164483 90776
rect 800 90096 163640 90376
rect 800 88472 164483 90096
rect 880 88192 164483 88472
rect 800 87520 164483 88192
rect 800 87240 163640 87520
rect 800 85888 164483 87240
rect 880 85608 164483 85888
rect 800 84800 164483 85608
rect 800 84520 163640 84800
rect 800 83440 164483 84520
rect 880 83160 164483 83440
rect 800 82080 164483 83160
rect 800 81800 163640 82080
rect 800 80856 164483 81800
rect 880 80576 164483 80856
rect 800 79224 164483 80576
rect 800 78944 163640 79224
rect 800 78272 164483 78944
rect 880 77992 164483 78272
rect 800 76504 164483 77992
rect 800 76224 163640 76504
rect 800 75688 164483 76224
rect 880 75408 164483 75688
rect 800 73648 164483 75408
rect 800 73368 163640 73648
rect 800 73104 164483 73368
rect 880 72824 164483 73104
rect 800 70928 164483 72824
rect 800 70648 163640 70928
rect 800 70520 164483 70648
rect 880 70240 164483 70520
rect 800 68208 164483 70240
rect 800 68072 163640 68208
rect 880 67928 163640 68072
rect 880 67792 164483 67928
rect 800 65488 164483 67792
rect 880 65352 164483 65488
rect 880 65208 163640 65352
rect 800 65072 163640 65208
rect 800 62904 164483 65072
rect 880 62632 164483 62904
rect 880 62624 163640 62632
rect 800 62352 163640 62624
rect 800 60320 164483 62352
rect 880 60040 164483 60320
rect 800 59776 164483 60040
rect 800 59496 163640 59776
rect 800 57736 164483 59496
rect 880 57456 164483 57736
rect 800 57056 164483 57456
rect 800 56776 163640 57056
rect 800 55152 164483 56776
rect 880 54872 164483 55152
rect 800 54200 164483 54872
rect 800 53920 163640 54200
rect 800 52568 164483 53920
rect 880 52288 164483 52568
rect 800 51480 164483 52288
rect 800 51200 163640 51480
rect 800 50120 164483 51200
rect 880 49840 164483 50120
rect 800 48760 164483 49840
rect 800 48480 163640 48760
rect 800 47536 164483 48480
rect 880 47256 164483 47536
rect 800 45904 164483 47256
rect 800 45624 163640 45904
rect 800 44952 164483 45624
rect 880 44672 164483 44952
rect 800 43184 164483 44672
rect 800 42904 163640 43184
rect 800 42368 164483 42904
rect 880 42088 164483 42368
rect 800 40328 164483 42088
rect 800 40048 163640 40328
rect 800 39784 164483 40048
rect 880 39504 164483 39784
rect 800 37608 164483 39504
rect 800 37328 163640 37608
rect 800 37200 164483 37328
rect 880 36920 164483 37200
rect 800 34888 164483 36920
rect 800 34752 163640 34888
rect 880 34608 163640 34752
rect 880 34472 164483 34608
rect 800 32168 164483 34472
rect 880 32032 164483 32168
rect 880 31888 163640 32032
rect 800 31752 163640 31888
rect 800 29584 164483 31752
rect 880 29312 164483 29584
rect 880 29304 163640 29312
rect 800 29032 163640 29304
rect 800 27000 164483 29032
rect 880 26720 164483 27000
rect 800 26456 164483 26720
rect 800 26176 163640 26456
rect 800 24416 164483 26176
rect 880 24136 164483 24416
rect 800 23736 164483 24136
rect 800 23456 163640 23736
rect 800 21832 164483 23456
rect 880 21552 164483 21832
rect 800 20880 164483 21552
rect 800 20600 163640 20880
rect 800 19248 164483 20600
rect 880 18968 164483 19248
rect 800 18160 164483 18968
rect 800 17880 163640 18160
rect 800 16800 164483 17880
rect 880 16520 164483 16800
rect 800 15440 164483 16520
rect 800 15160 163640 15440
rect 800 14216 164483 15160
rect 880 13936 164483 14216
rect 800 12584 164483 13936
rect 800 12304 163640 12584
rect 800 11632 164483 12304
rect 880 11352 164483 11632
rect 800 9864 164483 11352
rect 800 9584 163640 9864
rect 800 9048 164483 9584
rect 880 8768 164483 9048
rect 800 7008 164483 8768
rect 800 6728 163640 7008
rect 800 6464 164483 6728
rect 880 6184 164483 6464
rect 800 4288 164483 6184
rect 800 4008 163640 4288
rect 800 3880 164483 4008
rect 880 3600 164483 3880
rect 800 1568 164483 3600
rect 800 1432 163640 1568
rect 880 1288 163640 1432
rect 880 1152 164483 1288
rect 800 443 164483 1152
<< metal4 >>
rect 4208 2128 4528 164336
rect 19568 2128 19888 164336
rect 34928 2128 35248 164336
rect 50288 2128 50608 164336
rect 65648 2128 65968 164336
rect 81008 2128 81328 164336
rect 96368 2128 96688 164336
rect 111728 2128 112048 164336
rect 127088 2128 127408 164336
rect 142448 2128 142768 164336
rect 157808 2128 158128 164336
<< obsm4 >>
rect 4659 2048 19488 164117
rect 19968 2048 34848 164117
rect 35328 2048 50208 164117
rect 50688 2048 65568 164117
rect 66048 2048 80928 164117
rect 81408 2048 96288 164117
rect 96768 2048 111648 164117
rect 112128 2048 127008 164117
rect 127488 2048 142368 164117
rect 142848 2048 157728 164117
rect 158208 2048 163517 164117
rect 4659 443 163517 2048
<< labels >>
rlabel metal2 s 107566 0 107622 800 6 i_dout0[0]
port 1 nsew signal input
rlabel metal3 s 0 72904 800 73024 6 i_dout0[10]
port 2 nsew signal input
rlabel metal3 s 0 80656 800 80776 6 i_dout0[11]
port 3 nsew signal input
rlabel metal2 s 133602 165864 133658 166664 6 i_dout0[12]
port 4 nsew signal input
rlabel metal2 s 136546 165864 136602 166664 6 i_dout0[13]
port 5 nsew signal input
rlabel metal3 s 0 93440 800 93560 6 i_dout0[14]
port 6 nsew signal input
rlabel metal3 s 0 98608 800 98728 6 i_dout0[15]
port 7 nsew signal input
rlabel metal2 s 141422 165864 141478 166664 6 i_dout0[16]
port 8 nsew signal input
rlabel metal3 s 0 111392 800 111512 6 i_dout0[17]
port 9 nsew signal input
rlabel metal2 s 144826 0 144882 800 6 i_dout0[18]
port 10 nsew signal input
rlabel metal2 s 146298 165864 146354 166664 6 i_dout0[19]
port 11 nsew signal input
rlabel metal2 s 115938 165864 115994 166664 6 i_dout0[1]
port 12 nsew signal input
rlabel metal3 s 163720 129072 164520 129192 6 i_dout0[20]
port 13 nsew signal input
rlabel metal3 s 0 121592 800 121712 6 i_dout0[21]
port 14 nsew signal input
rlabel metal2 s 150622 0 150678 800 6 i_dout0[22]
port 15 nsew signal input
rlabel metal3 s 163720 137368 164520 137488 6 i_dout0[23]
port 16 nsew signal input
rlabel metal2 s 152186 165864 152242 166664 6 i_dout0[24]
port 17 nsew signal input
rlabel metal3 s 163720 148520 164520 148640 6 i_dout0[25]
port 18 nsew signal input
rlabel metal2 s 154394 0 154450 800 6 i_dout0[26]
port 19 nsew signal input
rlabel metal3 s 0 147296 800 147416 6 i_dout0[27]
port 20 nsew signal input
rlabel metal3 s 0 152328 800 152448 6 i_dout0[28]
port 21 nsew signal input
rlabel metal2 s 161110 0 161166 800 6 i_dout0[29]
port 22 nsew signal input
rlabel metal2 s 113270 0 113326 800 6 i_dout0[2]
port 23 nsew signal input
rlabel metal3 s 163720 159536 164520 159656 6 i_dout0[30]
port 24 nsew signal input
rlabel metal3 s 0 165248 800 165368 6 i_dout0[31]
port 25 nsew signal input
rlabel metal2 s 117134 0 117190 800 6 i_dout0[3]
port 26 nsew signal input
rlabel metal3 s 163720 42984 164520 43104 6 i_dout0[4]
port 27 nsew signal input
rlabel metal3 s 163720 54000 164520 54120 6 i_dout0[5]
port 28 nsew signal input
rlabel metal3 s 163720 62432 164520 62552 6 i_dout0[6]
port 29 nsew signal input
rlabel metal2 s 127622 0 127678 800 6 i_dout0[7]
port 30 nsew signal input
rlabel metal3 s 163720 73448 164520 73568 6 i_dout0[8]
port 31 nsew signal input
rlabel metal2 s 131670 165864 131726 166664 6 i_dout0[9]
port 32 nsew signal input
rlabel metal2 s 108486 0 108542 800 6 i_dout0_1[0]
port 33 nsew signal input
rlabel metal3 s 0 67872 800 67992 6 i_dout0_1[10]
port 34 nsew signal input
rlabel metal3 s 0 75488 800 75608 6 i_dout0_1[11]
port 35 nsew signal input
rlabel metal3 s 163720 92896 164520 93016 6 i_dout0_1[12]
port 36 nsew signal input
rlabel metal2 s 134614 165864 134670 166664 6 i_dout0_1[13]
port 37 nsew signal input
rlabel metal2 s 137558 165864 137614 166664 6 i_dout0_1[14]
port 38 nsew signal input
rlabel metal3 s 163720 104048 164520 104168 6 i_dout0_1[15]
port 39 nsew signal input
rlabel metal3 s 0 103640 800 103760 6 i_dout0_1[16]
port 40 nsew signal input
rlabel metal2 s 140042 0 140098 800 6 i_dout0_1[17]
port 41 nsew signal input
rlabel metal3 s 0 113976 800 114096 6 i_dout0_1[18]
port 42 nsew signal input
rlabel metal2 s 145378 165864 145434 166664 6 i_dout0_1[19]
port 43 nsew signal input
rlabel metal3 s 163720 9664 164520 9784 6 i_dout0_1[1]
port 44 nsew signal input
rlabel metal3 s 0 116560 800 116680 6 i_dout0_1[20]
port 45 nsew signal input
rlabel metal2 s 147310 165864 147366 166664 6 i_dout0_1[21]
port 46 nsew signal input
rlabel metal2 s 149242 165864 149298 166664 6 i_dout0_1[22]
port 47 nsew signal input
rlabel metal2 s 151266 165864 151322 166664 6 i_dout0_1[23]
port 48 nsew signal input
rlabel metal3 s 0 131928 800 132048 6 i_dout0_1[24]
port 49 nsew signal input
rlabel metal3 s 0 134512 800 134632 6 i_dout0_1[25]
port 50 nsew signal input
rlabel metal2 s 156142 165864 156198 166664 6 i_dout0_1[26]
port 51 nsew signal input
rlabel metal2 s 156326 0 156382 800 6 i_dout0_1[27]
port 52 nsew signal input
rlabel metal2 s 159086 165864 159142 166664 6 i_dout0_1[28]
port 53 nsew signal input
rlabel metal3 s 0 160080 800 160200 6 i_dout0_1[29]
port 54 nsew signal input
rlabel metal3 s 163720 17960 164520 18080 6 i_dout0_1[2]
port 55 nsew signal input
rlabel metal3 s 163720 156816 164520 156936 6 i_dout0_1[30]
port 56 nsew signal input
rlabel metal2 s 163042 0 163098 800 6 i_dout0_1[31]
port 57 nsew signal input
rlabel metal2 s 116122 0 116178 800 6 i_dout0_1[3]
port 58 nsew signal input
rlabel metal3 s 163720 37408 164520 37528 6 i_dout0_1[4]
port 59 nsew signal input
rlabel metal2 s 123850 165864 123906 166664 6 i_dout0_1[5]
port 60 nsew signal input
rlabel metal3 s 0 39584 800 39704 6 i_dout0_1[6]
port 61 nsew signal input
rlabel metal2 s 126702 0 126758 800 6 i_dout0_1[7]
port 62 nsew signal input
rlabel metal2 s 131486 0 131542 800 6 i_dout0_1[8]
port 63 nsew signal input
rlabel metal3 s 163720 81880 164520 82000 6 i_dout0_1[9]
port 64 nsew signal input
rlabel metal2 s 109498 0 109554 800 6 i_dout1[0]
port 65 nsew signal input
rlabel metal3 s 163720 87320 164520 87440 6 i_dout1[10]
port 66 nsew signal input
rlabel metal3 s 163720 90176 164520 90296 6 i_dout1[11]
port 67 nsew signal input
rlabel metal2 s 138110 0 138166 800 6 i_dout1[12]
port 68 nsew signal input
rlabel metal3 s 163720 95752 164520 95872 6 i_dout1[13]
port 69 nsew signal input
rlabel metal3 s 0 96024 800 96144 6 i_dout1[14]
port 70 nsew signal input
rlabel metal3 s 0 101192 800 101312 6 i_dout1[15]
port 71 nsew signal input
rlabel metal3 s 0 106224 800 106344 6 i_dout1[16]
port 72 nsew signal input
rlabel metal2 s 141974 0 142030 800 6 i_dout1[17]
port 73 nsew signal input
rlabel metal2 s 143354 165864 143410 166664 6 i_dout1[18]
port 74 nsew signal input
rlabel metal3 s 163720 120640 164520 120760 6 i_dout1[19]
port 75 nsew signal input
rlabel metal3 s 0 11432 800 11552 6 i_dout1[1]
port 76 nsew signal input
rlabel metal2 s 146758 0 146814 800 6 i_dout1[20]
port 77 nsew signal input
rlabel metal2 s 148322 165864 148378 166664 6 i_dout1[21]
port 78 nsew signal input
rlabel metal3 s 0 126760 800 126880 6 i_dout1[22]
port 79 nsew signal input
rlabel metal3 s 163720 140088 164520 140208 6 i_dout1[23]
port 80 nsew signal input
rlabel metal2 s 153198 165864 153254 166664 6 i_dout1[24]
port 81 nsew signal input
rlabel metal2 s 155130 165864 155186 166664 6 i_dout1[25]
port 82 nsew signal input
rlabel metal2 s 155406 0 155462 800 6 i_dout1[26]
port 83 nsew signal input
rlabel metal2 s 157246 0 157302 800 6 i_dout1[27]
port 84 nsew signal input
rlabel metal2 s 159178 0 159234 800 6 i_dout1[28]
port 85 nsew signal input
rlabel metal3 s 163720 153960 164520 154080 6 i_dout1[29]
port 86 nsew signal input
rlabel metal3 s 0 24216 800 24336 6 i_dout1[2]
port 87 nsew signal input
rlabel metal3 s 163720 162392 164520 162512 6 i_dout1[30]
port 88 nsew signal input
rlabel metal2 s 162950 165864 163006 166664 6 i_dout1[31]
port 89 nsew signal input
rlabel metal2 s 118054 0 118110 800 6 i_dout1[3]
port 90 nsew signal input
rlabel metal3 s 163720 45704 164520 45824 6 i_dout1[4]
port 91 nsew signal input
rlabel metal2 s 123850 0 123906 800 6 i_dout1[5]
port 92 nsew signal input
rlabel metal2 s 126702 165864 126758 166664 6 i_dout1[6]
port 93 nsew signal input
rlabel metal2 s 128542 0 128598 800 6 i_dout1[7]
port 94 nsew signal input
rlabel metal3 s 163720 76304 164520 76424 6 i_dout1[8]
port 95 nsew signal input
rlabel metal2 s 133326 0 133382 800 6 i_dout1[9]
port 96 nsew signal input
rlabel metal3 s 163720 1368 164520 1488 6 i_dout1_1[0]
port 97 nsew signal input
rlabel metal3 s 0 70320 800 70440 6 i_dout1_1[10]
port 98 nsew signal input
rlabel metal3 s 0 78072 800 78192 6 i_dout1_1[11]
port 99 nsew signal input
rlabel metal2 s 137190 0 137246 800 6 i_dout1_1[12]
port 100 nsew signal input
rlabel metal2 s 135534 165864 135590 166664 6 i_dout1_1[13]
port 101 nsew signal input
rlabel metal2 s 138478 165864 138534 166664 6 i_dout1_1[14]
port 102 nsew signal input
rlabel metal2 s 139490 165864 139546 166664 6 i_dout1_1[15]
port 103 nsew signal input
rlabel metal3 s 163720 109624 164520 109744 6 i_dout1_1[16]
port 104 nsew signal input
rlabel metal2 s 141054 0 141110 800 6 i_dout1_1[17]
port 105 nsew signal input
rlabel metal2 s 143906 0 143962 800 6 i_dout1_1[18]
port 106 nsew signal input
rlabel metal3 s 163720 117920 164520 118040 6 i_dout1_1[19]
port 107 nsew signal input
rlabel metal2 s 111338 0 111394 800 6 i_dout1_1[1]
port 108 nsew signal input
rlabel metal2 s 145838 0 145894 800 6 i_dout1_1[20]
port 109 nsew signal input
rlabel metal2 s 148690 0 148746 800 6 i_dout1_1[21]
port 110 nsew signal input
rlabel metal2 s 149610 0 149666 800 6 i_dout1_1[22]
port 111 nsew signal input
rlabel metal2 s 151542 0 151598 800 6 i_dout1_1[23]
port 112 nsew signal input
rlabel metal3 s 163720 145664 164520 145784 6 i_dout1_1[24]
port 113 nsew signal input
rlabel metal3 s 0 136960 800 137080 6 i_dout1_1[25]
port 114 nsew signal input
rlabel metal3 s 163720 151240 164520 151360 6 i_dout1_1[26]
port 115 nsew signal input
rlabel metal3 s 0 144712 800 144832 6 i_dout1_1[27]
port 116 nsew signal input
rlabel metal3 s 0 149880 800 150000 6 i_dout1_1[28]
port 117 nsew signal input
rlabel metal2 s 160190 0 160246 800 6 i_dout1_1[29]
port 118 nsew signal input
rlabel metal3 s 163720 20680 164520 20800 6 i_dout1_1[2]
port 119 nsew signal input
rlabel metal2 s 161018 165864 161074 166664 6 i_dout1_1[30]
port 120 nsew signal input
rlabel metal3 s 163720 165112 164520 165232 6 i_dout1_1[31]
port 121 nsew signal input
rlabel metal3 s 163720 26256 164520 26376 6 i_dout1_1[3]
port 122 nsew signal input
rlabel metal3 s 163720 40128 164520 40248 6 i_dout1_1[4]
port 123 nsew signal input
rlabel metal2 s 122838 0 122894 800 6 i_dout1_1[5]
port 124 nsew signal input
rlabel metal2 s 125690 0 125746 800 6 i_dout1_1[6]
port 125 nsew signal input
rlabel metal3 s 0 49920 800 50040 6 i_dout1_1[7]
port 126 nsew signal input
rlabel metal2 s 129646 165864 129702 166664 6 i_dout1_1[8]
port 127 nsew signal input
rlabel metal3 s 163720 84600 164520 84720 6 i_dout1_1[9]
port 128 nsew signal input
rlabel metal2 s 478 165864 534 166664 6 io_in[0]
port 129 nsew signal input
rlabel metal2 s 29826 165864 29882 166664 6 io_in[10]
port 130 nsew signal input
rlabel metal2 s 32770 165864 32826 166664 6 io_in[11]
port 131 nsew signal input
rlabel metal2 s 35714 165864 35770 166664 6 io_in[12]
port 132 nsew signal input
rlabel metal2 s 38658 165864 38714 166664 6 io_in[13]
port 133 nsew signal input
rlabel metal2 s 41602 165864 41658 166664 6 io_in[14]
port 134 nsew signal input
rlabel metal2 s 44454 165864 44510 166664 6 io_in[15]
port 135 nsew signal input
rlabel metal2 s 47398 165864 47454 166664 6 io_in[16]
port 136 nsew signal input
rlabel metal2 s 50342 165864 50398 166664 6 io_in[17]
port 137 nsew signal input
rlabel metal2 s 53286 165864 53342 166664 6 io_in[18]
port 138 nsew signal input
rlabel metal2 s 56230 165864 56286 166664 6 io_in[19]
port 139 nsew signal input
rlabel metal2 s 3330 165864 3386 166664 6 io_in[1]
port 140 nsew signal input
rlabel metal2 s 59174 165864 59230 166664 6 io_in[20]
port 141 nsew signal input
rlabel metal2 s 62118 165864 62174 166664 6 io_in[21]
port 142 nsew signal input
rlabel metal2 s 65062 165864 65118 166664 6 io_in[22]
port 143 nsew signal input
rlabel metal2 s 68006 165864 68062 166664 6 io_in[23]
port 144 nsew signal input
rlabel metal2 s 70950 165864 71006 166664 6 io_in[24]
port 145 nsew signal input
rlabel metal2 s 73894 165864 73950 166664 6 io_in[25]
port 146 nsew signal input
rlabel metal2 s 76838 165864 76894 166664 6 io_in[26]
port 147 nsew signal input
rlabel metal2 s 79782 165864 79838 166664 6 io_in[27]
port 148 nsew signal input
rlabel metal2 s 82726 165864 82782 166664 6 io_in[28]
port 149 nsew signal input
rlabel metal2 s 85578 165864 85634 166664 6 io_in[29]
port 150 nsew signal input
rlabel metal2 s 6274 165864 6330 166664 6 io_in[2]
port 151 nsew signal input
rlabel metal2 s 88522 165864 88578 166664 6 io_in[30]
port 152 nsew signal input
rlabel metal2 s 91466 165864 91522 166664 6 io_in[31]
port 153 nsew signal input
rlabel metal2 s 94410 165864 94466 166664 6 io_in[32]
port 154 nsew signal input
rlabel metal2 s 97354 165864 97410 166664 6 io_in[33]
port 155 nsew signal input
rlabel metal2 s 100298 165864 100354 166664 6 io_in[34]
port 156 nsew signal input
rlabel metal2 s 103242 165864 103298 166664 6 io_in[35]
port 157 nsew signal input
rlabel metal2 s 106186 165864 106242 166664 6 io_in[36]
port 158 nsew signal input
rlabel metal2 s 109130 165864 109186 166664 6 io_in[37]
port 159 nsew signal input
rlabel metal2 s 9218 165864 9274 166664 6 io_in[3]
port 160 nsew signal input
rlabel metal2 s 12162 165864 12218 166664 6 io_in[4]
port 161 nsew signal input
rlabel metal2 s 15106 165864 15162 166664 6 io_in[5]
port 162 nsew signal input
rlabel metal2 s 18050 165864 18106 166664 6 io_in[6]
port 163 nsew signal input
rlabel metal2 s 20994 165864 21050 166664 6 io_in[7]
port 164 nsew signal input
rlabel metal2 s 23938 165864 23994 166664 6 io_in[8]
port 165 nsew signal input
rlabel metal2 s 26882 165864 26938 166664 6 io_in[9]
port 166 nsew signal input
rlabel metal2 s 1398 165864 1454 166664 6 io_oeb[0]
port 167 nsew signal output
rlabel metal2 s 30746 165864 30802 166664 6 io_oeb[10]
port 168 nsew signal output
rlabel metal2 s 33690 165864 33746 166664 6 io_oeb[11]
port 169 nsew signal output
rlabel metal2 s 36634 165864 36690 166664 6 io_oeb[12]
port 170 nsew signal output
rlabel metal2 s 39578 165864 39634 166664 6 io_oeb[13]
port 171 nsew signal output
rlabel metal2 s 42522 165864 42578 166664 6 io_oeb[14]
port 172 nsew signal output
rlabel metal2 s 45466 165864 45522 166664 6 io_oeb[15]
port 173 nsew signal output
rlabel metal2 s 48410 165864 48466 166664 6 io_oeb[16]
port 174 nsew signal output
rlabel metal2 s 51354 165864 51410 166664 6 io_oeb[17]
port 175 nsew signal output
rlabel metal2 s 54298 165864 54354 166664 6 io_oeb[18]
port 176 nsew signal output
rlabel metal2 s 57242 165864 57298 166664 6 io_oeb[19]
port 177 nsew signal output
rlabel metal2 s 4342 165864 4398 166664 6 io_oeb[1]
port 178 nsew signal output
rlabel metal2 s 60186 165864 60242 166664 6 io_oeb[20]
port 179 nsew signal output
rlabel metal2 s 63130 165864 63186 166664 6 io_oeb[21]
port 180 nsew signal output
rlabel metal2 s 66074 165864 66130 166664 6 io_oeb[22]
port 181 nsew signal output
rlabel metal2 s 69018 165864 69074 166664 6 io_oeb[23]
port 182 nsew signal output
rlabel metal2 s 71870 165864 71926 166664 6 io_oeb[24]
port 183 nsew signal output
rlabel metal2 s 74814 165864 74870 166664 6 io_oeb[25]
port 184 nsew signal output
rlabel metal2 s 77758 165864 77814 166664 6 io_oeb[26]
port 185 nsew signal output
rlabel metal2 s 80702 165864 80758 166664 6 io_oeb[27]
port 186 nsew signal output
rlabel metal2 s 83646 165864 83702 166664 6 io_oeb[28]
port 187 nsew signal output
rlabel metal2 s 86590 165864 86646 166664 6 io_oeb[29]
port 188 nsew signal output
rlabel metal2 s 7286 165864 7342 166664 6 io_oeb[2]
port 189 nsew signal output
rlabel metal2 s 89534 165864 89590 166664 6 io_oeb[30]
port 190 nsew signal output
rlabel metal2 s 92478 165864 92534 166664 6 io_oeb[31]
port 191 nsew signal output
rlabel metal2 s 95422 165864 95478 166664 6 io_oeb[32]
port 192 nsew signal output
rlabel metal2 s 98366 165864 98422 166664 6 io_oeb[33]
port 193 nsew signal output
rlabel metal2 s 101310 165864 101366 166664 6 io_oeb[34]
port 194 nsew signal output
rlabel metal2 s 104254 165864 104310 166664 6 io_oeb[35]
port 195 nsew signal output
rlabel metal2 s 107198 165864 107254 166664 6 io_oeb[36]
port 196 nsew signal output
rlabel metal2 s 110142 165864 110198 166664 6 io_oeb[37]
port 197 nsew signal output
rlabel metal2 s 10230 165864 10286 166664 6 io_oeb[3]
port 198 nsew signal output
rlabel metal2 s 13174 165864 13230 166664 6 io_oeb[4]
port 199 nsew signal output
rlabel metal2 s 16118 165864 16174 166664 6 io_oeb[5]
port 200 nsew signal output
rlabel metal2 s 19062 165864 19118 166664 6 io_oeb[6]
port 201 nsew signal output
rlabel metal2 s 22006 165864 22062 166664 6 io_oeb[7]
port 202 nsew signal output
rlabel metal2 s 24950 165864 25006 166664 6 io_oeb[8]
port 203 nsew signal output
rlabel metal2 s 27894 165864 27950 166664 6 io_oeb[9]
port 204 nsew signal output
rlabel metal2 s 2410 165864 2466 166664 6 io_out[0]
port 205 nsew signal output
rlabel metal2 s 31758 165864 31814 166664 6 io_out[10]
port 206 nsew signal output
rlabel metal2 s 34702 165864 34758 166664 6 io_out[11]
port 207 nsew signal output
rlabel metal2 s 37646 165864 37702 166664 6 io_out[12]
port 208 nsew signal output
rlabel metal2 s 40590 165864 40646 166664 6 io_out[13]
port 209 nsew signal output
rlabel metal2 s 43534 165864 43590 166664 6 io_out[14]
port 210 nsew signal output
rlabel metal2 s 46478 165864 46534 166664 6 io_out[15]
port 211 nsew signal output
rlabel metal2 s 49422 165864 49478 166664 6 io_out[16]
port 212 nsew signal output
rlabel metal2 s 52366 165864 52422 166664 6 io_out[17]
port 213 nsew signal output
rlabel metal2 s 55310 165864 55366 166664 6 io_out[18]
port 214 nsew signal output
rlabel metal2 s 58162 165864 58218 166664 6 io_out[19]
port 215 nsew signal output
rlabel metal2 s 5354 165864 5410 166664 6 io_out[1]
port 216 nsew signal output
rlabel metal2 s 61106 165864 61162 166664 6 io_out[20]
port 217 nsew signal output
rlabel metal2 s 64050 165864 64106 166664 6 io_out[21]
port 218 nsew signal output
rlabel metal2 s 66994 165864 67050 166664 6 io_out[22]
port 219 nsew signal output
rlabel metal2 s 69938 165864 69994 166664 6 io_out[23]
port 220 nsew signal output
rlabel metal2 s 72882 165864 72938 166664 6 io_out[24]
port 221 nsew signal output
rlabel metal2 s 75826 165864 75882 166664 6 io_out[25]
port 222 nsew signal output
rlabel metal2 s 78770 165864 78826 166664 6 io_out[26]
port 223 nsew signal output
rlabel metal2 s 81714 165864 81770 166664 6 io_out[27]
port 224 nsew signal output
rlabel metal2 s 84658 165864 84714 166664 6 io_out[28]
port 225 nsew signal output
rlabel metal2 s 87602 165864 87658 166664 6 io_out[29]
port 226 nsew signal output
rlabel metal2 s 8298 165864 8354 166664 6 io_out[2]
port 227 nsew signal output
rlabel metal2 s 90546 165864 90602 166664 6 io_out[30]
port 228 nsew signal output
rlabel metal2 s 93490 165864 93546 166664 6 io_out[31]
port 229 nsew signal output
rlabel metal2 s 96434 165864 96490 166664 6 io_out[32]
port 230 nsew signal output
rlabel metal2 s 99286 165864 99342 166664 6 io_out[33]
port 231 nsew signal output
rlabel metal2 s 102230 165864 102286 166664 6 io_out[34]
port 232 nsew signal output
rlabel metal2 s 105174 165864 105230 166664 6 io_out[35]
port 233 nsew signal output
rlabel metal2 s 108118 165864 108174 166664 6 io_out[36]
port 234 nsew signal output
rlabel metal2 s 111062 165864 111118 166664 6 io_out[37]
port 235 nsew signal output
rlabel metal2 s 11242 165864 11298 166664 6 io_out[3]
port 236 nsew signal output
rlabel metal2 s 14186 165864 14242 166664 6 io_out[4]
port 237 nsew signal output
rlabel metal2 s 17038 165864 17094 166664 6 io_out[5]
port 238 nsew signal output
rlabel metal2 s 19982 165864 20038 166664 6 io_out[6]
port 239 nsew signal output
rlabel metal2 s 22926 165864 22982 166664 6 io_out[7]
port 240 nsew signal output
rlabel metal2 s 25870 165864 25926 166664 6 io_out[8]
port 241 nsew signal output
rlabel metal2 s 28814 165864 28870 166664 6 io_out[9]
port 242 nsew signal output
rlabel metal2 s 101770 0 101826 800 6 irq[0]
port 243 nsew signal output
rlabel metal2 s 102782 0 102838 800 6 irq[1]
port 244 nsew signal output
rlabel metal2 s 103702 0 103758 800 6 irq[2]
port 245 nsew signal output
rlabel metal2 s 114006 165864 114062 166664 6 o_addr1[0]
port 246 nsew signal output
rlabel metal3 s 0 14016 800 14136 6 o_addr1[1]
port 247 nsew signal output
rlabel metal3 s 0 26800 800 26920 6 o_addr1[2]
port 248 nsew signal output
rlabel metal2 s 120906 165864 120962 166664 6 o_addr1[3]
port 249 nsew signal output
rlabel metal2 s 120906 0 120962 800 6 o_addr1[4]
port 250 nsew signal output
rlabel metal3 s 163720 56856 164520 56976 6 o_addr1[5]
port 251 nsew signal output
rlabel metal2 s 127714 165864 127770 166664 6 o_addr1[6]
port 252 nsew signal output
rlabel metal2 s 128726 165864 128782 166664 6 o_addr1[7]
port 253 nsew signal output
rlabel metal3 s 0 57536 800 57656 6 o_addr1[8]
port 254 nsew signal output
rlabel metal2 s 112994 165864 113050 166664 6 o_addr1_1[0]
port 255 nsew signal output
rlabel metal3 s 163720 12384 164520 12504 6 o_addr1_1[1]
port 256 nsew signal output
rlabel metal2 s 114282 0 114338 800 6 o_addr1_1[2]
port 257 nsew signal output
rlabel metal3 s 163720 29112 164520 29232 6 o_addr1_1[3]
port 258 nsew signal output
rlabel metal3 s 163720 48560 164520 48680 6 o_addr1_1[4]
port 259 nsew signal output
rlabel metal2 s 124770 0 124826 800 6 o_addr1_1[5]
port 260 nsew signal output
rlabel metal3 s 0 42168 800 42288 6 o_addr1_1[6]
port 261 nsew signal output
rlabel metal2 s 129554 0 129610 800 6 o_addr1_1[7]
port 262 nsew signal output
rlabel metal3 s 163720 79024 164520 79144 6 o_addr1_1[8]
port 263 nsew signal output
rlabel metal2 s 112074 165864 112130 166664 6 o_csb0
port 264 nsew signal output
rlabel metal2 s 104714 0 104770 800 6 o_csb0_1
port 265 nsew signal output
rlabel metal3 s 0 1232 800 1352 6 o_csb1
port 266 nsew signal output
rlabel metal2 s 105634 0 105690 800 6 o_csb1_1
port 267 nsew signal output
rlabel metal2 s 115018 165864 115074 166664 6 o_din0[0]
port 268 nsew signal output
rlabel metal2 s 135258 0 135314 800 6 o_din0[10]
port 269 nsew signal output
rlabel metal3 s 0 83240 800 83360 6 o_din0[11]
port 270 nsew signal output
rlabel metal3 s 0 85688 800 85808 6 o_din0[12]
port 271 nsew signal output
rlabel metal3 s 0 90856 800 90976 6 o_din0[13]
port 272 nsew signal output
rlabel metal3 s 163720 101328 164520 101448 6 o_din0[14]
port 273 nsew signal output
rlabel metal2 s 140410 165864 140466 166664 6 o_din0[15]
port 274 nsew signal output
rlabel metal3 s 0 108808 800 108928 6 o_din0[16]
port 275 nsew signal output
rlabel metal2 s 142894 0 142950 800 6 o_din0[17]
port 276 nsew signal output
rlabel metal3 s 163720 115200 164520 115320 6 o_din0[18]
port 277 nsew signal output
rlabel metal3 s 163720 126216 164520 126336 6 o_din0[19]
port 278 nsew signal output
rlabel metal2 s 116950 165864 117006 166664 6 o_din0[1]
port 279 nsew signal output
rlabel metal3 s 0 119008 800 119128 6 o_din0[20]
port 280 nsew signal output
rlabel metal3 s 163720 131792 164520 131912 6 o_din0[21]
port 281 nsew signal output
rlabel metal3 s 163720 134648 164520 134768 6 o_din0[22]
port 282 nsew signal output
rlabel metal3 s 0 129344 800 129464 6 o_din0[23]
port 283 nsew signal output
rlabel metal2 s 154118 165864 154174 166664 6 o_din0[24]
port 284 nsew signal output
rlabel metal2 s 153474 0 153530 800 6 o_din0[25]
port 285 nsew signal output
rlabel metal2 s 157062 165864 157118 166664 6 o_din0[26]
port 286 nsew signal output
rlabel metal2 s 158258 0 158314 800 6 o_din0[27]
port 287 nsew signal output
rlabel metal3 s 0 157496 800 157616 6 o_din0[28]
port 288 nsew signal output
rlabel metal2 s 160006 165864 160062 166664 6 o_din0[29]
port 289 nsew signal output
rlabel metal3 s 163720 23536 164520 23656 6 o_din0[2]
port 290 nsew signal output
rlabel metal2 s 162030 165864 162086 166664 6 o_din0[30]
port 291 nsew signal output
rlabel metal2 s 163962 165864 164018 166664 6 o_din0[31]
port 292 nsew signal output
rlabel metal2 s 119066 0 119122 800 6 o_din0[3]
port 293 nsew signal output
rlabel metal2 s 122838 165864 122894 166664 6 o_din0[4]
port 294 nsew signal output
rlabel metal3 s 163720 59576 164520 59696 6 o_din0[5]
port 295 nsew signal output
rlabel metal3 s 0 44752 800 44872 6 o_din0[6]
port 296 nsew signal output
rlabel metal3 s 163720 70728 164520 70848 6 o_din0[7]
port 297 nsew signal output
rlabel metal3 s 0 60120 800 60240 6 o_din0[8]
port 298 nsew signal output
rlabel metal3 s 0 65288 800 65408 6 o_din0[9]
port 299 nsew signal output
rlabel metal3 s 163720 4088 164520 4208 6 o_din0_1[0]
port 300 nsew signal output
rlabel metal2 s 132590 165864 132646 166664 6 o_din0_1[10]
port 301 nsew signal output
rlabel metal2 s 136270 0 136326 800 6 o_din0_1[11]
port 302 nsew signal output
rlabel metal2 s 139122 0 139178 800 6 o_din0_1[12]
port 303 nsew signal output
rlabel metal3 s 0 88272 800 88392 6 o_din0_1[13]
port 304 nsew signal output
rlabel metal3 s 163720 98472 164520 98592 6 o_din0_1[14]
port 305 nsew signal output
rlabel metal3 s 163720 106768 164520 106888 6 o_din0_1[15]
port 306 nsew signal output
rlabel metal3 s 163720 112344 164520 112464 6 o_din0_1[16]
port 307 nsew signal output
rlabel metal2 s 142434 165864 142490 166664 6 o_din0_1[17]
port 308 nsew signal output
rlabel metal2 s 144366 165864 144422 166664 6 o_din0_1[18]
port 309 nsew signal output
rlabel metal3 s 163720 123496 164520 123616 6 o_din0_1[19]
port 310 nsew signal output
rlabel metal3 s 163720 15240 164520 15360 6 o_din0_1[1]
port 311 nsew signal output
rlabel metal2 s 147678 0 147734 800 6 o_din0_1[20]
port 312 nsew signal output
rlabel metal3 s 0 124176 800 124296 6 o_din0_1[21]
port 313 nsew signal output
rlabel metal2 s 150254 165864 150310 166664 6 o_din0_1[22]
port 314 nsew signal output
rlabel metal3 s 163720 142944 164520 143064 6 o_din0_1[23]
port 315 nsew signal output
rlabel metal2 s 152462 0 152518 800 6 o_din0_1[24]
port 316 nsew signal output
rlabel metal3 s 0 139544 800 139664 6 o_din0_1[25]
port 317 nsew signal output
rlabel metal3 s 0 142128 800 142248 6 o_din0_1[26]
port 318 nsew signal output
rlabel metal2 s 158074 165864 158130 166664 6 o_din0_1[27]
port 319 nsew signal output
rlabel metal3 s 0 154912 800 155032 6 o_din0_1[28]
port 320 nsew signal output
rlabel metal2 s 162030 0 162086 800 6 o_din0_1[29]
port 321 nsew signal output
rlabel metal2 s 115202 0 115258 800 6 o_din0_1[2]
port 322 nsew signal output
rlabel metal3 s 0 162664 800 162784 6 o_din0_1[30]
port 323 nsew signal output
rlabel metal2 s 163962 0 164018 800 6 o_din0_1[31]
port 324 nsew signal output
rlabel metal3 s 0 31968 800 32088 6 o_din0_1[3]
port 325 nsew signal output
rlabel metal2 s 121826 165864 121882 166664 6 o_din0_1[4]
port 326 nsew signal output
rlabel metal3 s 0 37000 800 37120 6 o_din0_1[5]
port 327 nsew signal output
rlabel metal3 s 163720 65152 164520 65272 6 o_din0_1[6]
port 328 nsew signal output
rlabel metal2 s 130474 0 130530 800 6 o_din0_1[7]
port 329 nsew signal output
rlabel metal2 s 132406 0 132462 800 6 o_din0_1[8]
port 330 nsew signal output
rlabel metal2 s 134338 0 134394 800 6 o_din0_1[9]
port 331 nsew signal output
rlabel metal3 s 0 6264 800 6384 6 o_waddr0[0]
port 332 nsew signal output
rlabel metal3 s 0 19048 800 19168 6 o_waddr0[1]
port 333 nsew signal output
rlabel metal3 s 0 29384 800 29504 6 o_waddr0[2]
port 334 nsew signal output
rlabel metal3 s 163720 31832 164520 31952 6 o_waddr0[3]
port 335 nsew signal output
rlabel metal3 s 163720 51280 164520 51400 6 o_waddr0[4]
port 336 nsew signal output
rlabel metal2 s 125782 165864 125838 166664 6 o_waddr0[5]
port 337 nsew signal output
rlabel metal3 s 0 47336 800 47456 6 o_waddr0[6]
port 338 nsew signal output
rlabel metal3 s 0 54952 800 55072 6 o_waddr0[7]
port 339 nsew signal output
rlabel metal3 s 0 62704 800 62824 6 o_waddr0[8]
port 340 nsew signal output
rlabel metal2 s 110418 0 110474 800 6 o_waddr0_1[0]
port 341 nsew signal output
rlabel metal3 s 0 16600 800 16720 6 o_waddr0_1[1]
port 342 nsew signal output
rlabel metal2 s 117962 165864 118018 166664 6 o_waddr0_1[2]
port 343 nsew signal output
rlabel metal2 s 119986 0 120042 800 6 o_waddr0_1[3]
port 344 nsew signal output
rlabel metal2 s 121918 0 121974 800 6 o_waddr0_1[4]
port 345 nsew signal output
rlabel metal2 s 124770 165864 124826 166664 6 o_waddr0_1[5]
port 346 nsew signal output
rlabel metal3 s 163720 68008 164520 68128 6 o_waddr0_1[6]
port 347 nsew signal output
rlabel metal3 s 0 52368 800 52488 6 o_waddr0_1[7]
port 348 nsew signal output
rlabel metal2 s 130658 165864 130714 166664 6 o_waddr0_1[8]
port 349 nsew signal output
rlabel metal3 s 0 3680 800 3800 6 o_web0
port 350 nsew signal output
rlabel metal2 s 106554 0 106610 800 6 o_web0_1
port 351 nsew signal output
rlabel metal3 s 0 8848 800 8968 6 o_wmask0[0]
port 352 nsew signal output
rlabel metal3 s 0 21632 800 21752 6 o_wmask0[1]
port 353 nsew signal output
rlabel metal2 s 119894 165864 119950 166664 6 o_wmask0[2]
port 354 nsew signal output
rlabel metal3 s 163720 34688 164520 34808 6 o_wmask0[3]
port 355 nsew signal output
rlabel metal3 s 163720 6808 164520 6928 6 o_wmask0_1[0]
port 356 nsew signal output
rlabel metal2 s 112350 0 112406 800 6 o_wmask0_1[1]
port 357 nsew signal output
rlabel metal2 s 118882 165864 118938 166664 6 o_wmask0_1[2]
port 358 nsew signal output
rlabel metal3 s 0 34552 800 34672 6 o_wmask0_1[3]
port 359 nsew signal output
rlabel metal4 s 4208 2128 4528 164336 6 vccd1
port 360 nsew power input
rlabel metal4 s 34928 2128 35248 164336 6 vccd1
port 360 nsew power input
rlabel metal4 s 65648 2128 65968 164336 6 vccd1
port 360 nsew power input
rlabel metal4 s 96368 2128 96688 164336 6 vccd1
port 360 nsew power input
rlabel metal4 s 127088 2128 127408 164336 6 vccd1
port 360 nsew power input
rlabel metal4 s 157808 2128 158128 164336 6 vccd1
port 360 nsew power input
rlabel metal4 s 19568 2128 19888 164336 6 vssd1
port 361 nsew ground input
rlabel metal4 s 50288 2128 50608 164336 6 vssd1
port 361 nsew ground input
rlabel metal4 s 81008 2128 81328 164336 6 vssd1
port 361 nsew ground input
rlabel metal4 s 111728 2128 112048 164336 6 vssd1
port 361 nsew ground input
rlabel metal4 s 142448 2128 142768 164336 6 vssd1
port 361 nsew ground input
rlabel metal2 s 478 0 534 800 6 wb_clk_i
port 362 nsew signal input
rlabel metal2 s 1398 0 1454 800 6 wb_rst_i
port 363 nsew signal input
rlabel metal2 s 2318 0 2374 800 6 wbs_ack_o
port 364 nsew signal output
rlabel metal2 s 6182 0 6238 800 6 wbs_adr_i[0]
port 365 nsew signal input
rlabel metal2 s 38658 0 38714 800 6 wbs_adr_i[10]
port 366 nsew signal input
rlabel metal2 s 41602 0 41658 800 6 wbs_adr_i[11]
port 367 nsew signal input
rlabel metal2 s 44454 0 44510 800 6 wbs_adr_i[12]
port 368 nsew signal input
rlabel metal2 s 47306 0 47362 800 6 wbs_adr_i[13]
port 369 nsew signal input
rlabel metal2 s 50158 0 50214 800 6 wbs_adr_i[14]
port 370 nsew signal input
rlabel metal2 s 53010 0 53066 800 6 wbs_adr_i[15]
port 371 nsew signal input
rlabel metal2 s 55862 0 55918 800 6 wbs_adr_i[16]
port 372 nsew signal input
rlabel metal2 s 58806 0 58862 800 6 wbs_adr_i[17]
port 373 nsew signal input
rlabel metal2 s 61658 0 61714 800 6 wbs_adr_i[18]
port 374 nsew signal input
rlabel metal2 s 64510 0 64566 800 6 wbs_adr_i[19]
port 375 nsew signal input
rlabel metal2 s 9954 0 10010 800 6 wbs_adr_i[1]
port 376 nsew signal input
rlabel metal2 s 67362 0 67418 800 6 wbs_adr_i[20]
port 377 nsew signal input
rlabel metal2 s 70214 0 70270 800 6 wbs_adr_i[21]
port 378 nsew signal input
rlabel metal2 s 73158 0 73214 800 6 wbs_adr_i[22]
port 379 nsew signal input
rlabel metal2 s 76010 0 76066 800 6 wbs_adr_i[23]
port 380 nsew signal input
rlabel metal2 s 78862 0 78918 800 6 wbs_adr_i[24]
port 381 nsew signal input
rlabel metal2 s 81714 0 81770 800 6 wbs_adr_i[25]
port 382 nsew signal input
rlabel metal2 s 84566 0 84622 800 6 wbs_adr_i[26]
port 383 nsew signal input
rlabel metal2 s 87418 0 87474 800 6 wbs_adr_i[27]
port 384 nsew signal input
rlabel metal2 s 90362 0 90418 800 6 wbs_adr_i[28]
port 385 nsew signal input
rlabel metal2 s 93214 0 93270 800 6 wbs_adr_i[29]
port 386 nsew signal input
rlabel metal2 s 13818 0 13874 800 6 wbs_adr_i[2]
port 387 nsew signal input
rlabel metal2 s 96066 0 96122 800 6 wbs_adr_i[30]
port 388 nsew signal input
rlabel metal2 s 98918 0 98974 800 6 wbs_adr_i[31]
port 389 nsew signal input
rlabel metal2 s 17682 0 17738 800 6 wbs_adr_i[3]
port 390 nsew signal input
rlabel metal2 s 21454 0 21510 800 6 wbs_adr_i[4]
port 391 nsew signal input
rlabel metal2 s 24306 0 24362 800 6 wbs_adr_i[5]
port 392 nsew signal input
rlabel metal2 s 27250 0 27306 800 6 wbs_adr_i[6]
port 393 nsew signal input
rlabel metal2 s 30102 0 30158 800 6 wbs_adr_i[7]
port 394 nsew signal input
rlabel metal2 s 32954 0 33010 800 6 wbs_adr_i[8]
port 395 nsew signal input
rlabel metal2 s 35806 0 35862 800 6 wbs_adr_i[9]
port 396 nsew signal input
rlabel metal2 s 3330 0 3386 800 6 wbs_cyc_i
port 397 nsew signal input
rlabel metal2 s 7102 0 7158 800 6 wbs_dat_i[0]
port 398 nsew signal input
rlabel metal2 s 39670 0 39726 800 6 wbs_dat_i[10]
port 399 nsew signal input
rlabel metal2 s 42522 0 42578 800 6 wbs_dat_i[11]
port 400 nsew signal input
rlabel metal2 s 45374 0 45430 800 6 wbs_dat_i[12]
port 401 nsew signal input
rlabel metal2 s 48226 0 48282 800 6 wbs_dat_i[13]
port 402 nsew signal input
rlabel metal2 s 51078 0 51134 800 6 wbs_dat_i[14]
port 403 nsew signal input
rlabel metal2 s 54022 0 54078 800 6 wbs_dat_i[15]
port 404 nsew signal input
rlabel metal2 s 56874 0 56930 800 6 wbs_dat_i[16]
port 405 nsew signal input
rlabel metal2 s 59726 0 59782 800 6 wbs_dat_i[17]
port 406 nsew signal input
rlabel metal2 s 62578 0 62634 800 6 wbs_dat_i[18]
port 407 nsew signal input
rlabel metal2 s 65430 0 65486 800 6 wbs_dat_i[19]
port 408 nsew signal input
rlabel metal2 s 10966 0 11022 800 6 wbs_dat_i[1]
port 409 nsew signal input
rlabel metal2 s 68374 0 68430 800 6 wbs_dat_i[20]
port 410 nsew signal input
rlabel metal2 s 71226 0 71282 800 6 wbs_dat_i[21]
port 411 nsew signal input
rlabel metal2 s 74078 0 74134 800 6 wbs_dat_i[22]
port 412 nsew signal input
rlabel metal2 s 76930 0 76986 800 6 wbs_dat_i[23]
port 413 nsew signal input
rlabel metal2 s 79782 0 79838 800 6 wbs_dat_i[24]
port 414 nsew signal input
rlabel metal2 s 82726 0 82782 800 6 wbs_dat_i[25]
port 415 nsew signal input
rlabel metal2 s 85578 0 85634 800 6 wbs_dat_i[26]
port 416 nsew signal input
rlabel metal2 s 88430 0 88486 800 6 wbs_dat_i[27]
port 417 nsew signal input
rlabel metal2 s 91282 0 91338 800 6 wbs_dat_i[28]
port 418 nsew signal input
rlabel metal2 s 94134 0 94190 800 6 wbs_dat_i[29]
port 419 nsew signal input
rlabel metal2 s 14738 0 14794 800 6 wbs_dat_i[2]
port 420 nsew signal input
rlabel metal2 s 96986 0 97042 800 6 wbs_dat_i[30]
port 421 nsew signal input
rlabel metal2 s 99930 0 99986 800 6 wbs_dat_i[31]
port 422 nsew signal input
rlabel metal2 s 18602 0 18658 800 6 wbs_dat_i[3]
port 423 nsew signal input
rlabel metal2 s 22466 0 22522 800 6 wbs_dat_i[4]
port 424 nsew signal input
rlabel metal2 s 25318 0 25374 800 6 wbs_dat_i[5]
port 425 nsew signal input
rlabel metal2 s 28170 0 28226 800 6 wbs_dat_i[6]
port 426 nsew signal input
rlabel metal2 s 31022 0 31078 800 6 wbs_dat_i[7]
port 427 nsew signal input
rlabel metal2 s 33874 0 33930 800 6 wbs_dat_i[8]
port 428 nsew signal input
rlabel metal2 s 36818 0 36874 800 6 wbs_dat_i[9]
port 429 nsew signal input
rlabel metal2 s 8114 0 8170 800 6 wbs_dat_o[0]
port 430 nsew signal output
rlabel metal2 s 40590 0 40646 800 6 wbs_dat_o[10]
port 431 nsew signal output
rlabel metal2 s 43442 0 43498 800 6 wbs_dat_o[11]
port 432 nsew signal output
rlabel metal2 s 46294 0 46350 800 6 wbs_dat_o[12]
port 433 nsew signal output
rlabel metal2 s 49238 0 49294 800 6 wbs_dat_o[13]
port 434 nsew signal output
rlabel metal2 s 52090 0 52146 800 6 wbs_dat_o[14]
port 435 nsew signal output
rlabel metal2 s 54942 0 54998 800 6 wbs_dat_o[15]
port 436 nsew signal output
rlabel metal2 s 57794 0 57850 800 6 wbs_dat_o[16]
port 437 nsew signal output
rlabel metal2 s 60646 0 60702 800 6 wbs_dat_o[17]
port 438 nsew signal output
rlabel metal2 s 63590 0 63646 800 6 wbs_dat_o[18]
port 439 nsew signal output
rlabel metal2 s 66442 0 66498 800 6 wbs_dat_o[19]
port 440 nsew signal output
rlabel metal2 s 11886 0 11942 800 6 wbs_dat_o[1]
port 441 nsew signal output
rlabel metal2 s 69294 0 69350 800 6 wbs_dat_o[20]
port 442 nsew signal output
rlabel metal2 s 72146 0 72202 800 6 wbs_dat_o[21]
port 443 nsew signal output
rlabel metal2 s 74998 0 75054 800 6 wbs_dat_o[22]
port 444 nsew signal output
rlabel metal2 s 77942 0 77998 800 6 wbs_dat_o[23]
port 445 nsew signal output
rlabel metal2 s 80794 0 80850 800 6 wbs_dat_o[24]
port 446 nsew signal output
rlabel metal2 s 83646 0 83702 800 6 wbs_dat_o[25]
port 447 nsew signal output
rlabel metal2 s 86498 0 86554 800 6 wbs_dat_o[26]
port 448 nsew signal output
rlabel metal2 s 89350 0 89406 800 6 wbs_dat_o[27]
port 449 nsew signal output
rlabel metal2 s 92202 0 92258 800 6 wbs_dat_o[28]
port 450 nsew signal output
rlabel metal2 s 95146 0 95202 800 6 wbs_dat_o[29]
port 451 nsew signal output
rlabel metal2 s 15750 0 15806 800 6 wbs_dat_o[2]
port 452 nsew signal output
rlabel metal2 s 97998 0 98054 800 6 wbs_dat_o[30]
port 453 nsew signal output
rlabel metal2 s 100850 0 100906 800 6 wbs_dat_o[31]
port 454 nsew signal output
rlabel metal2 s 19522 0 19578 800 6 wbs_dat_o[3]
port 455 nsew signal output
rlabel metal2 s 23386 0 23442 800 6 wbs_dat_o[4]
port 456 nsew signal output
rlabel metal2 s 26238 0 26294 800 6 wbs_dat_o[5]
port 457 nsew signal output
rlabel metal2 s 29090 0 29146 800 6 wbs_dat_o[6]
port 458 nsew signal output
rlabel metal2 s 32034 0 32090 800 6 wbs_dat_o[7]
port 459 nsew signal output
rlabel metal2 s 34886 0 34942 800 6 wbs_dat_o[8]
port 460 nsew signal output
rlabel metal2 s 37738 0 37794 800 6 wbs_dat_o[9]
port 461 nsew signal output
rlabel metal2 s 9034 0 9090 800 6 wbs_sel_i[0]
port 462 nsew signal input
rlabel metal2 s 12898 0 12954 800 6 wbs_sel_i[1]
port 463 nsew signal input
rlabel metal2 s 16670 0 16726 800 6 wbs_sel_i[2]
port 464 nsew signal input
rlabel metal2 s 20534 0 20590 800 6 wbs_sel_i[3]
port 465 nsew signal input
rlabel metal2 s 4250 0 4306 800 6 wbs_stb_i
port 466 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 wbs_we_i
port 467 nsew signal input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 164520 166664
string LEFview TRUE
string GDS_FILE /project/openlane/user_proj/runs/user_proj/results/magic/user_proj.gds
string GDS_END 79876404
string GDS_START 1378264
<< end >>

