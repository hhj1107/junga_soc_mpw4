magic
tech sky130A
magscale 1 2
timestamp 1640471712
<< obsli1 >>
rect 1104 2159 163731 164305
<< obsm1 >>
rect 474 8 164114 164336
<< metal2 >>
rect 478 165957 534 166757
rect 1398 165957 1454 166757
rect 2318 165957 2374 166757
rect 3330 165957 3386 166757
rect 4250 165957 4306 166757
rect 5262 165957 5318 166757
rect 6182 165957 6238 166757
rect 7102 165957 7158 166757
rect 8114 165957 8170 166757
rect 9034 165957 9090 166757
rect 10046 165957 10102 166757
rect 10966 165957 11022 166757
rect 11886 165957 11942 166757
rect 12898 165957 12954 166757
rect 13818 165957 13874 166757
rect 14830 165957 14886 166757
rect 15750 165957 15806 166757
rect 16670 165957 16726 166757
rect 17682 165957 17738 166757
rect 18602 165957 18658 166757
rect 19614 165957 19670 166757
rect 20534 165957 20590 166757
rect 21454 165957 21510 166757
rect 22466 165957 22522 166757
rect 23386 165957 23442 166757
rect 24398 165957 24454 166757
rect 25318 165957 25374 166757
rect 26238 165957 26294 166757
rect 27250 165957 27306 166757
rect 28170 165957 28226 166757
rect 29182 165957 29238 166757
rect 30102 165957 30158 166757
rect 31022 165957 31078 166757
rect 32034 165957 32090 166757
rect 32954 165957 33010 166757
rect 33966 165957 34022 166757
rect 34886 165957 34942 166757
rect 35806 165957 35862 166757
rect 36818 165957 36874 166757
rect 37738 165957 37794 166757
rect 38750 165957 38806 166757
rect 39670 165957 39726 166757
rect 40590 165957 40646 166757
rect 41602 165957 41658 166757
rect 42522 165957 42578 166757
rect 43534 165957 43590 166757
rect 44454 165957 44510 166757
rect 45374 165957 45430 166757
rect 46386 165957 46442 166757
rect 47306 165957 47362 166757
rect 48318 165957 48374 166757
rect 49238 165957 49294 166757
rect 50158 165957 50214 166757
rect 51170 165957 51226 166757
rect 52090 165957 52146 166757
rect 53102 165957 53158 166757
rect 54022 165957 54078 166757
rect 54942 165957 54998 166757
rect 55954 165957 56010 166757
rect 56874 165957 56930 166757
rect 57886 165957 57942 166757
rect 58806 165957 58862 166757
rect 59726 165957 59782 166757
rect 60738 165957 60794 166757
rect 61658 165957 61714 166757
rect 62670 165957 62726 166757
rect 63590 165957 63646 166757
rect 64510 165957 64566 166757
rect 65522 165957 65578 166757
rect 66442 165957 66498 166757
rect 67454 165957 67510 166757
rect 68374 165957 68430 166757
rect 69294 165957 69350 166757
rect 70306 165957 70362 166757
rect 71226 165957 71282 166757
rect 72238 165957 72294 166757
rect 73158 165957 73214 166757
rect 74078 165957 74134 166757
rect 75090 165957 75146 166757
rect 76010 165957 76066 166757
rect 77022 165957 77078 166757
rect 77942 165957 77998 166757
rect 78862 165957 78918 166757
rect 79874 165957 79930 166757
rect 80794 165957 80850 166757
rect 81806 165957 81862 166757
rect 82726 165957 82782 166757
rect 83646 165957 83702 166757
rect 84658 165957 84714 166757
rect 85578 165957 85634 166757
rect 86590 165957 86646 166757
rect 87510 165957 87566 166757
rect 88430 165957 88486 166757
rect 89442 165957 89498 166757
rect 90362 165957 90418 166757
rect 91374 165957 91430 166757
rect 92294 165957 92350 166757
rect 93214 165957 93270 166757
rect 94226 165957 94282 166757
rect 95146 165957 95202 166757
rect 96158 165957 96214 166757
rect 97078 165957 97134 166757
rect 97998 165957 98054 166757
rect 99010 165957 99066 166757
rect 99930 165957 99986 166757
rect 100942 165957 100998 166757
rect 101862 165957 101918 166757
rect 102782 165957 102838 166757
rect 103794 165957 103850 166757
rect 104714 165957 104770 166757
rect 105726 165957 105782 166757
rect 106646 165957 106702 166757
rect 107566 165957 107622 166757
rect 108578 165957 108634 166757
rect 109498 165957 109554 166757
rect 110510 165957 110566 166757
rect 111430 165957 111486 166757
rect 112350 165957 112406 166757
rect 113362 165957 113418 166757
rect 114282 165957 114338 166757
rect 115294 165957 115350 166757
rect 116214 165957 116270 166757
rect 117134 165957 117190 166757
rect 118146 165957 118202 166757
rect 119066 165957 119122 166757
rect 120078 165957 120134 166757
rect 120998 165957 121054 166757
rect 121918 165957 121974 166757
rect 122930 165957 122986 166757
rect 123850 165957 123906 166757
rect 124862 165957 124918 166757
rect 125782 165957 125838 166757
rect 126702 165957 126758 166757
rect 127714 165957 127770 166757
rect 128634 165957 128690 166757
rect 129646 165957 129702 166757
rect 130566 165957 130622 166757
rect 131486 165957 131542 166757
rect 132498 165957 132554 166757
rect 133418 165957 133474 166757
rect 134430 165957 134486 166757
rect 135350 165957 135406 166757
rect 136270 165957 136326 166757
rect 137282 165957 137338 166757
rect 138202 165957 138258 166757
rect 139214 165957 139270 166757
rect 140134 165957 140190 166757
rect 141054 165957 141110 166757
rect 142066 165957 142122 166757
rect 142986 165957 143042 166757
rect 143998 165957 144054 166757
rect 144918 165957 144974 166757
rect 145838 165957 145894 166757
rect 146850 165957 146906 166757
rect 147770 165957 147826 166757
rect 148782 165957 148838 166757
rect 149702 165957 149758 166757
rect 150622 165957 150678 166757
rect 151634 165957 151690 166757
rect 152554 165957 152610 166757
rect 153566 165957 153622 166757
rect 154486 165957 154542 166757
rect 155406 165957 155462 166757
rect 156418 165957 156474 166757
rect 157338 165957 157394 166757
rect 158350 165957 158406 166757
rect 159270 165957 159326 166757
rect 160190 165957 160246 166757
rect 161202 165957 161258 166757
rect 162122 165957 162178 166757
rect 163134 165957 163190 166757
rect 164054 165957 164110 166757
rect 478 0 534 800
rect 1398 0 1454 800
rect 2410 0 2466 800
rect 3422 0 3478 800
rect 4434 0 4490 800
rect 5446 0 5502 800
rect 6458 0 6514 800
rect 7470 0 7526 800
rect 8482 0 8538 800
rect 9494 0 9550 800
rect 10506 0 10562 800
rect 11518 0 11574 800
rect 12530 0 12586 800
rect 13542 0 13598 800
rect 14554 0 14610 800
rect 15566 0 15622 800
rect 16578 0 16634 800
rect 17590 0 17646 800
rect 18602 0 18658 800
rect 19614 0 19670 800
rect 20626 0 20682 800
rect 21638 0 21694 800
rect 22650 0 22706 800
rect 23662 0 23718 800
rect 24674 0 24730 800
rect 25686 0 25742 800
rect 26698 0 26754 800
rect 27710 0 27766 800
rect 28722 0 28778 800
rect 29734 0 29790 800
rect 30746 0 30802 800
rect 31758 0 31814 800
rect 32770 0 32826 800
rect 33782 0 33838 800
rect 34794 0 34850 800
rect 35806 0 35862 800
rect 36818 0 36874 800
rect 37830 0 37886 800
rect 38842 0 38898 800
rect 39854 0 39910 800
rect 40866 0 40922 800
rect 41786 0 41842 800
rect 42798 0 42854 800
rect 43810 0 43866 800
rect 44822 0 44878 800
rect 45834 0 45890 800
rect 46846 0 46902 800
rect 47858 0 47914 800
rect 48870 0 48926 800
rect 49882 0 49938 800
rect 50894 0 50950 800
rect 51906 0 51962 800
rect 52918 0 52974 800
rect 53930 0 53986 800
rect 54942 0 54998 800
rect 55954 0 56010 800
rect 56966 0 57022 800
rect 57978 0 58034 800
rect 58990 0 59046 800
rect 60002 0 60058 800
rect 61014 0 61070 800
rect 62026 0 62082 800
rect 63038 0 63094 800
rect 64050 0 64106 800
rect 65062 0 65118 800
rect 66074 0 66130 800
rect 67086 0 67142 800
rect 68098 0 68154 800
rect 69110 0 69166 800
rect 70122 0 70178 800
rect 71134 0 71190 800
rect 72146 0 72202 800
rect 73158 0 73214 800
rect 74170 0 74226 800
rect 75182 0 75238 800
rect 76194 0 76250 800
rect 77206 0 77262 800
rect 78218 0 78274 800
rect 79230 0 79286 800
rect 80242 0 80298 800
rect 81254 0 81310 800
rect 82266 0 82322 800
rect 83186 0 83242 800
rect 84198 0 84254 800
rect 85210 0 85266 800
rect 86222 0 86278 800
rect 87234 0 87290 800
rect 88246 0 88302 800
rect 89258 0 89314 800
rect 90270 0 90326 800
rect 91282 0 91338 800
rect 92294 0 92350 800
rect 93306 0 93362 800
rect 94318 0 94374 800
rect 95330 0 95386 800
rect 96342 0 96398 800
rect 97354 0 97410 800
rect 98366 0 98422 800
rect 99378 0 99434 800
rect 100390 0 100446 800
rect 101402 0 101458 800
rect 102414 0 102470 800
rect 103426 0 103482 800
rect 104438 0 104494 800
rect 105450 0 105506 800
rect 106462 0 106518 800
rect 107474 0 107530 800
rect 108486 0 108542 800
rect 109498 0 109554 800
rect 110510 0 110566 800
rect 111522 0 111578 800
rect 112534 0 112590 800
rect 113546 0 113602 800
rect 114558 0 114614 800
rect 115570 0 115626 800
rect 116582 0 116638 800
rect 117594 0 117650 800
rect 118606 0 118662 800
rect 119618 0 119674 800
rect 120630 0 120686 800
rect 121642 0 121698 800
rect 122654 0 122710 800
rect 123666 0 123722 800
rect 124586 0 124642 800
rect 125598 0 125654 800
rect 126610 0 126666 800
rect 127622 0 127678 800
rect 128634 0 128690 800
rect 129646 0 129702 800
rect 130658 0 130714 800
rect 131670 0 131726 800
rect 132682 0 132738 800
rect 133694 0 133750 800
rect 134706 0 134762 800
rect 135718 0 135774 800
rect 136730 0 136786 800
rect 137742 0 137798 800
rect 138754 0 138810 800
rect 139766 0 139822 800
rect 140778 0 140834 800
rect 141790 0 141846 800
rect 142802 0 142858 800
rect 143814 0 143870 800
rect 144826 0 144882 800
rect 145838 0 145894 800
rect 146850 0 146906 800
rect 147862 0 147918 800
rect 148874 0 148930 800
rect 149886 0 149942 800
rect 150898 0 150954 800
rect 151910 0 151966 800
rect 152922 0 152978 800
rect 153934 0 153990 800
rect 154946 0 155002 800
rect 155958 0 156014 800
rect 156970 0 157026 800
rect 157982 0 158038 800
rect 158994 0 159050 800
rect 160006 0 160062 800
rect 161018 0 161074 800
rect 162030 0 162086 800
rect 163042 0 163098 800
rect 164054 0 164110 800
<< obsm2 >>
rect 18 165901 422 166002
rect 590 165901 1342 166002
rect 1510 165901 2262 166002
rect 2430 165901 3274 166002
rect 3442 165901 4194 166002
rect 4362 165901 5206 166002
rect 5374 165901 6126 166002
rect 6294 165901 7046 166002
rect 7214 165901 8058 166002
rect 8226 165901 8978 166002
rect 9146 165901 9990 166002
rect 10158 165901 10910 166002
rect 11078 165901 11830 166002
rect 11998 165901 12842 166002
rect 13010 165901 13762 166002
rect 13930 165901 14774 166002
rect 14942 165901 15694 166002
rect 15862 165901 16614 166002
rect 16782 165901 17626 166002
rect 17794 165901 18546 166002
rect 18714 165901 19558 166002
rect 19726 165901 20478 166002
rect 20646 165901 21398 166002
rect 21566 165901 22410 166002
rect 22578 165901 23330 166002
rect 23498 165901 24342 166002
rect 24510 165901 25262 166002
rect 25430 165901 26182 166002
rect 26350 165901 27194 166002
rect 27362 165901 28114 166002
rect 28282 165901 29126 166002
rect 29294 165901 30046 166002
rect 30214 165901 30966 166002
rect 31134 165901 31978 166002
rect 32146 165901 32898 166002
rect 33066 165901 33910 166002
rect 34078 165901 34830 166002
rect 34998 165901 35750 166002
rect 35918 165901 36762 166002
rect 36930 165901 37682 166002
rect 37850 165901 38694 166002
rect 38862 165901 39614 166002
rect 39782 165901 40534 166002
rect 40702 165901 41546 166002
rect 41714 165901 42466 166002
rect 42634 165901 43478 166002
rect 43646 165901 44398 166002
rect 44566 165901 45318 166002
rect 45486 165901 46330 166002
rect 46498 165901 47250 166002
rect 47418 165901 48262 166002
rect 48430 165901 49182 166002
rect 49350 165901 50102 166002
rect 50270 165901 51114 166002
rect 51282 165901 52034 166002
rect 52202 165901 53046 166002
rect 53214 165901 53966 166002
rect 54134 165901 54886 166002
rect 55054 165901 55898 166002
rect 56066 165901 56818 166002
rect 56986 165901 57830 166002
rect 57998 165901 58750 166002
rect 58918 165901 59670 166002
rect 59838 165901 60682 166002
rect 60850 165901 61602 166002
rect 61770 165901 62614 166002
rect 62782 165901 63534 166002
rect 63702 165901 64454 166002
rect 64622 165901 65466 166002
rect 65634 165901 66386 166002
rect 66554 165901 67398 166002
rect 67566 165901 68318 166002
rect 68486 165901 69238 166002
rect 69406 165901 70250 166002
rect 70418 165901 71170 166002
rect 71338 165901 72182 166002
rect 72350 165901 73102 166002
rect 73270 165901 74022 166002
rect 74190 165901 75034 166002
rect 75202 165901 75954 166002
rect 76122 165901 76966 166002
rect 77134 165901 77886 166002
rect 78054 165901 78806 166002
rect 78974 165901 79818 166002
rect 79986 165901 80738 166002
rect 80906 165901 81750 166002
rect 81918 165901 82670 166002
rect 82838 165901 83590 166002
rect 83758 165901 84602 166002
rect 84770 165901 85522 166002
rect 85690 165901 86534 166002
rect 86702 165901 87454 166002
rect 87622 165901 88374 166002
rect 88542 165901 89386 166002
rect 89554 165901 90306 166002
rect 90474 165901 91318 166002
rect 91486 165901 92238 166002
rect 92406 165901 93158 166002
rect 93326 165901 94170 166002
rect 94338 165901 95090 166002
rect 95258 165901 96102 166002
rect 96270 165901 97022 166002
rect 97190 165901 97942 166002
rect 98110 165901 98954 166002
rect 99122 165901 99874 166002
rect 100042 165901 100886 166002
rect 101054 165901 101806 166002
rect 101974 165901 102726 166002
rect 102894 165901 103738 166002
rect 103906 165901 104658 166002
rect 104826 165901 105670 166002
rect 105838 165901 106590 166002
rect 106758 165901 107510 166002
rect 107678 165901 108522 166002
rect 108690 165901 109442 166002
rect 109610 165901 110454 166002
rect 110622 165901 111374 166002
rect 111542 165901 112294 166002
rect 112462 165901 113306 166002
rect 113474 165901 114226 166002
rect 114394 165901 115238 166002
rect 115406 165901 116158 166002
rect 116326 165901 117078 166002
rect 117246 165901 118090 166002
rect 118258 165901 119010 166002
rect 119178 165901 120022 166002
rect 120190 165901 120942 166002
rect 121110 165901 121862 166002
rect 122030 165901 122874 166002
rect 123042 165901 123794 166002
rect 123962 165901 124806 166002
rect 124974 165901 125726 166002
rect 125894 165901 126646 166002
rect 126814 165901 127658 166002
rect 127826 165901 128578 166002
rect 128746 165901 129590 166002
rect 129758 165901 130510 166002
rect 130678 165901 131430 166002
rect 131598 165901 132442 166002
rect 132610 165901 133362 166002
rect 133530 165901 134374 166002
rect 134542 165901 135294 166002
rect 135462 165901 136214 166002
rect 136382 165901 137226 166002
rect 137394 165901 138146 166002
rect 138314 165901 139158 166002
rect 139326 165901 140078 166002
rect 140246 165901 140998 166002
rect 141166 165901 142010 166002
rect 142178 165901 142930 166002
rect 143098 165901 143942 166002
rect 144110 165901 144862 166002
rect 145030 165901 145782 166002
rect 145950 165901 146794 166002
rect 146962 165901 147714 166002
rect 147882 165901 148726 166002
rect 148894 165901 149646 166002
rect 149814 165901 150566 166002
rect 150734 165901 151578 166002
rect 151746 165901 152498 166002
rect 152666 165901 153510 166002
rect 153678 165901 154430 166002
rect 154598 165901 155350 166002
rect 155518 165901 156362 166002
rect 156530 165901 157282 166002
rect 157450 165901 158294 166002
rect 158462 165901 159214 166002
rect 159382 165901 160134 166002
rect 160302 165901 161146 166002
rect 161314 165901 162066 166002
rect 162234 165901 163078 166002
rect 163246 165901 163998 166002
rect 18 856 164108 165901
rect 18 2 422 856
rect 590 2 1342 856
rect 1510 2 2354 856
rect 2522 2 3366 856
rect 3534 2 4378 856
rect 4546 2 5390 856
rect 5558 2 6402 856
rect 6570 2 7414 856
rect 7582 2 8426 856
rect 8594 2 9438 856
rect 9606 2 10450 856
rect 10618 2 11462 856
rect 11630 2 12474 856
rect 12642 2 13486 856
rect 13654 2 14498 856
rect 14666 2 15510 856
rect 15678 2 16522 856
rect 16690 2 17534 856
rect 17702 2 18546 856
rect 18714 2 19558 856
rect 19726 2 20570 856
rect 20738 2 21582 856
rect 21750 2 22594 856
rect 22762 2 23606 856
rect 23774 2 24618 856
rect 24786 2 25630 856
rect 25798 2 26642 856
rect 26810 2 27654 856
rect 27822 2 28666 856
rect 28834 2 29678 856
rect 29846 2 30690 856
rect 30858 2 31702 856
rect 31870 2 32714 856
rect 32882 2 33726 856
rect 33894 2 34738 856
rect 34906 2 35750 856
rect 35918 2 36762 856
rect 36930 2 37774 856
rect 37942 2 38786 856
rect 38954 2 39798 856
rect 39966 2 40810 856
rect 40978 2 41730 856
rect 41898 2 42742 856
rect 42910 2 43754 856
rect 43922 2 44766 856
rect 44934 2 45778 856
rect 45946 2 46790 856
rect 46958 2 47802 856
rect 47970 2 48814 856
rect 48982 2 49826 856
rect 49994 2 50838 856
rect 51006 2 51850 856
rect 52018 2 52862 856
rect 53030 2 53874 856
rect 54042 2 54886 856
rect 55054 2 55898 856
rect 56066 2 56910 856
rect 57078 2 57922 856
rect 58090 2 58934 856
rect 59102 2 59946 856
rect 60114 2 60958 856
rect 61126 2 61970 856
rect 62138 2 62982 856
rect 63150 2 63994 856
rect 64162 2 65006 856
rect 65174 2 66018 856
rect 66186 2 67030 856
rect 67198 2 68042 856
rect 68210 2 69054 856
rect 69222 2 70066 856
rect 70234 2 71078 856
rect 71246 2 72090 856
rect 72258 2 73102 856
rect 73270 2 74114 856
rect 74282 2 75126 856
rect 75294 2 76138 856
rect 76306 2 77150 856
rect 77318 2 78162 856
rect 78330 2 79174 856
rect 79342 2 80186 856
rect 80354 2 81198 856
rect 81366 2 82210 856
rect 82378 2 83130 856
rect 83298 2 84142 856
rect 84310 2 85154 856
rect 85322 2 86166 856
rect 86334 2 87178 856
rect 87346 2 88190 856
rect 88358 2 89202 856
rect 89370 2 90214 856
rect 90382 2 91226 856
rect 91394 2 92238 856
rect 92406 2 93250 856
rect 93418 2 94262 856
rect 94430 2 95274 856
rect 95442 2 96286 856
rect 96454 2 97298 856
rect 97466 2 98310 856
rect 98478 2 99322 856
rect 99490 2 100334 856
rect 100502 2 101346 856
rect 101514 2 102358 856
rect 102526 2 103370 856
rect 103538 2 104382 856
rect 104550 2 105394 856
rect 105562 2 106406 856
rect 106574 2 107418 856
rect 107586 2 108430 856
rect 108598 2 109442 856
rect 109610 2 110454 856
rect 110622 2 111466 856
rect 111634 2 112478 856
rect 112646 2 113490 856
rect 113658 2 114502 856
rect 114670 2 115514 856
rect 115682 2 116526 856
rect 116694 2 117538 856
rect 117706 2 118550 856
rect 118718 2 119562 856
rect 119730 2 120574 856
rect 120742 2 121586 856
rect 121754 2 122598 856
rect 122766 2 123610 856
rect 123778 2 124530 856
rect 124698 2 125542 856
rect 125710 2 126554 856
rect 126722 2 127566 856
rect 127734 2 128578 856
rect 128746 2 129590 856
rect 129758 2 130602 856
rect 130770 2 131614 856
rect 131782 2 132626 856
rect 132794 2 133638 856
rect 133806 2 134650 856
rect 134818 2 135662 856
rect 135830 2 136674 856
rect 136842 2 137686 856
rect 137854 2 138698 856
rect 138866 2 139710 856
rect 139878 2 140722 856
rect 140890 2 141734 856
rect 141902 2 142746 856
rect 142914 2 143758 856
rect 143926 2 144770 856
rect 144938 2 145782 856
rect 145950 2 146794 856
rect 146962 2 147806 856
rect 147974 2 148818 856
rect 148986 2 149830 856
rect 149998 2 150842 856
rect 151010 2 151854 856
rect 152022 2 152866 856
rect 153034 2 153878 856
rect 154046 2 154890 856
rect 155058 2 155902 856
rect 156070 2 156914 856
rect 157082 2 157926 856
rect 158094 2 158938 856
rect 159106 2 159950 856
rect 160118 2 160962 856
rect 161130 2 161974 856
rect 162142 2 162986 856
rect 163154 2 163998 856
<< metal3 >>
rect 0 165384 800 165504
rect 163813 165112 164613 165232
rect 0 163072 800 163192
rect 163813 162256 164613 162376
rect 0 160760 800 160880
rect 163813 159400 164613 159520
rect 0 158448 800 158568
rect 163813 156544 164613 156664
rect 0 156136 800 156256
rect 0 153824 800 153944
rect 163813 153688 164613 153808
rect 0 151512 800 151632
rect 163813 150832 164613 150952
rect 0 149200 800 149320
rect 163813 147976 164613 148096
rect 0 146888 800 147008
rect 163813 144984 164613 145104
rect 0 144576 800 144696
rect 0 142264 800 142384
rect 163813 142128 164613 142248
rect 0 139952 800 140072
rect 163813 139272 164613 139392
rect 0 137640 800 137760
rect 163813 136416 164613 136536
rect 0 135328 800 135448
rect 163813 133560 164613 133680
rect 0 133016 800 133136
rect 0 130704 800 130824
rect 163813 130704 164613 130824
rect 0 128392 800 128512
rect 163813 127848 164613 127968
rect 0 126080 800 126200
rect 163813 124856 164613 124976
rect 0 123768 800 123888
rect 163813 122000 164613 122120
rect 0 121456 800 121576
rect 0 119144 800 119264
rect 163813 119144 164613 119264
rect 0 116832 800 116952
rect 163813 116288 164613 116408
rect 0 114520 800 114640
rect 163813 113432 164613 113552
rect 0 112208 800 112328
rect 163813 110576 164613 110696
rect 0 109896 800 110016
rect 0 107584 800 107704
rect 163813 107720 164613 107840
rect 0 105272 800 105392
rect 163813 104728 164613 104848
rect 0 102960 800 103080
rect 163813 101872 164613 101992
rect 0 100648 800 100768
rect 163813 99016 164613 99136
rect 0 98336 800 98456
rect 0 96024 800 96144
rect 163813 96160 164613 96280
rect 0 93712 800 93832
rect 163813 93304 164613 93424
rect 0 91400 800 91520
rect 163813 90448 164613 90568
rect 0 89088 800 89208
rect 163813 87592 164613 87712
rect 0 86776 800 86896
rect 163813 84736 164613 84856
rect 0 84464 800 84584
rect 0 82016 800 82136
rect 163813 81744 164613 81864
rect 0 79704 800 79824
rect 163813 78888 164613 79008
rect 0 77392 800 77512
rect 163813 76032 164613 76152
rect 0 75080 800 75200
rect 163813 73176 164613 73296
rect 0 72768 800 72888
rect 0 70456 800 70576
rect 163813 70320 164613 70440
rect 0 68144 800 68264
rect 163813 67464 164613 67584
rect 0 65832 800 65952
rect 163813 64608 164613 64728
rect 0 63520 800 63640
rect 163813 61616 164613 61736
rect 0 61208 800 61328
rect 0 58896 800 59016
rect 163813 58760 164613 58880
rect 0 56584 800 56704
rect 163813 55904 164613 56024
rect 0 54272 800 54392
rect 163813 53048 164613 53168
rect 0 51960 800 52080
rect 163813 50192 164613 50312
rect 0 49648 800 49768
rect 0 47336 800 47456
rect 163813 47336 164613 47456
rect 0 45024 800 45144
rect 163813 44480 164613 44600
rect 0 42712 800 42832
rect 163813 41488 164613 41608
rect 0 40400 800 40520
rect 163813 38632 164613 38752
rect 0 38088 800 38208
rect 0 35776 800 35896
rect 163813 35776 164613 35896
rect 0 33464 800 33584
rect 163813 32920 164613 33040
rect 0 31152 800 31272
rect 163813 30064 164613 30184
rect 0 28840 800 28960
rect 163813 27208 164613 27328
rect 0 26528 800 26648
rect 0 24216 800 24336
rect 163813 24352 164613 24472
rect 0 21904 800 22024
rect 163813 21360 164613 21480
rect 0 19592 800 19712
rect 163813 18504 164613 18624
rect 0 17280 800 17400
rect 163813 15648 164613 15768
rect 0 14968 800 15088
rect 0 12656 800 12776
rect 163813 12792 164613 12912
rect 0 10344 800 10464
rect 163813 9936 164613 10056
rect 0 8032 800 8152
rect 163813 7080 164613 7200
rect 0 5720 800 5840
rect 163813 4224 164613 4344
rect 0 3408 800 3528
rect 163813 1368 164613 1488
rect 0 1096 800 1216
<< obsm3 >>
rect 13 165032 163733 165205
rect 13 163272 163813 165032
rect 880 162992 163813 163272
rect 13 162456 163813 162992
rect 13 162176 163733 162456
rect 13 160960 163813 162176
rect 880 160680 163813 160960
rect 13 159600 163813 160680
rect 13 159320 163733 159600
rect 13 158648 163813 159320
rect 880 158368 163813 158648
rect 13 156744 163813 158368
rect 13 156464 163733 156744
rect 13 156336 163813 156464
rect 880 156056 163813 156336
rect 13 154024 163813 156056
rect 880 153888 163813 154024
rect 880 153744 163733 153888
rect 13 153608 163733 153744
rect 13 151712 163813 153608
rect 880 151432 163813 151712
rect 13 151032 163813 151432
rect 13 150752 163733 151032
rect 13 149400 163813 150752
rect 880 149120 163813 149400
rect 13 148176 163813 149120
rect 13 147896 163733 148176
rect 13 147088 163813 147896
rect 880 146808 163813 147088
rect 13 145184 163813 146808
rect 13 144904 163733 145184
rect 13 144776 163813 144904
rect 880 144496 163813 144776
rect 13 142464 163813 144496
rect 880 142328 163813 142464
rect 880 142184 163733 142328
rect 13 142048 163733 142184
rect 13 140152 163813 142048
rect 880 139872 163813 140152
rect 13 139472 163813 139872
rect 13 139192 163733 139472
rect 13 137840 163813 139192
rect 880 137560 163813 137840
rect 13 136616 163813 137560
rect 13 136336 163733 136616
rect 13 135528 163813 136336
rect 880 135248 163813 135528
rect 13 133760 163813 135248
rect 13 133480 163733 133760
rect 13 133216 163813 133480
rect 880 132936 163813 133216
rect 13 130904 163813 132936
rect 880 130624 163733 130904
rect 13 128592 163813 130624
rect 880 128312 163813 128592
rect 13 128048 163813 128312
rect 13 127768 163733 128048
rect 13 126280 163813 127768
rect 880 126000 163813 126280
rect 13 125056 163813 126000
rect 13 124776 163733 125056
rect 13 123968 163813 124776
rect 880 123688 163813 123968
rect 13 122200 163813 123688
rect 13 121920 163733 122200
rect 13 121656 163813 121920
rect 880 121376 163813 121656
rect 13 119344 163813 121376
rect 880 119064 163733 119344
rect 13 117032 163813 119064
rect 880 116752 163813 117032
rect 13 116488 163813 116752
rect 13 116208 163733 116488
rect 13 114720 163813 116208
rect 880 114440 163813 114720
rect 13 113632 163813 114440
rect 13 113352 163733 113632
rect 13 112408 163813 113352
rect 880 112128 163813 112408
rect 13 110776 163813 112128
rect 13 110496 163733 110776
rect 13 110096 163813 110496
rect 880 109816 163813 110096
rect 13 107920 163813 109816
rect 13 107784 163733 107920
rect 880 107640 163733 107784
rect 880 107504 163813 107640
rect 13 105472 163813 107504
rect 880 105192 163813 105472
rect 13 104928 163813 105192
rect 13 104648 163733 104928
rect 13 103160 163813 104648
rect 880 102880 163813 103160
rect 13 102072 163813 102880
rect 13 101792 163733 102072
rect 13 100848 163813 101792
rect 880 100568 163813 100848
rect 13 99216 163813 100568
rect 13 98936 163733 99216
rect 13 98536 163813 98936
rect 880 98256 163813 98536
rect 13 96360 163813 98256
rect 13 96224 163733 96360
rect 880 96080 163733 96224
rect 880 95944 163813 96080
rect 13 93912 163813 95944
rect 880 93632 163813 93912
rect 13 93504 163813 93632
rect 13 93224 163733 93504
rect 13 91600 163813 93224
rect 880 91320 163813 91600
rect 13 90648 163813 91320
rect 13 90368 163733 90648
rect 13 89288 163813 90368
rect 880 89008 163813 89288
rect 13 87792 163813 89008
rect 13 87512 163733 87792
rect 13 86976 163813 87512
rect 880 86696 163813 86976
rect 13 84936 163813 86696
rect 13 84664 163733 84936
rect 880 84656 163733 84664
rect 880 84384 163813 84656
rect 13 82216 163813 84384
rect 880 81944 163813 82216
rect 880 81936 163733 81944
rect 13 81664 163733 81936
rect 13 79904 163813 81664
rect 880 79624 163813 79904
rect 13 79088 163813 79624
rect 13 78808 163733 79088
rect 13 77592 163813 78808
rect 880 77312 163813 77592
rect 13 76232 163813 77312
rect 13 75952 163733 76232
rect 13 75280 163813 75952
rect 880 75000 163813 75280
rect 13 73376 163813 75000
rect 13 73096 163733 73376
rect 13 72968 163813 73096
rect 880 72688 163813 72968
rect 13 70656 163813 72688
rect 880 70520 163813 70656
rect 880 70376 163733 70520
rect 13 70240 163733 70376
rect 13 68344 163813 70240
rect 880 68064 163813 68344
rect 13 67664 163813 68064
rect 13 67384 163733 67664
rect 13 66032 163813 67384
rect 880 65752 163813 66032
rect 13 64808 163813 65752
rect 13 64528 163733 64808
rect 13 63720 163813 64528
rect 880 63440 163813 63720
rect 13 61816 163813 63440
rect 13 61536 163733 61816
rect 13 61408 163813 61536
rect 880 61128 163813 61408
rect 13 59096 163813 61128
rect 880 58960 163813 59096
rect 880 58816 163733 58960
rect 13 58680 163733 58816
rect 13 56784 163813 58680
rect 880 56504 163813 56784
rect 13 56104 163813 56504
rect 13 55824 163733 56104
rect 13 54472 163813 55824
rect 880 54192 163813 54472
rect 13 53248 163813 54192
rect 13 52968 163733 53248
rect 13 52160 163813 52968
rect 880 51880 163813 52160
rect 13 50392 163813 51880
rect 13 50112 163733 50392
rect 13 49848 163813 50112
rect 880 49568 163813 49848
rect 13 47536 163813 49568
rect 880 47256 163733 47536
rect 13 45224 163813 47256
rect 880 44944 163813 45224
rect 13 44680 163813 44944
rect 13 44400 163733 44680
rect 13 42912 163813 44400
rect 880 42632 163813 42912
rect 13 41688 163813 42632
rect 13 41408 163733 41688
rect 13 40600 163813 41408
rect 880 40320 163813 40600
rect 13 38832 163813 40320
rect 13 38552 163733 38832
rect 13 38288 163813 38552
rect 880 38008 163813 38288
rect 13 35976 163813 38008
rect 880 35696 163733 35976
rect 13 33664 163813 35696
rect 880 33384 163813 33664
rect 13 33120 163813 33384
rect 13 32840 163733 33120
rect 13 31352 163813 32840
rect 880 31072 163813 31352
rect 13 30264 163813 31072
rect 13 29984 163733 30264
rect 13 29040 163813 29984
rect 880 28760 163813 29040
rect 13 27408 163813 28760
rect 13 27128 163733 27408
rect 13 26728 163813 27128
rect 880 26448 163813 26728
rect 13 24552 163813 26448
rect 13 24416 163733 24552
rect 880 24272 163733 24416
rect 880 24136 163813 24272
rect 13 22104 163813 24136
rect 880 21824 163813 22104
rect 13 21560 163813 21824
rect 13 21280 163733 21560
rect 13 19792 163813 21280
rect 880 19512 163813 19792
rect 13 18704 163813 19512
rect 13 18424 163733 18704
rect 13 17480 163813 18424
rect 880 17200 163813 17480
rect 13 15848 163813 17200
rect 13 15568 163733 15848
rect 13 15168 163813 15568
rect 880 14888 163813 15168
rect 13 12992 163813 14888
rect 13 12856 163733 12992
rect 880 12712 163733 12856
rect 880 12576 163813 12712
rect 13 10544 163813 12576
rect 880 10264 163813 10544
rect 13 10136 163813 10264
rect 13 9856 163733 10136
rect 13 8232 163813 9856
rect 880 7952 163813 8232
rect 13 7280 163813 7952
rect 13 7000 163733 7280
rect 13 5920 163813 7000
rect 880 5640 163813 5920
rect 13 4424 163813 5640
rect 13 4144 163733 4424
rect 13 3608 163813 4144
rect 880 3328 163813 3608
rect 13 1568 163813 3328
rect 13 1296 163733 1568
rect 880 1288 163733 1296
rect 880 1016 163813 1288
rect 13 35 163813 1016
<< metal4 >>
rect 4208 2128 4528 164336
rect 19568 2128 19888 164336
rect 34928 2128 35248 164336
rect 50288 2128 50608 164336
rect 65648 2128 65968 164336
rect 81008 2128 81328 164336
rect 96368 2128 96688 164336
rect 111728 2128 112048 164336
rect 127088 2128 127408 164336
rect 142448 2128 142768 164336
rect 157808 2128 158128 164336
<< obsm4 >>
rect 243 2048 4128 163981
rect 4608 2048 19488 163981
rect 19968 2048 34848 163981
rect 35328 2048 50208 163981
rect 50688 2048 65568 163981
rect 66048 2048 80928 163981
rect 81408 2048 96288 163981
rect 96768 2048 111648 163981
rect 112128 2048 127008 163981
rect 127488 2048 142368 163981
rect 142848 2048 146405 163981
rect 243 1939 146405 2048
<< labels >>
rlabel metal3 s 163813 4224 164613 4344 6 i_dout0[0]
port 1 nsew signal input
rlabel metal2 s 134430 165957 134486 166757 6 i_dout0[10]
port 2 nsew signal input
rlabel metal2 s 137742 0 137798 800 6 i_dout0[11]
port 3 nsew signal input
rlabel metal2 s 137282 165957 137338 166757 6 i_dout0[12]
port 4 nsew signal input
rlabel metal2 s 141790 0 141846 800 6 i_dout0[13]
port 5 nsew signal input
rlabel metal3 s 163813 93304 164613 93424 6 i_dout0[14]
port 6 nsew signal input
rlabel metal2 s 144826 0 144882 800 6 i_dout0[15]
port 7 nsew signal input
rlabel metal3 s 0 96024 800 96144 6 i_dout0[16]
port 8 nsew signal input
rlabel metal3 s 163813 101872 164613 101992 6 i_dout0[17]
port 9 nsew signal input
rlabel metal3 s 163813 110576 164613 110696 6 i_dout0[18]
port 10 nsew signal input
rlabel metal3 s 163813 119144 164613 119264 6 i_dout0[19]
port 11 nsew signal input
rlabel metal3 s 163813 9936 164613 10056 6 i_dout0[1]
port 12 nsew signal input
rlabel metal3 s 163813 124856 164613 124976 6 i_dout0[20]
port 13 nsew signal input
rlabel metal3 s 163813 130704 164613 130824 6 i_dout0[21]
port 14 nsew signal input
rlabel metal3 s 0 119144 800 119264 6 i_dout0[22]
port 15 nsew signal input
rlabel metal2 s 152922 0 152978 800 6 i_dout0[23]
port 16 nsew signal input
rlabel metal3 s 163813 142128 164613 142248 6 i_dout0[24]
port 17 nsew signal input
rlabel metal3 s 163813 144984 164613 145104 6 i_dout0[25]
port 18 nsew signal input
rlabel metal3 s 163813 150832 164613 150952 6 i_dout0[26]
port 19 nsew signal input
rlabel metal3 s 0 142264 800 142384 6 i_dout0[27]
port 20 nsew signal input
rlabel metal2 s 160006 0 160062 800 6 i_dout0[28]
port 21 nsew signal input
rlabel metal2 s 161202 165957 161258 166757 6 i_dout0[29]
port 22 nsew signal input
rlabel metal2 s 116214 165957 116270 166757 6 i_dout0[2]
port 23 nsew signal input
rlabel metal3 s 0 160760 800 160880 6 i_dout0[30]
port 24 nsew signal input
rlabel metal2 s 163134 165957 163190 166757 6 i_dout0[31]
port 25 nsew signal input
rlabel metal3 s 163813 24352 164613 24472 6 i_dout0[3]
port 26 nsew signal input
rlabel metal3 s 163813 35776 164613 35896 6 i_dout0[4]
port 27 nsew signal input
rlabel metal2 s 121918 165957 121974 166757 6 i_dout0[5]
port 28 nsew signal input
rlabel metal2 s 131670 0 131726 800 6 i_dout0[6]
port 29 nsew signal input
rlabel metal3 s 0 56584 800 56704 6 i_dout0[7]
port 30 nsew signal input
rlabel metal2 s 128634 165957 128690 166757 6 i_dout0[8]
port 31 nsew signal input
rlabel metal3 s 163813 78888 164613 79008 6 i_dout0[9]
port 32 nsew signal input
rlabel metal2 s 110510 165957 110566 166757 6 i_dout0_1[0]
port 33 nsew signal input
rlabel metal2 s 132498 165957 132554 166757 6 i_dout0_1[10]
port 34 nsew signal input
rlabel metal3 s 0 75080 800 75200 6 i_dout0_1[11]
port 35 nsew signal input
rlabel metal3 s 0 82016 800 82136 6 i_dout0_1[12]
port 36 nsew signal input
rlabel metal2 s 140778 0 140834 800 6 i_dout0_1[13]
port 37 nsew signal input
rlabel metal2 s 142802 0 142858 800 6 i_dout0_1[14]
port 38 nsew signal input
rlabel metal2 s 142066 165957 142122 166757 6 i_dout0_1[15]
port 39 nsew signal input
rlabel metal2 s 143998 165957 144054 166757 6 i_dout0_1[16]
port 40 nsew signal input
rlabel metal3 s 163813 99016 164613 99136 6 i_dout0_1[17]
port 41 nsew signal input
rlabel metal3 s 0 102960 800 103080 6 i_dout0_1[18]
port 42 nsew signal input
rlabel metal3 s 0 105272 800 105392 6 i_dout0_1[19]
port 43 nsew signal input
rlabel metal3 s 0 12656 800 12776 6 i_dout0_1[1]
port 44 nsew signal input
rlabel metal3 s 0 109896 800 110016 6 i_dout0_1[20]
port 45 nsew signal input
rlabel metal2 s 151634 165957 151690 166757 6 i_dout0_1[21]
port 46 nsew signal input
rlabel metal2 s 150898 0 150954 800 6 i_dout0_1[22]
port 47 nsew signal input
rlabel metal2 s 152554 165957 152610 166757 6 i_dout0_1[23]
port 48 nsew signal input
rlabel metal3 s 163813 139272 164613 139392 6 i_dout0_1[24]
port 49 nsew signal input
rlabel metal3 s 0 133016 800 133136 6 i_dout0_1[25]
port 50 nsew signal input
rlabel metal3 s 0 135328 800 135448 6 i_dout0_1[26]
port 51 nsew signal input
rlabel metal3 s 0 139952 800 140072 6 i_dout0_1[27]
port 52 nsew signal input
rlabel metal2 s 157982 0 158038 800 6 i_dout0_1[28]
port 53 nsew signal input
rlabel metal2 s 160190 165957 160246 166757 6 i_dout0_1[29]
port 54 nsew signal input
rlabel metal3 s 163813 15648 164613 15768 6 i_dout0_1[2]
port 55 nsew signal input
rlabel metal3 s 0 156136 800 156256 6 i_dout0_1[30]
port 56 nsew signal input
rlabel metal3 s 0 163072 800 163192 6 i_dout0_1[31]
port 57 nsew signal input
rlabel metal3 s 0 24216 800 24336 6 i_dout0_1[3]
port 58 nsew signal input
rlabel metal3 s 0 33464 800 33584 6 i_dout0_1[4]
port 59 nsew signal input
rlabel metal2 s 120998 165957 121054 166757 6 i_dout0_1[5]
port 60 nsew signal input
rlabel metal2 s 123850 165957 123906 166757 6 i_dout0_1[6]
port 61 nsew signal input
rlabel metal3 s 0 54272 800 54392 6 i_dout0_1[7]
port 62 nsew signal input
rlabel metal2 s 127714 165957 127770 166757 6 i_dout0_1[8]
port 63 nsew signal input
rlabel metal3 s 163813 76032 164613 76152 6 i_dout0_1[9]
port 64 nsew signal input
rlabel metal2 s 111430 165957 111486 166757 6 i_dout1[0]
port 65 nsew signal input
rlabel metal2 s 135350 165957 135406 166757 6 i_dout1[10]
port 66 nsew signal input
rlabel metal2 s 136270 165957 136326 166757 6 i_dout1[11]
port 67 nsew signal input
rlabel metal2 s 138202 165957 138258 166757 6 i_dout1[12]
port 68 nsew signal input
rlabel metal3 s 163813 87592 164613 87712 6 i_dout1[13]
port 69 nsew signal input
rlabel metal2 s 143814 0 143870 800 6 i_dout1[14]
port 70 nsew signal input
rlabel metal3 s 0 91400 800 91520 6 i_dout1[15]
port 71 nsew signal input
rlabel metal3 s 0 98336 800 98456 6 i_dout1[16]
port 72 nsew signal input
rlabel metal2 s 146850 0 146906 800 6 i_dout1[17]
port 73 nsew signal input
rlabel metal3 s 163813 113432 164613 113552 6 i_dout1[18]
port 74 nsew signal input
rlabel metal2 s 148782 165957 148838 166757 6 i_dout1[19]
port 75 nsew signal input
rlabel metal3 s 0 14968 800 15088 6 i_dout1[1]
port 76 nsew signal input
rlabel metal3 s 0 112208 800 112328 6 i_dout1[20]
port 77 nsew signal input
rlabel metal2 s 148874 0 148930 800 6 i_dout1[21]
port 78 nsew signal input
rlabel metal2 s 151910 0 151966 800 6 i_dout1[22]
port 79 nsew signal input
rlabel metal3 s 0 126080 800 126200 6 i_dout1[23]
port 80 nsew signal input
rlabel metal2 s 154946 0 155002 800 6 i_dout1[24]
port 81 nsew signal input
rlabel metal2 s 155406 165957 155462 166757 6 i_dout1[25]
port 82 nsew signal input
rlabel metal2 s 156970 0 157026 800 6 i_dout1[26]
port 83 nsew signal input
rlabel metal3 s 163813 159400 164613 159520 6 i_dout1[27]
port 84 nsew signal input
rlabel metal3 s 0 144576 800 144696 6 i_dout1[28]
port 85 nsew signal input
rlabel metal3 s 163813 162256 164613 162376 6 i_dout1[29]
port 86 nsew signal input
rlabel metal2 s 122654 0 122710 800 6 i_dout1[2]
port 87 nsew signal input
rlabel metal2 s 161018 0 161074 800 6 i_dout1[30]
port 88 nsew signal input
rlabel metal3 s 0 165384 800 165504 6 i_dout1[31]
port 89 nsew signal input
rlabel metal3 s 0 26528 800 26648 6 i_dout1[3]
port 90 nsew signal input
rlabel metal2 s 129646 0 129702 800 6 i_dout1[4]
port 91 nsew signal input
rlabel metal3 s 0 40400 800 40520 6 i_dout1[5]
port 92 nsew signal input
rlabel metal3 s 163813 55904 164613 56024 6 i_dout1[6]
port 93 nsew signal input
rlabel metal3 s 163813 61616 164613 61736 6 i_dout1[7]
port 94 nsew signal input
rlabel metal2 s 129646 165957 129702 166757 6 i_dout1[8]
port 95 nsew signal input
rlabel metal3 s 163813 81744 164613 81864 6 i_dout1[9]
port 96 nsew signal input
rlabel metal3 s 0 5720 800 5840 6 i_dout1_1[0]
port 97 nsew signal input
rlabel metal2 s 133418 165957 133474 166757 6 i_dout1_1[10]
port 98 nsew signal input
rlabel metal3 s 0 77392 800 77512 6 i_dout1_1[11]
port 99 nsew signal input
rlabel metal3 s 0 84464 800 84584 6 i_dout1_1[12]
port 100 nsew signal input
rlabel metal3 s 0 86776 800 86896 6 i_dout1_1[13]
port 101 nsew signal input
rlabel metal3 s 163813 90448 164613 90568 6 i_dout1_1[14]
port 102 nsew signal input
rlabel metal2 s 142986 165957 143042 166757 6 i_dout1_1[15]
port 103 nsew signal input
rlabel metal3 s 163813 96160 164613 96280 6 i_dout1_1[16]
port 104 nsew signal input
rlabel metal3 s 0 100648 800 100768 6 i_dout1_1[17]
port 105 nsew signal input
rlabel metal2 s 146850 165957 146906 166757 6 i_dout1_1[18]
port 106 nsew signal input
rlabel metal3 s 163813 116288 164613 116408 6 i_dout1_1[19]
port 107 nsew signal input
rlabel metal2 s 112350 165957 112406 166757 6 i_dout1_1[1]
port 108 nsew signal input
rlabel metal3 s 163813 122000 164613 122120 6 i_dout1_1[20]
port 109 nsew signal input
rlabel metal3 s 0 114520 800 114640 6 i_dout1_1[21]
port 110 nsew signal input
rlabel metal3 s 163813 133560 164613 133680 6 i_dout1_1[22]
port 111 nsew signal input
rlabel metal2 s 153566 165957 153622 166757 6 i_dout1_1[23]
port 112 nsew signal input
rlabel metal2 s 153934 0 153990 800 6 i_dout1_1[24]
port 113 nsew signal input
rlabel metal2 s 155958 0 156014 800 6 i_dout1_1[25]
port 114 nsew signal input
rlabel metal3 s 163813 147976 164613 148096 6 i_dout1_1[26]
port 115 nsew signal input
rlabel metal3 s 163813 156544 164613 156664 6 i_dout1_1[27]
port 116 nsew signal input
rlabel metal2 s 158994 0 159050 800 6 i_dout1_1[28]
port 117 nsew signal input
rlabel metal3 s 0 151512 800 151632 6 i_dout1_1[29]
port 118 nsew signal input
rlabel metal2 s 121642 0 121698 800 6 i_dout1_1[2]
port 119 nsew signal input
rlabel metal3 s 0 158448 800 158568 6 i_dout1_1[30]
port 120 nsew signal input
rlabel metal2 s 163042 0 163098 800 6 i_dout1_1[31]
port 121 nsew signal input
rlabel metal2 s 125598 0 125654 800 6 i_dout1_1[3]
port 122 nsew signal input
rlabel metal3 s 163813 32920 164613 33040 6 i_dout1_1[4]
port 123 nsew signal input
rlabel metal3 s 0 38088 800 38208 6 i_dout1_1[5]
port 124 nsew signal input
rlabel metal3 s 0 45024 800 45144 6 i_dout1_1[6]
port 125 nsew signal input
rlabel metal2 s 125782 165957 125838 166757 6 i_dout1_1[7]
port 126 nsew signal input
rlabel metal2 s 134706 0 134762 800 6 i_dout1_1[8]
port 127 nsew signal input
rlabel metal3 s 0 65832 800 65952 6 i_dout1_1[9]
port 128 nsew signal input
rlabel metal2 s 478 165957 534 166757 6 io_in[0]
port 129 nsew signal input
rlabel metal2 s 29182 165957 29238 166757 6 io_in[10]
port 130 nsew signal input
rlabel metal2 s 32034 165957 32090 166757 6 io_in[11]
port 131 nsew signal input
rlabel metal2 s 34886 165957 34942 166757 6 io_in[12]
port 132 nsew signal input
rlabel metal2 s 37738 165957 37794 166757 6 io_in[13]
port 133 nsew signal input
rlabel metal2 s 40590 165957 40646 166757 6 io_in[14]
port 134 nsew signal input
rlabel metal2 s 43534 165957 43590 166757 6 io_in[15]
port 135 nsew signal input
rlabel metal2 s 46386 165957 46442 166757 6 io_in[16]
port 136 nsew signal input
rlabel metal2 s 49238 165957 49294 166757 6 io_in[17]
port 137 nsew signal input
rlabel metal2 s 52090 165957 52146 166757 6 io_in[18]
port 138 nsew signal input
rlabel metal2 s 54942 165957 54998 166757 6 io_in[19]
port 139 nsew signal input
rlabel metal2 s 3330 165957 3386 166757 6 io_in[1]
port 140 nsew signal input
rlabel metal2 s 57886 165957 57942 166757 6 io_in[20]
port 141 nsew signal input
rlabel metal2 s 60738 165957 60794 166757 6 io_in[21]
port 142 nsew signal input
rlabel metal2 s 63590 165957 63646 166757 6 io_in[22]
port 143 nsew signal input
rlabel metal2 s 66442 165957 66498 166757 6 io_in[23]
port 144 nsew signal input
rlabel metal2 s 69294 165957 69350 166757 6 io_in[24]
port 145 nsew signal input
rlabel metal2 s 72238 165957 72294 166757 6 io_in[25]
port 146 nsew signal input
rlabel metal2 s 75090 165957 75146 166757 6 io_in[26]
port 147 nsew signal input
rlabel metal2 s 77942 165957 77998 166757 6 io_in[27]
port 148 nsew signal input
rlabel metal2 s 80794 165957 80850 166757 6 io_in[28]
port 149 nsew signal input
rlabel metal2 s 83646 165957 83702 166757 6 io_in[29]
port 150 nsew signal input
rlabel metal2 s 6182 165957 6238 166757 6 io_in[2]
port 151 nsew signal input
rlabel metal2 s 86590 165957 86646 166757 6 io_in[30]
port 152 nsew signal input
rlabel metal2 s 89442 165957 89498 166757 6 io_in[31]
port 153 nsew signal input
rlabel metal2 s 92294 165957 92350 166757 6 io_in[32]
port 154 nsew signal input
rlabel metal2 s 95146 165957 95202 166757 6 io_in[33]
port 155 nsew signal input
rlabel metal2 s 97998 165957 98054 166757 6 io_in[34]
port 156 nsew signal input
rlabel metal2 s 100942 165957 100998 166757 6 io_in[35]
port 157 nsew signal input
rlabel metal2 s 103794 165957 103850 166757 6 io_in[36]
port 158 nsew signal input
rlabel metal2 s 106646 165957 106702 166757 6 io_in[37]
port 159 nsew signal input
rlabel metal2 s 9034 165957 9090 166757 6 io_in[3]
port 160 nsew signal input
rlabel metal2 s 11886 165957 11942 166757 6 io_in[4]
port 161 nsew signal input
rlabel metal2 s 14830 165957 14886 166757 6 io_in[5]
port 162 nsew signal input
rlabel metal2 s 17682 165957 17738 166757 6 io_in[6]
port 163 nsew signal input
rlabel metal2 s 20534 165957 20590 166757 6 io_in[7]
port 164 nsew signal input
rlabel metal2 s 23386 165957 23442 166757 6 io_in[8]
port 165 nsew signal input
rlabel metal2 s 26238 165957 26294 166757 6 io_in[9]
port 166 nsew signal input
rlabel metal2 s 1398 165957 1454 166757 6 io_oeb[0]
port 167 nsew signal output
rlabel metal2 s 30102 165957 30158 166757 6 io_oeb[10]
port 168 nsew signal output
rlabel metal2 s 32954 165957 33010 166757 6 io_oeb[11]
port 169 nsew signal output
rlabel metal2 s 35806 165957 35862 166757 6 io_oeb[12]
port 170 nsew signal output
rlabel metal2 s 38750 165957 38806 166757 6 io_oeb[13]
port 171 nsew signal output
rlabel metal2 s 41602 165957 41658 166757 6 io_oeb[14]
port 172 nsew signal output
rlabel metal2 s 44454 165957 44510 166757 6 io_oeb[15]
port 173 nsew signal output
rlabel metal2 s 47306 165957 47362 166757 6 io_oeb[16]
port 174 nsew signal output
rlabel metal2 s 50158 165957 50214 166757 6 io_oeb[17]
port 175 nsew signal output
rlabel metal2 s 53102 165957 53158 166757 6 io_oeb[18]
port 176 nsew signal output
rlabel metal2 s 55954 165957 56010 166757 6 io_oeb[19]
port 177 nsew signal output
rlabel metal2 s 4250 165957 4306 166757 6 io_oeb[1]
port 178 nsew signal output
rlabel metal2 s 58806 165957 58862 166757 6 io_oeb[20]
port 179 nsew signal output
rlabel metal2 s 61658 165957 61714 166757 6 io_oeb[21]
port 180 nsew signal output
rlabel metal2 s 64510 165957 64566 166757 6 io_oeb[22]
port 181 nsew signal output
rlabel metal2 s 67454 165957 67510 166757 6 io_oeb[23]
port 182 nsew signal output
rlabel metal2 s 70306 165957 70362 166757 6 io_oeb[24]
port 183 nsew signal output
rlabel metal2 s 73158 165957 73214 166757 6 io_oeb[25]
port 184 nsew signal output
rlabel metal2 s 76010 165957 76066 166757 6 io_oeb[26]
port 185 nsew signal output
rlabel metal2 s 78862 165957 78918 166757 6 io_oeb[27]
port 186 nsew signal output
rlabel metal2 s 81806 165957 81862 166757 6 io_oeb[28]
port 187 nsew signal output
rlabel metal2 s 84658 165957 84714 166757 6 io_oeb[29]
port 188 nsew signal output
rlabel metal2 s 7102 165957 7158 166757 6 io_oeb[2]
port 189 nsew signal output
rlabel metal2 s 87510 165957 87566 166757 6 io_oeb[30]
port 190 nsew signal output
rlabel metal2 s 90362 165957 90418 166757 6 io_oeb[31]
port 191 nsew signal output
rlabel metal2 s 93214 165957 93270 166757 6 io_oeb[32]
port 192 nsew signal output
rlabel metal2 s 96158 165957 96214 166757 6 io_oeb[33]
port 193 nsew signal output
rlabel metal2 s 99010 165957 99066 166757 6 io_oeb[34]
port 194 nsew signal output
rlabel metal2 s 101862 165957 101918 166757 6 io_oeb[35]
port 195 nsew signal output
rlabel metal2 s 104714 165957 104770 166757 6 io_oeb[36]
port 196 nsew signal output
rlabel metal2 s 107566 165957 107622 166757 6 io_oeb[37]
port 197 nsew signal output
rlabel metal2 s 10046 165957 10102 166757 6 io_oeb[3]
port 198 nsew signal output
rlabel metal2 s 12898 165957 12954 166757 6 io_oeb[4]
port 199 nsew signal output
rlabel metal2 s 15750 165957 15806 166757 6 io_oeb[5]
port 200 nsew signal output
rlabel metal2 s 18602 165957 18658 166757 6 io_oeb[6]
port 201 nsew signal output
rlabel metal2 s 21454 165957 21510 166757 6 io_oeb[7]
port 202 nsew signal output
rlabel metal2 s 24398 165957 24454 166757 6 io_oeb[8]
port 203 nsew signal output
rlabel metal2 s 27250 165957 27306 166757 6 io_oeb[9]
port 204 nsew signal output
rlabel metal2 s 2318 165957 2374 166757 6 io_out[0]
port 205 nsew signal output
rlabel metal2 s 31022 165957 31078 166757 6 io_out[10]
port 206 nsew signal output
rlabel metal2 s 33966 165957 34022 166757 6 io_out[11]
port 207 nsew signal output
rlabel metal2 s 36818 165957 36874 166757 6 io_out[12]
port 208 nsew signal output
rlabel metal2 s 39670 165957 39726 166757 6 io_out[13]
port 209 nsew signal output
rlabel metal2 s 42522 165957 42578 166757 6 io_out[14]
port 210 nsew signal output
rlabel metal2 s 45374 165957 45430 166757 6 io_out[15]
port 211 nsew signal output
rlabel metal2 s 48318 165957 48374 166757 6 io_out[16]
port 212 nsew signal output
rlabel metal2 s 51170 165957 51226 166757 6 io_out[17]
port 213 nsew signal output
rlabel metal2 s 54022 165957 54078 166757 6 io_out[18]
port 214 nsew signal output
rlabel metal2 s 56874 165957 56930 166757 6 io_out[19]
port 215 nsew signal output
rlabel metal2 s 5262 165957 5318 166757 6 io_out[1]
port 216 nsew signal output
rlabel metal2 s 59726 165957 59782 166757 6 io_out[20]
port 217 nsew signal output
rlabel metal2 s 62670 165957 62726 166757 6 io_out[21]
port 218 nsew signal output
rlabel metal2 s 65522 165957 65578 166757 6 io_out[22]
port 219 nsew signal output
rlabel metal2 s 68374 165957 68430 166757 6 io_out[23]
port 220 nsew signal output
rlabel metal2 s 71226 165957 71282 166757 6 io_out[24]
port 221 nsew signal output
rlabel metal2 s 74078 165957 74134 166757 6 io_out[25]
port 222 nsew signal output
rlabel metal2 s 77022 165957 77078 166757 6 io_out[26]
port 223 nsew signal output
rlabel metal2 s 79874 165957 79930 166757 6 io_out[27]
port 224 nsew signal output
rlabel metal2 s 82726 165957 82782 166757 6 io_out[28]
port 225 nsew signal output
rlabel metal2 s 85578 165957 85634 166757 6 io_out[29]
port 226 nsew signal output
rlabel metal2 s 8114 165957 8170 166757 6 io_out[2]
port 227 nsew signal output
rlabel metal2 s 88430 165957 88486 166757 6 io_out[30]
port 228 nsew signal output
rlabel metal2 s 91374 165957 91430 166757 6 io_out[31]
port 229 nsew signal output
rlabel metal2 s 94226 165957 94282 166757 6 io_out[32]
port 230 nsew signal output
rlabel metal2 s 97078 165957 97134 166757 6 io_out[33]
port 231 nsew signal output
rlabel metal2 s 99930 165957 99986 166757 6 io_out[34]
port 232 nsew signal output
rlabel metal2 s 102782 165957 102838 166757 6 io_out[35]
port 233 nsew signal output
rlabel metal2 s 105726 165957 105782 166757 6 io_out[36]
port 234 nsew signal output
rlabel metal2 s 108578 165957 108634 166757 6 io_out[37]
port 235 nsew signal output
rlabel metal2 s 10966 165957 11022 166757 6 io_out[3]
port 236 nsew signal output
rlabel metal2 s 13818 165957 13874 166757 6 io_out[4]
port 237 nsew signal output
rlabel metal2 s 16670 165957 16726 166757 6 io_out[5]
port 238 nsew signal output
rlabel metal2 s 19614 165957 19670 166757 6 io_out[6]
port 239 nsew signal output
rlabel metal2 s 22466 165957 22522 166757 6 io_out[7]
port 240 nsew signal output
rlabel metal2 s 25318 165957 25374 166757 6 io_out[8]
port 241 nsew signal output
rlabel metal2 s 28170 165957 28226 166757 6 io_out[9]
port 242 nsew signal output
rlabel metal2 s 107474 0 107530 800 6 irq[0]
port 243 nsew signal output
rlabel metal2 s 108486 0 108542 800 6 irq[1]
port 244 nsew signal output
rlabel metal2 s 109498 0 109554 800 6 irq[2]
port 245 nsew signal output
rlabel metal2 s 112534 0 112590 800 6 o_addr1[0]
port 246 nsew signal output
rlabel metal3 s 163813 12792 164613 12912 6 o_addr1[1]
port 247 nsew signal output
rlabel metal2 s 123666 0 123722 800 6 o_addr1[2]
port 248 nsew signal output
rlabel metal2 s 127622 0 127678 800 6 o_addr1[3]
port 249 nsew signal output
rlabel metal3 s 0 35776 800 35896 6 o_addr1[4]
port 250 nsew signal output
rlabel metal2 s 122930 165957 122986 166757 6 o_addr1[5]
port 251 nsew signal output
rlabel metal3 s 0 47336 800 47456 6 o_addr1[6]
port 252 nsew signal output
rlabel metal3 s 163813 64608 164613 64728 6 o_addr1[7]
port 253 nsew signal output
rlabel metal2 s 130566 165957 130622 166757 6 o_addr1[8]
port 254 nsew signal output
rlabel metal3 s 0 8032 800 8152 6 o_addr1_1[0]
port 255 nsew signal output
rlabel metal2 s 113362 165957 113418 166757 6 o_addr1_1[1]
port 256 nsew signal output
rlabel metal3 s 0 17280 800 17400 6 o_addr1_1[2]
port 257 nsew signal output
rlabel metal2 s 126610 0 126666 800 6 o_addr1_1[3]
port 258 nsew signal output
rlabel metal3 s 163813 38632 164613 38752 6 o_addr1_1[4]
port 259 nsew signal output
rlabel metal3 s 0 42712 800 42832 6 o_addr1_1[5]
port 260 nsew signal output
rlabel metal3 s 163813 58760 164613 58880 6 o_addr1_1[6]
port 261 nsew signal output
rlabel metal2 s 126702 165957 126758 166757 6 o_addr1_1[7]
port 262 nsew signal output
rlabel metal2 s 135718 0 135774 800 6 o_addr1_1[8]
port 263 nsew signal output
rlabel metal3 s 163813 1368 164613 1488 6 o_csb0
port 264 nsew signal output
rlabel metal2 s 110510 0 110566 800 6 o_csb0_1
port 265 nsew signal output
rlabel metal2 s 109498 165957 109554 166757 6 o_csb1
port 266 nsew signal output
rlabel metal3 s 0 1096 800 1216 6 o_csb1_1
port 267 nsew signal output
rlabel metal2 s 113546 0 113602 800 6 o_din0[0]
port 268 nsew signal output
rlabel metal3 s 0 72768 800 72888 6 o_din0[10]
port 269 nsew signal output
rlabel metal3 s 0 79704 800 79824 6 o_din0[11]
port 270 nsew signal output
rlabel metal3 s 163813 84736 164613 84856 6 o_din0[12]
port 271 nsew signal output
rlabel metal2 s 140134 165957 140190 166757 6 o_din0[13]
port 272 nsew signal output
rlabel metal2 s 141054 165957 141110 166757 6 o_din0[14]
port 273 nsew signal output
rlabel metal3 s 0 93712 800 93832 6 o_din0[15]
port 274 nsew signal output
rlabel metal2 s 145838 165957 145894 166757 6 o_din0[16]
port 275 nsew signal output
rlabel metal3 s 163813 107720 164613 107840 6 o_din0[17]
port 276 nsew signal output
rlabel metal2 s 147862 0 147918 800 6 o_din0[18]
port 277 nsew signal output
rlabel metal2 s 149702 165957 149758 166757 6 o_din0[19]
port 278 nsew signal output
rlabel metal2 s 118606 0 118662 800 6 o_din0[1]
port 279 nsew signal output
rlabel metal3 s 163813 127848 164613 127968 6 o_din0[20]
port 280 nsew signal output
rlabel metal2 s 149886 0 149942 800 6 o_din0[21]
port 281 nsew signal output
rlabel metal3 s 0 123768 800 123888 6 o_din0[22]
port 282 nsew signal output
rlabel metal3 s 0 128392 800 128512 6 o_din0[23]
port 283 nsew signal output
rlabel metal2 s 154486 165957 154542 166757 6 o_din0[24]
port 284 nsew signal output
rlabel metal2 s 157338 165957 157394 166757 6 o_din0[25]
port 285 nsew signal output
rlabel metal3 s 163813 153688 164613 153808 6 o_din0[26]
port 286 nsew signal output
rlabel metal2 s 159270 165957 159326 166757 6 o_din0[27]
port 287 nsew signal output
rlabel metal3 s 0 149200 800 149320 6 o_din0[28]
port 288 nsew signal output
rlabel metal3 s 0 153824 800 153944 6 o_din0[29]
port 289 nsew signal output
rlabel metal3 s 163813 21360 164613 21480 6 o_din0[2]
port 290 nsew signal output
rlabel metal2 s 162030 0 162086 800 6 o_din0[30]
port 291 nsew signal output
rlabel metal2 s 164054 165957 164110 166757 6 o_din0[31]
port 292 nsew signal output
rlabel metal3 s 163813 27208 164613 27328 6 o_din0[3]
port 293 nsew signal output
rlabel metal2 s 120078 165957 120134 166757 6 o_din0[4]
port 294 nsew signal output
rlabel metal2 s 130658 0 130714 800 6 o_din0[5]
port 295 nsew signal output
rlabel metal2 s 124862 165957 124918 166757 6 o_din0[6]
port 296 nsew signal output
rlabel metal3 s 0 61208 800 61328 6 o_din0[7]
port 297 nsew signal output
rlabel metal2 s 131486 165957 131542 166757 6 o_din0[8]
port 298 nsew signal output
rlabel metal3 s 0 70456 800 70576 6 o_din0[9]
port 299 nsew signal output
rlabel metal3 s 0 10344 800 10464 6 o_din0_1[0]
port 300 nsew signal output
rlabel metal2 s 136730 0 136786 800 6 o_din0_1[10]
port 301 nsew signal output
rlabel metal2 s 138754 0 138810 800 6 o_din0_1[11]
port 302 nsew signal output
rlabel metal2 s 139766 0 139822 800 6 o_din0_1[12]
port 303 nsew signal output
rlabel metal2 s 139214 165957 139270 166757 6 o_din0_1[13]
port 304 nsew signal output
rlabel metal3 s 0 89088 800 89208 6 o_din0_1[14]
port 305 nsew signal output
rlabel metal2 s 145838 0 145894 800 6 o_din0_1[15]
port 306 nsew signal output
rlabel metal2 s 144918 165957 144974 166757 6 o_din0_1[16]
port 307 nsew signal output
rlabel metal3 s 163813 104728 164613 104848 6 o_din0_1[17]
port 308 nsew signal output
rlabel metal2 s 147770 165957 147826 166757 6 o_din0_1[18]
port 309 nsew signal output
rlabel metal3 s 0 107584 800 107704 6 o_din0_1[19]
port 310 nsew signal output
rlabel metal2 s 117594 0 117650 800 6 o_din0_1[1]
port 311 nsew signal output
rlabel metal2 s 150622 165957 150678 166757 6 o_din0_1[20]
port 312 nsew signal output
rlabel metal3 s 0 116832 800 116952 6 o_din0_1[21]
port 313 nsew signal output
rlabel metal3 s 0 121456 800 121576 6 o_din0_1[22]
port 314 nsew signal output
rlabel metal3 s 163813 136416 164613 136536 6 o_din0_1[23]
port 315 nsew signal output
rlabel metal3 s 0 130704 800 130824 6 o_din0_1[24]
port 316 nsew signal output
rlabel metal2 s 156418 165957 156474 166757 6 o_din0_1[25]
port 317 nsew signal output
rlabel metal3 s 0 137640 800 137760 6 o_din0_1[26]
port 318 nsew signal output
rlabel metal2 s 158350 165957 158406 166757 6 o_din0_1[27]
port 319 nsew signal output
rlabel metal3 s 0 146888 800 147008 6 o_din0_1[28]
port 320 nsew signal output
rlabel metal2 s 162122 165957 162178 166757 6 o_din0_1[29]
port 321 nsew signal output
rlabel metal3 s 163813 18504 164613 18624 6 o_din0_1[2]
port 322 nsew signal output
rlabel metal3 s 163813 165112 164613 165232 6 o_din0_1[30]
port 323 nsew signal output
rlabel metal2 s 164054 0 164110 800 6 o_din0_1[31]
port 324 nsew signal output
rlabel metal2 s 118146 165957 118202 166757 6 o_din0_1[3]
port 325 nsew signal output
rlabel metal2 s 119066 165957 119122 166757 6 o_din0_1[4]
port 326 nsew signal output
rlabel metal3 s 163813 47336 164613 47456 6 o_din0_1[5]
port 327 nsew signal output
rlabel metal3 s 0 49648 800 49768 6 o_din0_1[6]
port 328 nsew signal output
rlabel metal3 s 0 58896 800 59016 6 o_din0_1[7]
port 329 nsew signal output
rlabel metal3 s 163813 70320 164613 70440 6 o_din0_1[8]
port 330 nsew signal output
rlabel metal3 s 0 68144 800 68264 6 o_din0_1[9]
port 331 nsew signal output
rlabel metal3 s 163813 7080 164613 7200 6 o_waddr0[0]
port 332 nsew signal output
rlabel metal2 s 115294 165957 115350 166757 6 o_waddr0[1]
port 333 nsew signal output
rlabel metal2 s 124586 0 124642 800 6 o_waddr0[2]
port 334 nsew signal output
rlabel metal3 s 163813 30064 164613 30184 6 o_waddr0[3]
port 335 nsew signal output
rlabel metal3 s 163813 44480 164613 44600 6 o_waddr0[4]
port 336 nsew signal output
rlabel metal3 s 163813 53048 164613 53168 6 o_waddr0[5]
port 337 nsew signal output
rlabel metal3 s 0 51960 800 52080 6 o_waddr0[6]
port 338 nsew signal output
rlabel metal3 s 163813 67464 164613 67584 6 o_waddr0[7]
port 339 nsew signal output
rlabel metal3 s 0 63520 800 63640 6 o_waddr0[8]
port 340 nsew signal output
rlabel metal2 s 114558 0 114614 800 6 o_waddr0_1[0]
port 341 nsew signal output
rlabel metal2 s 114282 165957 114338 166757 6 o_waddr0_1[1]
port 342 nsew signal output
rlabel metal3 s 0 19592 800 19712 6 o_waddr0_1[2]
port 343 nsew signal output
rlabel metal2 s 128634 0 128690 800 6 o_waddr0_1[3]
port 344 nsew signal output
rlabel metal3 s 163813 41488 164613 41608 6 o_waddr0_1[4]
port 345 nsew signal output
rlabel metal3 s 163813 50192 164613 50312 6 o_waddr0_1[5]
port 346 nsew signal output
rlabel metal2 s 132682 0 132738 800 6 o_waddr0_1[6]
port 347 nsew signal output
rlabel metal2 s 133694 0 133750 800 6 o_waddr0_1[7]
port 348 nsew signal output
rlabel metal3 s 163813 73176 164613 73296 6 o_waddr0_1[8]
port 349 nsew signal output
rlabel metal3 s 0 3408 800 3528 6 o_web0
port 350 nsew signal output
rlabel metal2 s 111522 0 111578 800 6 o_web0_1
port 351 nsew signal output
rlabel metal2 s 115570 0 115626 800 6 o_wmask0[0]
port 352 nsew signal output
rlabel metal2 s 120630 0 120686 800 6 o_wmask0[1]
port 353 nsew signal output
rlabel metal2 s 117134 165957 117190 166757 6 o_wmask0[2]
port 354 nsew signal output
rlabel metal3 s 0 31152 800 31272 6 o_wmask0[3]
port 355 nsew signal output
rlabel metal2 s 116582 0 116638 800 6 o_wmask0_1[0]
port 356 nsew signal output
rlabel metal2 s 119618 0 119674 800 6 o_wmask0_1[1]
port 357 nsew signal output
rlabel metal3 s 0 21904 800 22024 6 o_wmask0_1[2]
port 358 nsew signal output
rlabel metal3 s 0 28840 800 28960 6 o_wmask0_1[3]
port 359 nsew signal output
rlabel metal4 s 4208 2128 4528 164336 6 vccd1
port 360 nsew power input
rlabel metal4 s 34928 2128 35248 164336 6 vccd1
port 360 nsew power input
rlabel metal4 s 65648 2128 65968 164336 6 vccd1
port 360 nsew power input
rlabel metal4 s 96368 2128 96688 164336 6 vccd1
port 360 nsew power input
rlabel metal4 s 127088 2128 127408 164336 6 vccd1
port 360 nsew power input
rlabel metal4 s 157808 2128 158128 164336 6 vccd1
port 360 nsew power input
rlabel metal4 s 19568 2128 19888 164336 6 vssd1
port 361 nsew ground input
rlabel metal4 s 50288 2128 50608 164336 6 vssd1
port 361 nsew ground input
rlabel metal4 s 81008 2128 81328 164336 6 vssd1
port 361 nsew ground input
rlabel metal4 s 111728 2128 112048 164336 6 vssd1
port 361 nsew ground input
rlabel metal4 s 142448 2128 142768 164336 6 vssd1
port 361 nsew ground input
rlabel metal2 s 478 0 534 800 6 wb_clk_i
port 362 nsew signal input
rlabel metal2 s 1398 0 1454 800 6 wb_rst_i
port 363 nsew signal input
rlabel metal2 s 2410 0 2466 800 6 wbs_ack_o
port 364 nsew signal output
rlabel metal2 s 6458 0 6514 800 6 wbs_adr_i[0]
port 365 nsew signal input
rlabel metal2 s 40866 0 40922 800 6 wbs_adr_i[10]
port 366 nsew signal input
rlabel metal2 s 43810 0 43866 800 6 wbs_adr_i[11]
port 367 nsew signal input
rlabel metal2 s 46846 0 46902 800 6 wbs_adr_i[12]
port 368 nsew signal input
rlabel metal2 s 49882 0 49938 800 6 wbs_adr_i[13]
port 369 nsew signal input
rlabel metal2 s 52918 0 52974 800 6 wbs_adr_i[14]
port 370 nsew signal input
rlabel metal2 s 55954 0 56010 800 6 wbs_adr_i[15]
port 371 nsew signal input
rlabel metal2 s 58990 0 59046 800 6 wbs_adr_i[16]
port 372 nsew signal input
rlabel metal2 s 62026 0 62082 800 6 wbs_adr_i[17]
port 373 nsew signal input
rlabel metal2 s 65062 0 65118 800 6 wbs_adr_i[18]
port 374 nsew signal input
rlabel metal2 s 68098 0 68154 800 6 wbs_adr_i[19]
port 375 nsew signal input
rlabel metal2 s 10506 0 10562 800 6 wbs_adr_i[1]
port 376 nsew signal input
rlabel metal2 s 71134 0 71190 800 6 wbs_adr_i[20]
port 377 nsew signal input
rlabel metal2 s 74170 0 74226 800 6 wbs_adr_i[21]
port 378 nsew signal input
rlabel metal2 s 77206 0 77262 800 6 wbs_adr_i[22]
port 379 nsew signal input
rlabel metal2 s 80242 0 80298 800 6 wbs_adr_i[23]
port 380 nsew signal input
rlabel metal2 s 83186 0 83242 800 6 wbs_adr_i[24]
port 381 nsew signal input
rlabel metal2 s 86222 0 86278 800 6 wbs_adr_i[25]
port 382 nsew signal input
rlabel metal2 s 89258 0 89314 800 6 wbs_adr_i[26]
port 383 nsew signal input
rlabel metal2 s 92294 0 92350 800 6 wbs_adr_i[27]
port 384 nsew signal input
rlabel metal2 s 95330 0 95386 800 6 wbs_adr_i[28]
port 385 nsew signal input
rlabel metal2 s 98366 0 98422 800 6 wbs_adr_i[29]
port 386 nsew signal input
rlabel metal2 s 14554 0 14610 800 6 wbs_adr_i[2]
port 387 nsew signal input
rlabel metal2 s 101402 0 101458 800 6 wbs_adr_i[30]
port 388 nsew signal input
rlabel metal2 s 104438 0 104494 800 6 wbs_adr_i[31]
port 389 nsew signal input
rlabel metal2 s 18602 0 18658 800 6 wbs_adr_i[3]
port 390 nsew signal input
rlabel metal2 s 22650 0 22706 800 6 wbs_adr_i[4]
port 391 nsew signal input
rlabel metal2 s 25686 0 25742 800 6 wbs_adr_i[5]
port 392 nsew signal input
rlabel metal2 s 28722 0 28778 800 6 wbs_adr_i[6]
port 393 nsew signal input
rlabel metal2 s 31758 0 31814 800 6 wbs_adr_i[7]
port 394 nsew signal input
rlabel metal2 s 34794 0 34850 800 6 wbs_adr_i[8]
port 395 nsew signal input
rlabel metal2 s 37830 0 37886 800 6 wbs_adr_i[9]
port 396 nsew signal input
rlabel metal2 s 3422 0 3478 800 6 wbs_cyc_i
port 397 nsew signal input
rlabel metal2 s 7470 0 7526 800 6 wbs_dat_i[0]
port 398 nsew signal input
rlabel metal2 s 41786 0 41842 800 6 wbs_dat_i[10]
port 399 nsew signal input
rlabel metal2 s 44822 0 44878 800 6 wbs_dat_i[11]
port 400 nsew signal input
rlabel metal2 s 47858 0 47914 800 6 wbs_dat_i[12]
port 401 nsew signal input
rlabel metal2 s 50894 0 50950 800 6 wbs_dat_i[13]
port 402 nsew signal input
rlabel metal2 s 53930 0 53986 800 6 wbs_dat_i[14]
port 403 nsew signal input
rlabel metal2 s 56966 0 57022 800 6 wbs_dat_i[15]
port 404 nsew signal input
rlabel metal2 s 60002 0 60058 800 6 wbs_dat_i[16]
port 405 nsew signal input
rlabel metal2 s 63038 0 63094 800 6 wbs_dat_i[17]
port 406 nsew signal input
rlabel metal2 s 66074 0 66130 800 6 wbs_dat_i[18]
port 407 nsew signal input
rlabel metal2 s 69110 0 69166 800 6 wbs_dat_i[19]
port 408 nsew signal input
rlabel metal2 s 11518 0 11574 800 6 wbs_dat_i[1]
port 409 nsew signal input
rlabel metal2 s 72146 0 72202 800 6 wbs_dat_i[20]
port 410 nsew signal input
rlabel metal2 s 75182 0 75238 800 6 wbs_dat_i[21]
port 411 nsew signal input
rlabel metal2 s 78218 0 78274 800 6 wbs_dat_i[22]
port 412 nsew signal input
rlabel metal2 s 81254 0 81310 800 6 wbs_dat_i[23]
port 413 nsew signal input
rlabel metal2 s 84198 0 84254 800 6 wbs_dat_i[24]
port 414 nsew signal input
rlabel metal2 s 87234 0 87290 800 6 wbs_dat_i[25]
port 415 nsew signal input
rlabel metal2 s 90270 0 90326 800 6 wbs_dat_i[26]
port 416 nsew signal input
rlabel metal2 s 93306 0 93362 800 6 wbs_dat_i[27]
port 417 nsew signal input
rlabel metal2 s 96342 0 96398 800 6 wbs_dat_i[28]
port 418 nsew signal input
rlabel metal2 s 99378 0 99434 800 6 wbs_dat_i[29]
port 419 nsew signal input
rlabel metal2 s 15566 0 15622 800 6 wbs_dat_i[2]
port 420 nsew signal input
rlabel metal2 s 102414 0 102470 800 6 wbs_dat_i[30]
port 421 nsew signal input
rlabel metal2 s 105450 0 105506 800 6 wbs_dat_i[31]
port 422 nsew signal input
rlabel metal2 s 19614 0 19670 800 6 wbs_dat_i[3]
port 423 nsew signal input
rlabel metal2 s 23662 0 23718 800 6 wbs_dat_i[4]
port 424 nsew signal input
rlabel metal2 s 26698 0 26754 800 6 wbs_dat_i[5]
port 425 nsew signal input
rlabel metal2 s 29734 0 29790 800 6 wbs_dat_i[6]
port 426 nsew signal input
rlabel metal2 s 32770 0 32826 800 6 wbs_dat_i[7]
port 427 nsew signal input
rlabel metal2 s 35806 0 35862 800 6 wbs_dat_i[8]
port 428 nsew signal input
rlabel metal2 s 38842 0 38898 800 6 wbs_dat_i[9]
port 429 nsew signal input
rlabel metal2 s 8482 0 8538 800 6 wbs_dat_o[0]
port 430 nsew signal output
rlabel metal2 s 42798 0 42854 800 6 wbs_dat_o[10]
port 431 nsew signal output
rlabel metal2 s 45834 0 45890 800 6 wbs_dat_o[11]
port 432 nsew signal output
rlabel metal2 s 48870 0 48926 800 6 wbs_dat_o[12]
port 433 nsew signal output
rlabel metal2 s 51906 0 51962 800 6 wbs_dat_o[13]
port 434 nsew signal output
rlabel metal2 s 54942 0 54998 800 6 wbs_dat_o[14]
port 435 nsew signal output
rlabel metal2 s 57978 0 58034 800 6 wbs_dat_o[15]
port 436 nsew signal output
rlabel metal2 s 61014 0 61070 800 6 wbs_dat_o[16]
port 437 nsew signal output
rlabel metal2 s 64050 0 64106 800 6 wbs_dat_o[17]
port 438 nsew signal output
rlabel metal2 s 67086 0 67142 800 6 wbs_dat_o[18]
port 439 nsew signal output
rlabel metal2 s 70122 0 70178 800 6 wbs_dat_o[19]
port 440 nsew signal output
rlabel metal2 s 12530 0 12586 800 6 wbs_dat_o[1]
port 441 nsew signal output
rlabel metal2 s 73158 0 73214 800 6 wbs_dat_o[20]
port 442 nsew signal output
rlabel metal2 s 76194 0 76250 800 6 wbs_dat_o[21]
port 443 nsew signal output
rlabel metal2 s 79230 0 79286 800 6 wbs_dat_o[22]
port 444 nsew signal output
rlabel metal2 s 82266 0 82322 800 6 wbs_dat_o[23]
port 445 nsew signal output
rlabel metal2 s 85210 0 85266 800 6 wbs_dat_o[24]
port 446 nsew signal output
rlabel metal2 s 88246 0 88302 800 6 wbs_dat_o[25]
port 447 nsew signal output
rlabel metal2 s 91282 0 91338 800 6 wbs_dat_o[26]
port 448 nsew signal output
rlabel metal2 s 94318 0 94374 800 6 wbs_dat_o[27]
port 449 nsew signal output
rlabel metal2 s 97354 0 97410 800 6 wbs_dat_o[28]
port 450 nsew signal output
rlabel metal2 s 100390 0 100446 800 6 wbs_dat_o[29]
port 451 nsew signal output
rlabel metal2 s 16578 0 16634 800 6 wbs_dat_o[2]
port 452 nsew signal output
rlabel metal2 s 103426 0 103482 800 6 wbs_dat_o[30]
port 453 nsew signal output
rlabel metal2 s 106462 0 106518 800 6 wbs_dat_o[31]
port 454 nsew signal output
rlabel metal2 s 20626 0 20682 800 6 wbs_dat_o[3]
port 455 nsew signal output
rlabel metal2 s 24674 0 24730 800 6 wbs_dat_o[4]
port 456 nsew signal output
rlabel metal2 s 27710 0 27766 800 6 wbs_dat_o[5]
port 457 nsew signal output
rlabel metal2 s 30746 0 30802 800 6 wbs_dat_o[6]
port 458 nsew signal output
rlabel metal2 s 33782 0 33838 800 6 wbs_dat_o[7]
port 459 nsew signal output
rlabel metal2 s 36818 0 36874 800 6 wbs_dat_o[8]
port 460 nsew signal output
rlabel metal2 s 39854 0 39910 800 6 wbs_dat_o[9]
port 461 nsew signal output
rlabel metal2 s 9494 0 9550 800 6 wbs_sel_i[0]
port 462 nsew signal input
rlabel metal2 s 13542 0 13598 800 6 wbs_sel_i[1]
port 463 nsew signal input
rlabel metal2 s 17590 0 17646 800 6 wbs_sel_i[2]
port 464 nsew signal input
rlabel metal2 s 21638 0 21694 800 6 wbs_sel_i[3]
port 465 nsew signal input
rlabel metal2 s 4434 0 4490 800 6 wbs_stb_i
port 466 nsew signal input
rlabel metal2 s 5446 0 5502 800 6 wbs_we_i
port 467 nsew signal input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 164613 166757
string LEFview TRUE
string GDS_FILE /local/caravel_user_project/openlane/user_proj/runs/user_proj/results/magic/user_proj.gds
string GDS_END 80001714
string GDS_START 1385536
<< end >>

