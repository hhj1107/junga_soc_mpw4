magic
tech sky130A
magscale 1 2
timestamp 1640400942
<< obsli1 >>
rect 857 2159 164191 164305
<< obsm1 >>
rect 290 8 164206 164336
<< metal2 >>
rect 386 165721 442 166521
rect 1214 165721 1270 166521
rect 2134 165721 2190 166521
rect 3054 165721 3110 166521
rect 3974 165721 4030 166521
rect 4894 165721 4950 166521
rect 5814 165721 5870 166521
rect 6734 165721 6790 166521
rect 7562 165721 7618 166521
rect 8482 165721 8538 166521
rect 9402 165721 9458 166521
rect 10322 165721 10378 166521
rect 11242 165721 11298 166521
rect 12162 165721 12218 166521
rect 13082 165721 13138 166521
rect 14002 165721 14058 166521
rect 14830 165721 14886 166521
rect 15750 165721 15806 166521
rect 16670 165721 16726 166521
rect 17590 165721 17646 166521
rect 18510 165721 18566 166521
rect 19430 165721 19486 166521
rect 20350 165721 20406 166521
rect 21270 165721 21326 166521
rect 22098 165721 22154 166521
rect 23018 165721 23074 166521
rect 23938 165721 23994 166521
rect 24858 165721 24914 166521
rect 25778 165721 25834 166521
rect 26698 165721 26754 166521
rect 27618 165721 27674 166521
rect 28538 165721 28594 166521
rect 29366 165721 29422 166521
rect 30286 165721 30342 166521
rect 31206 165721 31262 166521
rect 32126 165721 32182 166521
rect 33046 165721 33102 166521
rect 33966 165721 34022 166521
rect 34886 165721 34942 166521
rect 35806 165721 35862 166521
rect 36634 165721 36690 166521
rect 37554 165721 37610 166521
rect 38474 165721 38530 166521
rect 39394 165721 39450 166521
rect 40314 165721 40370 166521
rect 41234 165721 41290 166521
rect 42154 165721 42210 166521
rect 43074 165721 43130 166521
rect 43902 165721 43958 166521
rect 44822 165721 44878 166521
rect 45742 165721 45798 166521
rect 46662 165721 46718 166521
rect 47582 165721 47638 166521
rect 48502 165721 48558 166521
rect 49422 165721 49478 166521
rect 50342 165721 50398 166521
rect 51170 165721 51226 166521
rect 52090 165721 52146 166521
rect 53010 165721 53066 166521
rect 53930 165721 53986 166521
rect 54850 165721 54906 166521
rect 55770 165721 55826 166521
rect 56690 165721 56746 166521
rect 57518 165721 57574 166521
rect 58438 165721 58494 166521
rect 59358 165721 59414 166521
rect 60278 165721 60334 166521
rect 61198 165721 61254 166521
rect 62118 165721 62174 166521
rect 63038 165721 63094 166521
rect 63958 165721 64014 166521
rect 64786 165721 64842 166521
rect 65706 165721 65762 166521
rect 66626 165721 66682 166521
rect 67546 165721 67602 166521
rect 68466 165721 68522 166521
rect 69386 165721 69442 166521
rect 70306 165721 70362 166521
rect 71226 165721 71282 166521
rect 72054 165721 72110 166521
rect 72974 165721 73030 166521
rect 73894 165721 73950 166521
rect 74814 165721 74870 166521
rect 75734 165721 75790 166521
rect 76654 165721 76710 166521
rect 77574 165721 77630 166521
rect 78494 165721 78550 166521
rect 79322 165721 79378 166521
rect 80242 165721 80298 166521
rect 81162 165721 81218 166521
rect 82082 165721 82138 166521
rect 83002 165721 83058 166521
rect 83922 165721 83978 166521
rect 84842 165721 84898 166521
rect 85762 165721 85818 166521
rect 86590 165721 86646 166521
rect 87510 165721 87566 166521
rect 88430 165721 88486 166521
rect 89350 165721 89406 166521
rect 90270 165721 90326 166521
rect 91190 165721 91246 166521
rect 92110 165721 92166 166521
rect 93030 165721 93086 166521
rect 93858 165721 93914 166521
rect 94778 165721 94834 166521
rect 95698 165721 95754 166521
rect 96618 165721 96674 166521
rect 97538 165721 97594 166521
rect 98458 165721 98514 166521
rect 99378 165721 99434 166521
rect 100298 165721 100354 166521
rect 101126 165721 101182 166521
rect 102046 165721 102102 166521
rect 102966 165721 103022 166521
rect 103886 165721 103942 166521
rect 104806 165721 104862 166521
rect 105726 165721 105782 166521
rect 106646 165721 106702 166521
rect 107566 165721 107622 166521
rect 108394 165721 108450 166521
rect 109314 165721 109370 166521
rect 110234 165721 110290 166521
rect 111154 165721 111210 166521
rect 112074 165721 112130 166521
rect 112994 165721 113050 166521
rect 113914 165721 113970 166521
rect 114742 165721 114798 166521
rect 115662 165721 115718 166521
rect 116582 165721 116638 166521
rect 117502 165721 117558 166521
rect 118422 165721 118478 166521
rect 119342 165721 119398 166521
rect 120262 165721 120318 166521
rect 121182 165721 121238 166521
rect 122010 165721 122066 166521
rect 122930 165721 122986 166521
rect 123850 165721 123906 166521
rect 124770 165721 124826 166521
rect 125690 165721 125746 166521
rect 126610 165721 126666 166521
rect 127530 165721 127586 166521
rect 128450 165721 128506 166521
rect 129278 165721 129334 166521
rect 130198 165721 130254 166521
rect 131118 165721 131174 166521
rect 132038 165721 132094 166521
rect 132958 165721 133014 166521
rect 133878 165721 133934 166521
rect 134798 165721 134854 166521
rect 135718 165721 135774 166521
rect 136546 165721 136602 166521
rect 137466 165721 137522 166521
rect 138386 165721 138442 166521
rect 139306 165721 139362 166521
rect 140226 165721 140282 166521
rect 141146 165721 141202 166521
rect 142066 165721 142122 166521
rect 142986 165721 143042 166521
rect 143814 165721 143870 166521
rect 144734 165721 144790 166521
rect 145654 165721 145710 166521
rect 146574 165721 146630 166521
rect 147494 165721 147550 166521
rect 148414 165721 148470 166521
rect 149334 165721 149390 166521
rect 150254 165721 150310 166521
rect 151082 165721 151138 166521
rect 152002 165721 152058 166521
rect 152922 165721 152978 166521
rect 153842 165721 153898 166521
rect 154762 165721 154818 166521
rect 155682 165721 155738 166521
rect 156602 165721 156658 166521
rect 157522 165721 157578 166521
rect 158350 165721 158406 166521
rect 159270 165721 159326 166521
rect 160190 165721 160246 166521
rect 161110 165721 161166 166521
rect 162030 165721 162086 166521
rect 162950 165721 163006 166521
rect 163870 165721 163926 166521
rect 478 0 534 800
rect 1398 0 1454 800
rect 2318 0 2374 800
rect 3238 0 3294 800
rect 4158 0 4214 800
rect 5170 0 5226 800
rect 6090 0 6146 800
rect 7010 0 7066 800
rect 7930 0 7986 800
rect 8850 0 8906 800
rect 9862 0 9918 800
rect 10782 0 10838 800
rect 11702 0 11758 800
rect 12622 0 12678 800
rect 13542 0 13598 800
rect 14554 0 14610 800
rect 15474 0 15530 800
rect 16394 0 16450 800
rect 17314 0 17370 800
rect 18326 0 18382 800
rect 19246 0 19302 800
rect 20166 0 20222 800
rect 21086 0 21142 800
rect 22006 0 22062 800
rect 23018 0 23074 800
rect 23938 0 23994 800
rect 24858 0 24914 800
rect 25778 0 25834 800
rect 26698 0 26754 800
rect 27710 0 27766 800
rect 28630 0 28686 800
rect 29550 0 29606 800
rect 30470 0 30526 800
rect 31390 0 31446 800
rect 32402 0 32458 800
rect 33322 0 33378 800
rect 34242 0 34298 800
rect 35162 0 35218 800
rect 36174 0 36230 800
rect 37094 0 37150 800
rect 38014 0 38070 800
rect 38934 0 38990 800
rect 39854 0 39910 800
rect 40866 0 40922 800
rect 41786 0 41842 800
rect 42706 0 42762 800
rect 43626 0 43682 800
rect 44546 0 44602 800
rect 45558 0 45614 800
rect 46478 0 46534 800
rect 47398 0 47454 800
rect 48318 0 48374 800
rect 49238 0 49294 800
rect 50250 0 50306 800
rect 51170 0 51226 800
rect 52090 0 52146 800
rect 53010 0 53066 800
rect 54022 0 54078 800
rect 54942 0 54998 800
rect 55862 0 55918 800
rect 56782 0 56838 800
rect 57702 0 57758 800
rect 58714 0 58770 800
rect 59634 0 59690 800
rect 60554 0 60610 800
rect 61474 0 61530 800
rect 62394 0 62450 800
rect 63406 0 63462 800
rect 64326 0 64382 800
rect 65246 0 65302 800
rect 66166 0 66222 800
rect 67178 0 67234 800
rect 68098 0 68154 800
rect 69018 0 69074 800
rect 69938 0 69994 800
rect 70858 0 70914 800
rect 71870 0 71926 800
rect 72790 0 72846 800
rect 73710 0 73766 800
rect 74630 0 74686 800
rect 75550 0 75606 800
rect 76562 0 76618 800
rect 77482 0 77538 800
rect 78402 0 78458 800
rect 79322 0 79378 800
rect 80242 0 80298 800
rect 81254 0 81310 800
rect 82174 0 82230 800
rect 83094 0 83150 800
rect 84014 0 84070 800
rect 85026 0 85082 800
rect 85946 0 86002 800
rect 86866 0 86922 800
rect 87786 0 87842 800
rect 88706 0 88762 800
rect 89718 0 89774 800
rect 90638 0 90694 800
rect 91558 0 91614 800
rect 92478 0 92534 800
rect 93398 0 93454 800
rect 94410 0 94466 800
rect 95330 0 95386 800
rect 96250 0 96306 800
rect 97170 0 97226 800
rect 98090 0 98146 800
rect 99102 0 99158 800
rect 100022 0 100078 800
rect 100942 0 100998 800
rect 101862 0 101918 800
rect 102874 0 102930 800
rect 103794 0 103850 800
rect 104714 0 104770 800
rect 105634 0 105690 800
rect 106554 0 106610 800
rect 107566 0 107622 800
rect 108486 0 108542 800
rect 109406 0 109462 800
rect 110326 0 110382 800
rect 111246 0 111302 800
rect 112258 0 112314 800
rect 113178 0 113234 800
rect 114098 0 114154 800
rect 115018 0 115074 800
rect 116030 0 116086 800
rect 116950 0 117006 800
rect 117870 0 117926 800
rect 118790 0 118846 800
rect 119710 0 119766 800
rect 120722 0 120778 800
rect 121642 0 121698 800
rect 122562 0 122618 800
rect 123482 0 123538 800
rect 124402 0 124458 800
rect 125414 0 125470 800
rect 126334 0 126390 800
rect 127254 0 127310 800
rect 128174 0 128230 800
rect 129094 0 129150 800
rect 130106 0 130162 800
rect 131026 0 131082 800
rect 131946 0 132002 800
rect 132866 0 132922 800
rect 133878 0 133934 800
rect 134798 0 134854 800
rect 135718 0 135774 800
rect 136638 0 136694 800
rect 137558 0 137614 800
rect 138570 0 138626 800
rect 139490 0 139546 800
rect 140410 0 140466 800
rect 141330 0 141386 800
rect 142250 0 142306 800
rect 143262 0 143318 800
rect 144182 0 144238 800
rect 145102 0 145158 800
rect 146022 0 146078 800
rect 146942 0 146998 800
rect 147954 0 148010 800
rect 148874 0 148930 800
rect 149794 0 149850 800
rect 150714 0 150770 800
rect 151726 0 151782 800
rect 152646 0 152702 800
rect 153566 0 153622 800
rect 154486 0 154542 800
rect 155406 0 155462 800
rect 156418 0 156474 800
rect 157338 0 157394 800
rect 158258 0 158314 800
rect 159178 0 159234 800
rect 160098 0 160154 800
rect 161110 0 161166 800
rect 162030 0 162086 800
rect 162950 0 163006 800
rect 163870 0 163926 800
<< obsm2 >>
rect 18 165665 330 165866
rect 498 165665 1158 165866
rect 1326 165665 2078 165866
rect 2246 165665 2998 165866
rect 3166 165665 3918 165866
rect 4086 165665 4838 165866
rect 5006 165665 5758 165866
rect 5926 165665 6678 165866
rect 6846 165665 7506 165866
rect 7674 165665 8426 165866
rect 8594 165665 9346 165866
rect 9514 165665 10266 165866
rect 10434 165665 11186 165866
rect 11354 165665 12106 165866
rect 12274 165665 13026 165866
rect 13194 165665 13946 165866
rect 14114 165665 14774 165866
rect 14942 165665 15694 165866
rect 15862 165665 16614 165866
rect 16782 165665 17534 165866
rect 17702 165665 18454 165866
rect 18622 165665 19374 165866
rect 19542 165665 20294 165866
rect 20462 165665 21214 165866
rect 21382 165665 22042 165866
rect 22210 165665 22962 165866
rect 23130 165665 23882 165866
rect 24050 165665 24802 165866
rect 24970 165665 25722 165866
rect 25890 165665 26642 165866
rect 26810 165665 27562 165866
rect 27730 165665 28482 165866
rect 28650 165665 29310 165866
rect 29478 165665 30230 165866
rect 30398 165665 31150 165866
rect 31318 165665 32070 165866
rect 32238 165665 32990 165866
rect 33158 165665 33910 165866
rect 34078 165665 34830 165866
rect 34998 165665 35750 165866
rect 35918 165665 36578 165866
rect 36746 165665 37498 165866
rect 37666 165665 38418 165866
rect 38586 165665 39338 165866
rect 39506 165665 40258 165866
rect 40426 165665 41178 165866
rect 41346 165665 42098 165866
rect 42266 165665 43018 165866
rect 43186 165665 43846 165866
rect 44014 165665 44766 165866
rect 44934 165665 45686 165866
rect 45854 165665 46606 165866
rect 46774 165665 47526 165866
rect 47694 165665 48446 165866
rect 48614 165665 49366 165866
rect 49534 165665 50286 165866
rect 50454 165665 51114 165866
rect 51282 165665 52034 165866
rect 52202 165665 52954 165866
rect 53122 165665 53874 165866
rect 54042 165665 54794 165866
rect 54962 165665 55714 165866
rect 55882 165665 56634 165866
rect 56802 165665 57462 165866
rect 57630 165665 58382 165866
rect 58550 165665 59302 165866
rect 59470 165665 60222 165866
rect 60390 165665 61142 165866
rect 61310 165665 62062 165866
rect 62230 165665 62982 165866
rect 63150 165665 63902 165866
rect 64070 165665 64730 165866
rect 64898 165665 65650 165866
rect 65818 165665 66570 165866
rect 66738 165665 67490 165866
rect 67658 165665 68410 165866
rect 68578 165665 69330 165866
rect 69498 165665 70250 165866
rect 70418 165665 71170 165866
rect 71338 165665 71998 165866
rect 72166 165665 72918 165866
rect 73086 165665 73838 165866
rect 74006 165665 74758 165866
rect 74926 165665 75678 165866
rect 75846 165665 76598 165866
rect 76766 165665 77518 165866
rect 77686 165665 78438 165866
rect 78606 165665 79266 165866
rect 79434 165665 80186 165866
rect 80354 165665 81106 165866
rect 81274 165665 82026 165866
rect 82194 165665 82946 165866
rect 83114 165665 83866 165866
rect 84034 165665 84786 165866
rect 84954 165665 85706 165866
rect 85874 165665 86534 165866
rect 86702 165665 87454 165866
rect 87622 165665 88374 165866
rect 88542 165665 89294 165866
rect 89462 165665 90214 165866
rect 90382 165665 91134 165866
rect 91302 165665 92054 165866
rect 92222 165665 92974 165866
rect 93142 165665 93802 165866
rect 93970 165665 94722 165866
rect 94890 165665 95642 165866
rect 95810 165665 96562 165866
rect 96730 165665 97482 165866
rect 97650 165665 98402 165866
rect 98570 165665 99322 165866
rect 99490 165665 100242 165866
rect 100410 165665 101070 165866
rect 101238 165665 101990 165866
rect 102158 165665 102910 165866
rect 103078 165665 103830 165866
rect 103998 165665 104750 165866
rect 104918 165665 105670 165866
rect 105838 165665 106590 165866
rect 106758 165665 107510 165866
rect 107678 165665 108338 165866
rect 108506 165665 109258 165866
rect 109426 165665 110178 165866
rect 110346 165665 111098 165866
rect 111266 165665 112018 165866
rect 112186 165665 112938 165866
rect 113106 165665 113858 165866
rect 114026 165665 114686 165866
rect 114854 165665 115606 165866
rect 115774 165665 116526 165866
rect 116694 165665 117446 165866
rect 117614 165665 118366 165866
rect 118534 165665 119286 165866
rect 119454 165665 120206 165866
rect 120374 165665 121126 165866
rect 121294 165665 121954 165866
rect 122122 165665 122874 165866
rect 123042 165665 123794 165866
rect 123962 165665 124714 165866
rect 124882 165665 125634 165866
rect 125802 165665 126554 165866
rect 126722 165665 127474 165866
rect 127642 165665 128394 165866
rect 128562 165665 129222 165866
rect 129390 165665 130142 165866
rect 130310 165665 131062 165866
rect 131230 165665 131982 165866
rect 132150 165665 132902 165866
rect 133070 165665 133822 165866
rect 133990 165665 134742 165866
rect 134910 165665 135662 165866
rect 135830 165665 136490 165866
rect 136658 165665 137410 165866
rect 137578 165665 138330 165866
rect 138498 165665 139250 165866
rect 139418 165665 140170 165866
rect 140338 165665 141090 165866
rect 141258 165665 142010 165866
rect 142178 165665 142930 165866
rect 143098 165665 143758 165866
rect 143926 165665 144678 165866
rect 144846 165665 145598 165866
rect 145766 165665 146518 165866
rect 146686 165665 147438 165866
rect 147606 165665 148358 165866
rect 148526 165665 149278 165866
rect 149446 165665 150198 165866
rect 150366 165665 151026 165866
rect 151194 165665 151946 165866
rect 152114 165665 152866 165866
rect 153034 165665 153786 165866
rect 153954 165665 154706 165866
rect 154874 165665 155626 165866
rect 155794 165665 156546 165866
rect 156714 165665 157466 165866
rect 157634 165665 158294 165866
rect 158462 165665 159214 165866
rect 159382 165665 160134 165866
rect 160302 165665 161054 165866
rect 161222 165665 161974 165866
rect 162142 165665 162894 165866
rect 163062 165665 163814 165866
rect 163982 165665 164372 165866
rect 18 856 164372 165665
rect 18 2 422 856
rect 590 2 1342 856
rect 1510 2 2262 856
rect 2430 2 3182 856
rect 3350 2 4102 856
rect 4270 2 5114 856
rect 5282 2 6034 856
rect 6202 2 6954 856
rect 7122 2 7874 856
rect 8042 2 8794 856
rect 8962 2 9806 856
rect 9974 2 10726 856
rect 10894 2 11646 856
rect 11814 2 12566 856
rect 12734 2 13486 856
rect 13654 2 14498 856
rect 14666 2 15418 856
rect 15586 2 16338 856
rect 16506 2 17258 856
rect 17426 2 18270 856
rect 18438 2 19190 856
rect 19358 2 20110 856
rect 20278 2 21030 856
rect 21198 2 21950 856
rect 22118 2 22962 856
rect 23130 2 23882 856
rect 24050 2 24802 856
rect 24970 2 25722 856
rect 25890 2 26642 856
rect 26810 2 27654 856
rect 27822 2 28574 856
rect 28742 2 29494 856
rect 29662 2 30414 856
rect 30582 2 31334 856
rect 31502 2 32346 856
rect 32514 2 33266 856
rect 33434 2 34186 856
rect 34354 2 35106 856
rect 35274 2 36118 856
rect 36286 2 37038 856
rect 37206 2 37958 856
rect 38126 2 38878 856
rect 39046 2 39798 856
rect 39966 2 40810 856
rect 40978 2 41730 856
rect 41898 2 42650 856
rect 42818 2 43570 856
rect 43738 2 44490 856
rect 44658 2 45502 856
rect 45670 2 46422 856
rect 46590 2 47342 856
rect 47510 2 48262 856
rect 48430 2 49182 856
rect 49350 2 50194 856
rect 50362 2 51114 856
rect 51282 2 52034 856
rect 52202 2 52954 856
rect 53122 2 53966 856
rect 54134 2 54886 856
rect 55054 2 55806 856
rect 55974 2 56726 856
rect 56894 2 57646 856
rect 57814 2 58658 856
rect 58826 2 59578 856
rect 59746 2 60498 856
rect 60666 2 61418 856
rect 61586 2 62338 856
rect 62506 2 63350 856
rect 63518 2 64270 856
rect 64438 2 65190 856
rect 65358 2 66110 856
rect 66278 2 67122 856
rect 67290 2 68042 856
rect 68210 2 68962 856
rect 69130 2 69882 856
rect 70050 2 70802 856
rect 70970 2 71814 856
rect 71982 2 72734 856
rect 72902 2 73654 856
rect 73822 2 74574 856
rect 74742 2 75494 856
rect 75662 2 76506 856
rect 76674 2 77426 856
rect 77594 2 78346 856
rect 78514 2 79266 856
rect 79434 2 80186 856
rect 80354 2 81198 856
rect 81366 2 82118 856
rect 82286 2 83038 856
rect 83206 2 83958 856
rect 84126 2 84970 856
rect 85138 2 85890 856
rect 86058 2 86810 856
rect 86978 2 87730 856
rect 87898 2 88650 856
rect 88818 2 89662 856
rect 89830 2 90582 856
rect 90750 2 91502 856
rect 91670 2 92422 856
rect 92590 2 93342 856
rect 93510 2 94354 856
rect 94522 2 95274 856
rect 95442 2 96194 856
rect 96362 2 97114 856
rect 97282 2 98034 856
rect 98202 2 99046 856
rect 99214 2 99966 856
rect 100134 2 100886 856
rect 101054 2 101806 856
rect 101974 2 102818 856
rect 102986 2 103738 856
rect 103906 2 104658 856
rect 104826 2 105578 856
rect 105746 2 106498 856
rect 106666 2 107510 856
rect 107678 2 108430 856
rect 108598 2 109350 856
rect 109518 2 110270 856
rect 110438 2 111190 856
rect 111358 2 112202 856
rect 112370 2 113122 856
rect 113290 2 114042 856
rect 114210 2 114962 856
rect 115130 2 115974 856
rect 116142 2 116894 856
rect 117062 2 117814 856
rect 117982 2 118734 856
rect 118902 2 119654 856
rect 119822 2 120666 856
rect 120834 2 121586 856
rect 121754 2 122506 856
rect 122674 2 123426 856
rect 123594 2 124346 856
rect 124514 2 125358 856
rect 125526 2 126278 856
rect 126446 2 127198 856
rect 127366 2 128118 856
rect 128286 2 129038 856
rect 129206 2 130050 856
rect 130218 2 130970 856
rect 131138 2 131890 856
rect 132058 2 132810 856
rect 132978 2 133822 856
rect 133990 2 134742 856
rect 134910 2 135662 856
rect 135830 2 136582 856
rect 136750 2 137502 856
rect 137670 2 138514 856
rect 138682 2 139434 856
rect 139602 2 140354 856
rect 140522 2 141274 856
rect 141442 2 142194 856
rect 142362 2 143206 856
rect 143374 2 144126 856
rect 144294 2 145046 856
rect 145214 2 145966 856
rect 146134 2 146886 856
rect 147054 2 147898 856
rect 148066 2 148818 856
rect 148986 2 149738 856
rect 149906 2 150658 856
rect 150826 2 151670 856
rect 151838 2 152590 856
rect 152758 2 153510 856
rect 153678 2 154430 856
rect 154598 2 155350 856
rect 155518 2 156362 856
rect 156530 2 157282 856
rect 157450 2 158202 856
rect 158370 2 159122 856
rect 159290 2 160042 856
rect 160210 2 161054 856
rect 161222 2 161974 856
rect 162142 2 162894 856
rect 163062 2 163814 856
rect 163982 2 164372 856
<< metal3 >>
rect 0 164976 800 165096
rect 163577 164704 164377 164824
rect 0 162120 800 162240
rect 163577 161440 164377 161560
rect 0 159264 800 159384
rect 163577 158040 164377 158160
rect 0 156544 800 156664
rect 163577 154776 164377 154896
rect 0 153688 800 153808
rect 163577 151376 164377 151496
rect 0 150832 800 150952
rect 0 147976 800 148096
rect 163577 148112 164377 148232
rect 0 145256 800 145376
rect 163577 144712 164377 144832
rect 0 142400 800 142520
rect 163577 141448 164377 141568
rect 0 139544 800 139664
rect 163577 138048 164377 138168
rect 0 136688 800 136808
rect 163577 134784 164377 134904
rect 0 133968 800 134088
rect 163577 131384 164377 131504
rect 0 131112 800 131232
rect 0 128256 800 128376
rect 163577 128120 164377 128240
rect 0 125400 800 125520
rect 163577 124720 164377 124840
rect 0 122680 800 122800
rect 163577 121456 164377 121576
rect 0 119824 800 119944
rect 163577 118056 164377 118176
rect 0 116968 800 117088
rect 163577 114792 164377 114912
rect 0 114112 800 114232
rect 0 111392 800 111512
rect 163577 111392 164377 111512
rect 0 108536 800 108656
rect 163577 108128 164377 108248
rect 0 105680 800 105800
rect 163577 104728 164377 104848
rect 0 102824 800 102944
rect 163577 101464 164377 101584
rect 0 100104 800 100224
rect 163577 98064 164377 98184
rect 0 97248 800 97368
rect 163577 94800 164377 94920
rect 0 94392 800 94512
rect 0 91536 800 91656
rect 163577 91400 164377 91520
rect 0 88816 800 88936
rect 163577 88136 164377 88256
rect 0 85960 800 86080
rect 163577 84872 164377 84992
rect 0 83104 800 83224
rect 163577 81472 164377 81592
rect 0 80248 800 80368
rect 163577 78208 164377 78328
rect 0 77528 800 77648
rect 0 74672 800 74792
rect 163577 74808 164377 74928
rect 0 71816 800 71936
rect 163577 71544 164377 71664
rect 0 68960 800 69080
rect 163577 68144 164377 68264
rect 0 66240 800 66360
rect 163577 64880 164377 65000
rect 0 63384 800 63504
rect 163577 61480 164377 61600
rect 0 60528 800 60648
rect 163577 58216 164377 58336
rect 0 57672 800 57792
rect 0 54952 800 55072
rect 163577 54816 164377 54936
rect 0 52096 800 52216
rect 163577 51552 164377 51672
rect 0 49240 800 49360
rect 163577 48152 164377 48272
rect 0 46384 800 46504
rect 163577 44888 164377 45008
rect 0 43664 800 43784
rect 163577 41488 164377 41608
rect 0 40808 800 40928
rect 163577 38224 164377 38344
rect 0 37952 800 38072
rect 0 35096 800 35216
rect 163577 34824 164377 34944
rect 0 32376 800 32496
rect 163577 31560 164377 31680
rect 0 29520 800 29640
rect 163577 28160 164377 28280
rect 0 26664 800 26784
rect 163577 24896 164377 25016
rect 0 23808 800 23928
rect 163577 21496 164377 21616
rect 0 21088 800 21208
rect 0 18232 800 18352
rect 163577 18232 164377 18352
rect 0 15376 800 15496
rect 163577 14832 164377 14952
rect 0 12520 800 12640
rect 163577 11568 164377 11688
rect 0 9800 800 9920
rect 163577 8168 164377 8288
rect 0 6944 800 7064
rect 163577 4904 164377 5024
rect 0 4088 800 4208
rect 163577 1640 164377 1760
rect 0 1368 800 1488
<< obsm3 >>
rect 880 164904 164299 165069
rect 880 164896 163497 164904
rect 13 164624 163497 164896
rect 13 162320 164299 164624
rect 880 162040 164299 162320
rect 13 161640 164299 162040
rect 13 161360 163497 161640
rect 13 159464 164299 161360
rect 880 159184 164299 159464
rect 13 158240 164299 159184
rect 13 157960 163497 158240
rect 13 156744 164299 157960
rect 880 156464 164299 156744
rect 13 154976 164299 156464
rect 13 154696 163497 154976
rect 13 153888 164299 154696
rect 880 153608 164299 153888
rect 13 151576 164299 153608
rect 13 151296 163497 151576
rect 13 151032 164299 151296
rect 880 150752 164299 151032
rect 13 148312 164299 150752
rect 13 148176 163497 148312
rect 880 148032 163497 148176
rect 880 147896 164299 148032
rect 13 145456 164299 147896
rect 880 145176 164299 145456
rect 13 144912 164299 145176
rect 13 144632 163497 144912
rect 13 142600 164299 144632
rect 880 142320 164299 142600
rect 13 141648 164299 142320
rect 13 141368 163497 141648
rect 13 139744 164299 141368
rect 880 139464 164299 139744
rect 13 138248 164299 139464
rect 13 137968 163497 138248
rect 13 136888 164299 137968
rect 880 136608 164299 136888
rect 13 134984 164299 136608
rect 13 134704 163497 134984
rect 13 134168 164299 134704
rect 880 133888 164299 134168
rect 13 131584 164299 133888
rect 13 131312 163497 131584
rect 880 131304 163497 131312
rect 880 131032 164299 131304
rect 13 128456 164299 131032
rect 880 128320 164299 128456
rect 880 128176 163497 128320
rect 13 128040 163497 128176
rect 13 125600 164299 128040
rect 880 125320 164299 125600
rect 13 124920 164299 125320
rect 13 124640 163497 124920
rect 13 122880 164299 124640
rect 880 122600 164299 122880
rect 13 121656 164299 122600
rect 13 121376 163497 121656
rect 13 120024 164299 121376
rect 880 119744 164299 120024
rect 13 118256 164299 119744
rect 13 117976 163497 118256
rect 13 117168 164299 117976
rect 880 116888 164299 117168
rect 13 114992 164299 116888
rect 13 114712 163497 114992
rect 13 114312 164299 114712
rect 880 114032 164299 114312
rect 13 111592 164299 114032
rect 880 111312 163497 111592
rect 13 108736 164299 111312
rect 880 108456 164299 108736
rect 13 108328 164299 108456
rect 13 108048 163497 108328
rect 13 105880 164299 108048
rect 880 105600 164299 105880
rect 13 104928 164299 105600
rect 13 104648 163497 104928
rect 13 103024 164299 104648
rect 880 102744 164299 103024
rect 13 101664 164299 102744
rect 13 101384 163497 101664
rect 13 100304 164299 101384
rect 880 100024 164299 100304
rect 13 98264 164299 100024
rect 13 97984 163497 98264
rect 13 97448 164299 97984
rect 880 97168 164299 97448
rect 13 95000 164299 97168
rect 13 94720 163497 95000
rect 13 94592 164299 94720
rect 880 94312 164299 94592
rect 13 91736 164299 94312
rect 880 91600 164299 91736
rect 880 91456 163497 91600
rect 13 91320 163497 91456
rect 13 89016 164299 91320
rect 880 88736 164299 89016
rect 13 88336 164299 88736
rect 13 88056 163497 88336
rect 13 86160 164299 88056
rect 880 85880 164299 86160
rect 13 85072 164299 85880
rect 13 84792 163497 85072
rect 13 83304 164299 84792
rect 880 83024 164299 83304
rect 13 81672 164299 83024
rect 13 81392 163497 81672
rect 13 80448 164299 81392
rect 880 80168 164299 80448
rect 13 78408 164299 80168
rect 13 78128 163497 78408
rect 13 77728 164299 78128
rect 880 77448 164299 77728
rect 13 75008 164299 77448
rect 13 74872 163497 75008
rect 880 74728 163497 74872
rect 880 74592 164299 74728
rect 13 72016 164299 74592
rect 880 71744 164299 72016
rect 880 71736 163497 71744
rect 13 71464 163497 71736
rect 13 69160 164299 71464
rect 880 68880 164299 69160
rect 13 68344 164299 68880
rect 13 68064 163497 68344
rect 13 66440 164299 68064
rect 880 66160 164299 66440
rect 13 65080 164299 66160
rect 13 64800 163497 65080
rect 13 63584 164299 64800
rect 880 63304 164299 63584
rect 13 61680 164299 63304
rect 13 61400 163497 61680
rect 13 60728 164299 61400
rect 880 60448 164299 60728
rect 13 58416 164299 60448
rect 13 58136 163497 58416
rect 13 57872 164299 58136
rect 880 57592 164299 57872
rect 13 55152 164299 57592
rect 880 55016 164299 55152
rect 880 54872 163497 55016
rect 13 54736 163497 54872
rect 13 52296 164299 54736
rect 880 52016 164299 52296
rect 13 51752 164299 52016
rect 13 51472 163497 51752
rect 13 49440 164299 51472
rect 880 49160 164299 49440
rect 13 48352 164299 49160
rect 13 48072 163497 48352
rect 13 46584 164299 48072
rect 880 46304 164299 46584
rect 13 45088 164299 46304
rect 13 44808 163497 45088
rect 13 43864 164299 44808
rect 880 43584 164299 43864
rect 13 41688 164299 43584
rect 13 41408 163497 41688
rect 13 41008 164299 41408
rect 880 40728 164299 41008
rect 13 38424 164299 40728
rect 13 38152 163497 38424
rect 880 38144 163497 38152
rect 880 37872 164299 38144
rect 13 35296 164299 37872
rect 880 35024 164299 35296
rect 880 35016 163497 35024
rect 13 34744 163497 35016
rect 13 32576 164299 34744
rect 880 32296 164299 32576
rect 13 31760 164299 32296
rect 13 31480 163497 31760
rect 13 29720 164299 31480
rect 880 29440 164299 29720
rect 13 28360 164299 29440
rect 13 28080 163497 28360
rect 13 26864 164299 28080
rect 880 26584 164299 26864
rect 13 25096 164299 26584
rect 13 24816 163497 25096
rect 13 24008 164299 24816
rect 880 23728 164299 24008
rect 13 21696 164299 23728
rect 13 21416 163497 21696
rect 13 21288 164299 21416
rect 880 21008 164299 21288
rect 13 18432 164299 21008
rect 880 18152 163497 18432
rect 13 15576 164299 18152
rect 880 15296 164299 15576
rect 13 15032 164299 15296
rect 13 14752 163497 15032
rect 13 12720 164299 14752
rect 880 12440 164299 12720
rect 13 11768 164299 12440
rect 13 11488 163497 11768
rect 13 10000 164299 11488
rect 880 9720 164299 10000
rect 13 8368 164299 9720
rect 13 8088 163497 8368
rect 13 7144 164299 8088
rect 880 6864 164299 7144
rect 13 5104 164299 6864
rect 13 4824 163497 5104
rect 13 4288 164299 4824
rect 880 4008 164299 4288
rect 13 1840 164299 4008
rect 13 1568 163497 1840
rect 880 1560 163497 1568
rect 880 1288 164299 1560
rect 13 35 164299 1288
<< metal4 >>
rect 4208 2128 4528 164336
rect 19568 2128 19888 164336
rect 34928 2128 35248 164336
rect 50288 2128 50608 164336
rect 65648 2128 65968 164336
rect 81008 2128 81328 164336
rect 96368 2128 96688 164336
rect 111728 2128 112048 164336
rect 127088 2128 127408 164336
rect 142448 2128 142768 164336
rect 157808 2128 158128 164336
<< obsm4 >>
rect 427 2048 4128 163981
rect 4608 2048 19488 163981
rect 19968 2048 34848 163981
rect 35328 2048 50208 163981
rect 50688 2048 65568 163981
rect 66048 2048 80928 163981
rect 81408 2048 96288 163981
rect 96768 2048 111648 163981
rect 112128 2048 127008 163981
rect 127488 2048 142368 163981
rect 142848 2048 153213 163981
rect 427 987 153213 2048
<< labels >>
rlabel metal2 s 104806 165721 104862 166521 6 i_dout0[0]
port 1 nsew signal input
rlabel metal2 s 131118 165721 131174 166521 6 i_dout0[10]
port 2 nsew signal input
rlabel metal2 s 132958 165721 133014 166521 6 i_dout0[11]
port 3 nsew signal input
rlabel metal2 s 134798 165721 134854 166521 6 i_dout0[12]
port 4 nsew signal input
rlabel metal2 s 136546 165721 136602 166521 6 i_dout0[13]
port 5 nsew signal input
rlabel metal2 s 143262 0 143318 800 6 i_dout0[14]
port 6 nsew signal input
rlabel metal3 s 163577 111392 164377 111512 6 i_dout0[15]
port 7 nsew signal input
rlabel metal2 s 146942 0 146998 800 6 i_dout0[16]
port 8 nsew signal input
rlabel metal2 s 142986 165721 143042 166521 6 i_dout0[17]
port 9 nsew signal input
rlabel metal3 s 163577 121456 164377 121576 6 i_dout0[18]
port 10 nsew signal input
rlabel metal2 s 147494 165721 147550 166521 6 i_dout0[19]
port 11 nsew signal input
rlabel metal2 s 105634 0 105690 800 6 i_dout0[1]
port 12 nsew signal input
rlabel metal3 s 0 88816 800 88936 6 i_dout0[20]
port 13 nsew signal input
rlabel metal2 s 154486 0 154542 800 6 i_dout0[21]
port 14 nsew signal input
rlabel metal2 s 151082 165721 151138 166521 6 i_dout0[22]
port 15 nsew signal input
rlabel metal2 s 158258 0 158314 800 6 i_dout0[23]
port 16 nsew signal input
rlabel metal3 s 163577 138048 164377 138168 6 i_dout0[24]
port 17 nsew signal input
rlabel metal2 s 154762 165721 154818 166521 6 i_dout0[25]
port 18 nsew signal input
rlabel metal3 s 0 119824 800 119944 6 i_dout0[26]
port 19 nsew signal input
rlabel metal2 s 157522 165721 157578 166521 6 i_dout0[27]
port 20 nsew signal input
rlabel metal3 s 163577 161440 164377 161560 6 i_dout0[28]
port 21 nsew signal input
rlabel metal2 s 163870 0 163926 800 6 i_dout0[29]
port 22 nsew signal input
rlabel metal2 s 109406 0 109462 800 6 i_dout0[2]
port 23 nsew signal input
rlabel metal3 s 0 150832 800 150952 6 i_dout0[30]
port 24 nsew signal input
rlabel metal3 s 0 156544 800 156664 6 i_dout0[31]
port 25 nsew signal input
rlabel metal2 s 116030 0 116086 800 6 i_dout0[3]
port 26 nsew signal input
rlabel metal2 s 116582 165721 116638 166521 6 i_dout0[4]
port 27 nsew signal input
rlabel metal2 s 119342 165721 119398 166521 6 i_dout0[5]
port 28 nsew signal input
rlabel metal2 s 124402 0 124458 800 6 i_dout0[6]
port 29 nsew signal input
rlabel metal3 s 163577 68144 164377 68264 6 i_dout0[7]
port 30 nsew signal input
rlabel metal2 s 128174 0 128230 800 6 i_dout0[8]
port 31 nsew signal input
rlabel metal3 s 0 57672 800 57792 6 i_dout0[9]
port 32 nsew signal input
rlabel metal3 s 163577 8168 164377 8288 6 i_dout0_1[0]
port 33 nsew signal input
rlabel metal2 s 130198 165721 130254 166521 6 i_dout0_1[10]
port 34 nsew signal input
rlabel metal2 s 133878 0 133934 800 6 i_dout0_1[11]
port 35 nsew signal input
rlabel metal2 s 137558 0 137614 800 6 i_dout0_1[12]
port 36 nsew signal input
rlabel metal2 s 140410 0 140466 800 6 i_dout0_1[13]
port 37 nsew signal input
rlabel metal3 s 163577 104728 164377 104848 6 i_dout0_1[14]
port 38 nsew signal input
rlabel metal3 s 163577 108128 164377 108248 6 i_dout0_1[15]
port 39 nsew signal input
rlabel metal3 s 0 71816 800 71936 6 i_dout0_1[16]
port 40 nsew signal input
rlabel metal2 s 147954 0 148010 800 6 i_dout0_1[17]
port 41 nsew signal input
rlabel metal3 s 0 77528 800 77648 6 i_dout0_1[18]
port 42 nsew signal input
rlabel metal2 s 146574 165721 146630 166521 6 i_dout0_1[19]
port 43 nsew signal input
rlabel metal3 s 163577 21496 164377 21616 6 i_dout0_1[1]
port 44 nsew signal input
rlabel metal3 s 163577 128120 164377 128240 6 i_dout0_1[20]
port 45 nsew signal input
rlabel metal2 s 153566 0 153622 800 6 i_dout0_1[21]
port 46 nsew signal input
rlabel metal2 s 150254 165721 150310 166521 6 i_dout0_1[22]
port 47 nsew signal input
rlabel metal2 s 152922 165721 152978 166521 6 i_dout0_1[23]
port 48 nsew signal input
rlabel metal3 s 0 108536 800 108656 6 i_dout0_1[24]
port 49 nsew signal input
rlabel metal3 s 0 114112 800 114232 6 i_dout0_1[25]
port 50 nsew signal input
rlabel metal2 s 161110 0 161166 800 6 i_dout0_1[26]
port 51 nsew signal input
rlabel metal3 s 0 128256 800 128376 6 i_dout0_1[27]
port 52 nsew signal input
rlabel metal3 s 0 133968 800 134088 6 i_dout0_1[28]
port 53 nsew signal input
rlabel metal3 s 0 139544 800 139664 6 i_dout0_1[29]
port 54 nsew signal input
rlabel metal3 s 0 15376 800 15496 6 i_dout0_1[2]
port 55 nsew signal input
rlabel metal2 s 161110 165721 161166 166521 6 i_dout0_1[30]
port 56 nsew signal input
rlabel metal2 s 163870 165721 163926 166521 6 i_dout0_1[31]
port 57 nsew signal input
rlabel metal3 s 163577 34824 164377 34944 6 i_dout0_1[3]
port 58 nsew signal input
rlabel metal3 s 0 35096 800 35216 6 i_dout0_1[4]
port 59 nsew signal input
rlabel metal2 s 118422 165721 118478 166521 6 i_dout0_1[5]
port 60 nsew signal input
rlabel metal3 s 163577 54816 164377 54936 6 i_dout0_1[6]
port 61 nsew signal input
rlabel metal3 s 0 49240 800 49360 6 i_dout0_1[7]
port 62 nsew signal input
rlabel metal3 s 0 54952 800 55072 6 i_dout0_1[8]
port 63 nsew signal input
rlabel metal2 s 129278 165721 129334 166521 6 i_dout0_1[9]
port 64 nsew signal input
rlabel metal2 s 103794 0 103850 800 6 i_dout1[0]
port 65 nsew signal input
rlabel metal3 s 0 60528 800 60648 6 i_dout1[10]
port 66 nsew signal input
rlabel metal2 s 134798 0 134854 800 6 i_dout1[11]
port 67 nsew signal input
rlabel metal2 s 135718 165721 135774 166521 6 i_dout1[12]
port 68 nsew signal input
rlabel metal3 s 163577 101464 164377 101584 6 i_dout1[13]
port 69 nsew signal input
rlabel metal2 s 137466 165721 137522 166521 6 i_dout1[14]
port 70 nsew signal input
rlabel metal2 s 145102 0 145158 800 6 i_dout1[15]
port 71 nsew signal input
rlabel metal2 s 141146 165721 141202 166521 6 i_dout1[16]
port 72 nsew signal input
rlabel metal2 s 143814 165721 143870 166521 6 i_dout1[17]
port 73 nsew signal input
rlabel metal3 s 0 80248 800 80368 6 i_dout1[18]
port 74 nsew signal input
rlabel metal2 s 148414 165721 148470 166521 6 i_dout1[19]
port 75 nsew signal input
rlabel metal2 s 108394 165721 108450 166521 6 i_dout1[1]
port 76 nsew signal input
rlabel metal2 s 151726 0 151782 800 6 i_dout1[20]
port 77 nsew signal input
rlabel metal2 s 155406 0 155462 800 6 i_dout1[21]
port 78 nsew signal input
rlabel metal2 s 152002 165721 152058 166521 6 i_dout1[22]
port 79 nsew signal input
rlabel metal3 s 0 100104 800 100224 6 i_dout1[23]
port 80 nsew signal input
rlabel metal2 s 153842 165721 153898 166521 6 i_dout1[24]
port 81 nsew signal input
rlabel metal2 s 160098 0 160154 800 6 i_dout1[25]
port 82 nsew signal input
rlabel metal2 s 156602 165721 156658 166521 6 i_dout1[26]
port 83 nsew signal input
rlabel metal2 s 158350 165721 158406 166521 6 i_dout1[27]
port 84 nsew signal input
rlabel metal2 s 162030 0 162086 800 6 i_dout1[28]
port 85 nsew signal input
rlabel metal2 s 160190 165721 160246 166521 6 i_dout1[29]
port 86 nsew signal input
rlabel metal2 s 110326 0 110382 800 6 i_dout1[2]
port 87 nsew signal input
rlabel metal2 s 162030 165721 162086 166521 6 i_dout1[30]
port 88 nsew signal input
rlabel metal3 s 0 159264 800 159384 6 i_dout1[31]
port 89 nsew signal input
rlabel metal2 s 116950 0 117006 800 6 i_dout1[3]
port 90 nsew signal input
rlabel metal2 s 118790 0 118846 800 6 i_dout1[4]
port 91 nsew signal input
rlabel metal2 s 121642 0 121698 800 6 i_dout1[5]
port 92 nsew signal input
rlabel metal3 s 163577 61480 164377 61600 6 i_dout1[6]
port 93 nsew signal input
rlabel metal3 s 0 52096 800 52216 6 i_dout1[7]
port 94 nsew signal input
rlabel metal3 s 163577 81472 164377 81592 6 i_dout1[8]
port 95 nsew signal input
rlabel metal3 s 163577 91400 164377 91520 6 i_dout1[9]
port 96 nsew signal input
rlabel metal2 s 105726 165721 105782 166521 6 i_dout1_1[0]
port 97 nsew signal input
rlabel metal2 s 132866 0 132922 800 6 i_dout1_1[10]
port 98 nsew signal input
rlabel metal3 s 163577 98064 164377 98184 6 i_dout1_1[11]
port 99 nsew signal input
rlabel metal2 s 133878 165721 133934 166521 6 i_dout1_1[12]
port 100 nsew signal input
rlabel metal2 s 141330 0 141386 800 6 i_dout1_1[13]
port 101 nsew signal input
rlabel metal3 s 0 66240 800 66360 6 i_dout1_1[14]
port 102 nsew signal input
rlabel metal2 s 144182 0 144238 800 6 i_dout1_1[15]
port 103 nsew signal input
rlabel metal2 s 146022 0 146078 800 6 i_dout1_1[16]
port 104 nsew signal input
rlabel metal2 s 142066 165721 142122 166521 6 i_dout1_1[17]
port 105 nsew signal input
rlabel metal2 s 145654 165721 145710 166521 6 i_dout1_1[18]
port 106 nsew signal input
rlabel metal3 s 163577 124720 164377 124840 6 i_dout1_1[19]
port 107 nsew signal input
rlabel metal3 s 0 12520 800 12640 6 i_dout1_1[1]
port 108 nsew signal input
rlabel metal3 s 0 85960 800 86080 6 i_dout1_1[20]
port 109 nsew signal input
rlabel metal2 s 149334 165721 149390 166521 6 i_dout1_1[21]
port 110 nsew signal input
rlabel metal3 s 163577 131384 164377 131504 6 i_dout1_1[22]
port 111 nsew signal input
rlabel metal3 s 0 97248 800 97368 6 i_dout1_1[23]
port 112 nsew signal input
rlabel metal2 s 159178 0 159234 800 6 i_dout1_1[24]
port 113 nsew signal input
rlabel metal3 s 163577 144712 164377 144832 6 i_dout1_1[25]
port 114 nsew signal input
rlabel metal2 s 155682 165721 155738 166521 6 i_dout1_1[26]
port 115 nsew signal input
rlabel metal3 s 0 131112 800 131232 6 i_dout1_1[27]
port 116 nsew signal input
rlabel metal3 s 163577 158040 164377 158160 6 i_dout1_1[28]
port 117 nsew signal input
rlabel metal2 s 159270 165721 159326 166521 6 i_dout1_1[29]
port 118 nsew signal input
rlabel metal2 s 108486 0 108542 800 6 i_dout1_1[2]
port 119 nsew signal input
rlabel metal3 s 0 147976 800 148096 6 i_dout1_1[30]
port 120 nsew signal input
rlabel metal3 s 0 153688 800 153808 6 i_dout1_1[31]
port 121 nsew signal input
rlabel metal2 s 112994 165721 113050 166521 6 i_dout1_1[3]
port 122 nsew signal input
rlabel metal2 s 115662 165721 115718 166521 6 i_dout1_1[4]
port 123 nsew signal input
rlabel metal3 s 163577 48152 164377 48272 6 i_dout1_1[5]
port 124 nsew signal input
rlabel metal3 s 163577 58216 164377 58336 6 i_dout1_1[6]
port 125 nsew signal input
rlabel metal2 s 123850 165721 123906 166521 6 i_dout1_1[7]
port 126 nsew signal input
rlabel metal2 s 127254 0 127310 800 6 i_dout1_1[8]
port 127 nsew signal input
rlabel metal2 s 130106 0 130162 800 6 i_dout1_1[9]
port 128 nsew signal input
rlabel metal2 s 386 165721 442 166521 6 io_in[0]
port 129 nsew signal input
rlabel metal2 s 27618 165721 27674 166521 6 io_in[10]
port 130 nsew signal input
rlabel metal2 s 30286 165721 30342 166521 6 io_in[11]
port 131 nsew signal input
rlabel metal2 s 33046 165721 33102 166521 6 io_in[12]
port 132 nsew signal input
rlabel metal2 s 35806 165721 35862 166521 6 io_in[13]
port 133 nsew signal input
rlabel metal2 s 38474 165721 38530 166521 6 io_in[14]
port 134 nsew signal input
rlabel metal2 s 41234 165721 41290 166521 6 io_in[15]
port 135 nsew signal input
rlabel metal2 s 43902 165721 43958 166521 6 io_in[16]
port 136 nsew signal input
rlabel metal2 s 46662 165721 46718 166521 6 io_in[17]
port 137 nsew signal input
rlabel metal2 s 49422 165721 49478 166521 6 io_in[18]
port 138 nsew signal input
rlabel metal2 s 52090 165721 52146 166521 6 io_in[19]
port 139 nsew signal input
rlabel metal2 s 3054 165721 3110 166521 6 io_in[1]
port 140 nsew signal input
rlabel metal2 s 54850 165721 54906 166521 6 io_in[20]
port 141 nsew signal input
rlabel metal2 s 57518 165721 57574 166521 6 io_in[21]
port 142 nsew signal input
rlabel metal2 s 60278 165721 60334 166521 6 io_in[22]
port 143 nsew signal input
rlabel metal2 s 63038 165721 63094 166521 6 io_in[23]
port 144 nsew signal input
rlabel metal2 s 65706 165721 65762 166521 6 io_in[24]
port 145 nsew signal input
rlabel metal2 s 68466 165721 68522 166521 6 io_in[25]
port 146 nsew signal input
rlabel metal2 s 71226 165721 71282 166521 6 io_in[26]
port 147 nsew signal input
rlabel metal2 s 73894 165721 73950 166521 6 io_in[27]
port 148 nsew signal input
rlabel metal2 s 76654 165721 76710 166521 6 io_in[28]
port 149 nsew signal input
rlabel metal2 s 79322 165721 79378 166521 6 io_in[29]
port 150 nsew signal input
rlabel metal2 s 5814 165721 5870 166521 6 io_in[2]
port 151 nsew signal input
rlabel metal2 s 82082 165721 82138 166521 6 io_in[30]
port 152 nsew signal input
rlabel metal2 s 84842 165721 84898 166521 6 io_in[31]
port 153 nsew signal input
rlabel metal2 s 87510 165721 87566 166521 6 io_in[32]
port 154 nsew signal input
rlabel metal2 s 90270 165721 90326 166521 6 io_in[33]
port 155 nsew signal input
rlabel metal2 s 93030 165721 93086 166521 6 io_in[34]
port 156 nsew signal input
rlabel metal2 s 95698 165721 95754 166521 6 io_in[35]
port 157 nsew signal input
rlabel metal2 s 98458 165721 98514 166521 6 io_in[36]
port 158 nsew signal input
rlabel metal2 s 101126 165721 101182 166521 6 io_in[37]
port 159 nsew signal input
rlabel metal2 s 8482 165721 8538 166521 6 io_in[3]
port 160 nsew signal input
rlabel metal2 s 11242 165721 11298 166521 6 io_in[4]
port 161 nsew signal input
rlabel metal2 s 14002 165721 14058 166521 6 io_in[5]
port 162 nsew signal input
rlabel metal2 s 16670 165721 16726 166521 6 io_in[6]
port 163 nsew signal input
rlabel metal2 s 19430 165721 19486 166521 6 io_in[7]
port 164 nsew signal input
rlabel metal2 s 22098 165721 22154 166521 6 io_in[8]
port 165 nsew signal input
rlabel metal2 s 24858 165721 24914 166521 6 io_in[9]
port 166 nsew signal input
rlabel metal2 s 1214 165721 1270 166521 6 io_oeb[0]
port 167 nsew signal output
rlabel metal2 s 28538 165721 28594 166521 6 io_oeb[10]
port 168 nsew signal output
rlabel metal2 s 31206 165721 31262 166521 6 io_oeb[11]
port 169 nsew signal output
rlabel metal2 s 33966 165721 34022 166521 6 io_oeb[12]
port 170 nsew signal output
rlabel metal2 s 36634 165721 36690 166521 6 io_oeb[13]
port 171 nsew signal output
rlabel metal2 s 39394 165721 39450 166521 6 io_oeb[14]
port 172 nsew signal output
rlabel metal2 s 42154 165721 42210 166521 6 io_oeb[15]
port 173 nsew signal output
rlabel metal2 s 44822 165721 44878 166521 6 io_oeb[16]
port 174 nsew signal output
rlabel metal2 s 47582 165721 47638 166521 6 io_oeb[17]
port 175 nsew signal output
rlabel metal2 s 50342 165721 50398 166521 6 io_oeb[18]
port 176 nsew signal output
rlabel metal2 s 53010 165721 53066 166521 6 io_oeb[19]
port 177 nsew signal output
rlabel metal2 s 3974 165721 4030 166521 6 io_oeb[1]
port 178 nsew signal output
rlabel metal2 s 55770 165721 55826 166521 6 io_oeb[20]
port 179 nsew signal output
rlabel metal2 s 58438 165721 58494 166521 6 io_oeb[21]
port 180 nsew signal output
rlabel metal2 s 61198 165721 61254 166521 6 io_oeb[22]
port 181 nsew signal output
rlabel metal2 s 63958 165721 64014 166521 6 io_oeb[23]
port 182 nsew signal output
rlabel metal2 s 66626 165721 66682 166521 6 io_oeb[24]
port 183 nsew signal output
rlabel metal2 s 69386 165721 69442 166521 6 io_oeb[25]
port 184 nsew signal output
rlabel metal2 s 72054 165721 72110 166521 6 io_oeb[26]
port 185 nsew signal output
rlabel metal2 s 74814 165721 74870 166521 6 io_oeb[27]
port 186 nsew signal output
rlabel metal2 s 77574 165721 77630 166521 6 io_oeb[28]
port 187 nsew signal output
rlabel metal2 s 80242 165721 80298 166521 6 io_oeb[29]
port 188 nsew signal output
rlabel metal2 s 6734 165721 6790 166521 6 io_oeb[2]
port 189 nsew signal output
rlabel metal2 s 83002 165721 83058 166521 6 io_oeb[30]
port 190 nsew signal output
rlabel metal2 s 85762 165721 85818 166521 6 io_oeb[31]
port 191 nsew signal output
rlabel metal2 s 88430 165721 88486 166521 6 io_oeb[32]
port 192 nsew signal output
rlabel metal2 s 91190 165721 91246 166521 6 io_oeb[33]
port 193 nsew signal output
rlabel metal2 s 93858 165721 93914 166521 6 io_oeb[34]
port 194 nsew signal output
rlabel metal2 s 96618 165721 96674 166521 6 io_oeb[35]
port 195 nsew signal output
rlabel metal2 s 99378 165721 99434 166521 6 io_oeb[36]
port 196 nsew signal output
rlabel metal2 s 102046 165721 102102 166521 6 io_oeb[37]
port 197 nsew signal output
rlabel metal2 s 9402 165721 9458 166521 6 io_oeb[3]
port 198 nsew signal output
rlabel metal2 s 12162 165721 12218 166521 6 io_oeb[4]
port 199 nsew signal output
rlabel metal2 s 14830 165721 14886 166521 6 io_oeb[5]
port 200 nsew signal output
rlabel metal2 s 17590 165721 17646 166521 6 io_oeb[6]
port 201 nsew signal output
rlabel metal2 s 20350 165721 20406 166521 6 io_oeb[7]
port 202 nsew signal output
rlabel metal2 s 23018 165721 23074 166521 6 io_oeb[8]
port 203 nsew signal output
rlabel metal2 s 25778 165721 25834 166521 6 io_oeb[9]
port 204 nsew signal output
rlabel metal2 s 2134 165721 2190 166521 6 io_out[0]
port 205 nsew signal output
rlabel metal2 s 29366 165721 29422 166521 6 io_out[10]
port 206 nsew signal output
rlabel metal2 s 32126 165721 32182 166521 6 io_out[11]
port 207 nsew signal output
rlabel metal2 s 34886 165721 34942 166521 6 io_out[12]
port 208 nsew signal output
rlabel metal2 s 37554 165721 37610 166521 6 io_out[13]
port 209 nsew signal output
rlabel metal2 s 40314 165721 40370 166521 6 io_out[14]
port 210 nsew signal output
rlabel metal2 s 43074 165721 43130 166521 6 io_out[15]
port 211 nsew signal output
rlabel metal2 s 45742 165721 45798 166521 6 io_out[16]
port 212 nsew signal output
rlabel metal2 s 48502 165721 48558 166521 6 io_out[17]
port 213 nsew signal output
rlabel metal2 s 51170 165721 51226 166521 6 io_out[18]
port 214 nsew signal output
rlabel metal2 s 53930 165721 53986 166521 6 io_out[19]
port 215 nsew signal output
rlabel metal2 s 4894 165721 4950 166521 6 io_out[1]
port 216 nsew signal output
rlabel metal2 s 56690 165721 56746 166521 6 io_out[20]
port 217 nsew signal output
rlabel metal2 s 59358 165721 59414 166521 6 io_out[21]
port 218 nsew signal output
rlabel metal2 s 62118 165721 62174 166521 6 io_out[22]
port 219 nsew signal output
rlabel metal2 s 64786 165721 64842 166521 6 io_out[23]
port 220 nsew signal output
rlabel metal2 s 67546 165721 67602 166521 6 io_out[24]
port 221 nsew signal output
rlabel metal2 s 70306 165721 70362 166521 6 io_out[25]
port 222 nsew signal output
rlabel metal2 s 72974 165721 73030 166521 6 io_out[26]
port 223 nsew signal output
rlabel metal2 s 75734 165721 75790 166521 6 io_out[27]
port 224 nsew signal output
rlabel metal2 s 78494 165721 78550 166521 6 io_out[28]
port 225 nsew signal output
rlabel metal2 s 81162 165721 81218 166521 6 io_out[29]
port 226 nsew signal output
rlabel metal2 s 7562 165721 7618 166521 6 io_out[2]
port 227 nsew signal output
rlabel metal2 s 83922 165721 83978 166521 6 io_out[30]
port 228 nsew signal output
rlabel metal2 s 86590 165721 86646 166521 6 io_out[31]
port 229 nsew signal output
rlabel metal2 s 89350 165721 89406 166521 6 io_out[32]
port 230 nsew signal output
rlabel metal2 s 92110 165721 92166 166521 6 io_out[33]
port 231 nsew signal output
rlabel metal2 s 94778 165721 94834 166521 6 io_out[34]
port 232 nsew signal output
rlabel metal2 s 97538 165721 97594 166521 6 io_out[35]
port 233 nsew signal output
rlabel metal2 s 100298 165721 100354 166521 6 io_out[36]
port 234 nsew signal output
rlabel metal2 s 102966 165721 103022 166521 6 io_out[37]
port 235 nsew signal output
rlabel metal2 s 10322 165721 10378 166521 6 io_out[3]
port 236 nsew signal output
rlabel metal2 s 13082 165721 13138 166521 6 io_out[4]
port 237 nsew signal output
rlabel metal2 s 15750 165721 15806 166521 6 io_out[5]
port 238 nsew signal output
rlabel metal2 s 18510 165721 18566 166521 6 io_out[6]
port 239 nsew signal output
rlabel metal2 s 21270 165721 21326 166521 6 io_out[7]
port 240 nsew signal output
rlabel metal2 s 23938 165721 23994 166521 6 io_out[8]
port 241 nsew signal output
rlabel metal2 s 26698 165721 26754 166521 6 io_out[9]
port 242 nsew signal output
rlabel metal2 s 100022 0 100078 800 6 irq[0]
port 243 nsew signal output
rlabel metal2 s 100942 0 100998 800 6 irq[1]
port 244 nsew signal output
rlabel metal2 s 101862 0 101918 800 6 irq[2]
port 245 nsew signal output
rlabel metal3 s 163577 14832 164377 14952 6 o_addr1[0]
port 246 nsew signal output
rlabel metal2 s 109314 165721 109370 166521 6 o_addr1[1]
port 247 nsew signal output
rlabel metal2 s 111246 0 111302 800 6 o_addr1[2]
port 248 nsew signal output
rlabel metal2 s 113914 165721 113970 166521 6 o_addr1[3]
port 249 nsew signal output
rlabel metal2 s 119710 0 119766 800 6 o_addr1[4]
port 250 nsew signal output
rlabel metal2 s 122562 0 122618 800 6 o_addr1[5]
port 251 nsew signal output
rlabel metal2 s 122010 165721 122066 166521 6 o_addr1[6]
port 252 nsew signal output
rlabel metal3 s 163577 71544 164377 71664 6 o_addr1[7]
port 253 nsew signal output
rlabel metal3 s 163577 84872 164377 84992 6 o_addr1[8]
port 254 nsew signal output
rlabel metal3 s 163577 11568 164377 11688 6 o_addr1_1[0]
port 255 nsew signal output
rlabel metal3 s 163577 24896 164377 25016 6 o_addr1_1[1]
port 256 nsew signal output
rlabel metal3 s 0 18232 800 18352 6 o_addr1_1[2]
port 257 nsew signal output
rlabel metal3 s 163577 38224 164377 38344 6 o_addr1_1[3]
port 258 nsew signal output
rlabel metal3 s 163577 41488 164377 41608 6 o_addr1_1[4]
port 259 nsew signal output
rlabel metal3 s 163577 51552 164377 51672 6 o_addr1_1[5]
port 260 nsew signal output
rlabel metal2 s 125414 0 125470 800 6 o_addr1_1[6]
port 261 nsew signal output
rlabel metal2 s 126334 0 126390 800 6 o_addr1_1[7]
port 262 nsew signal output
rlabel metal2 s 129094 0 129150 800 6 o_addr1_1[8]
port 263 nsew signal output
rlabel metal3 s 163577 1640 164377 1760 6 o_csb0
port 264 nsew signal output
rlabel metal3 s 0 1368 800 1488 6 o_csb0_1
port 265 nsew signal output
rlabel metal3 s 163577 4904 164377 5024 6 o_csb1
port 266 nsew signal output
rlabel metal2 s 103886 165721 103942 166521 6 o_csb1_1
port 267 nsew signal output
rlabel metal2 s 106646 165721 106702 166521 6 o_din0[0]
port 268 nsew signal output
rlabel metal2 s 132038 165721 132094 166521 6 o_din0[10]
port 269 nsew signal output
rlabel metal2 s 136638 0 136694 800 6 o_din0[11]
port 270 nsew signal output
rlabel metal2 s 139490 0 139546 800 6 o_din0[12]
port 271 nsew signal output
rlabel metal3 s 0 63384 800 63504 6 o_din0[13]
port 272 nsew signal output
rlabel metal3 s 0 68960 800 69080 6 o_din0[14]
port 273 nsew signal output
rlabel metal2 s 140226 165721 140282 166521 6 o_din0[15]
port 274 nsew signal output
rlabel metal3 s 0 74672 800 74792 6 o_din0[16]
port 275 nsew signal output
rlabel metal3 s 163577 118056 164377 118176 6 o_din0[17]
port 276 nsew signal output
rlabel metal2 s 149794 0 149850 800 6 o_din0[18]
port 277 nsew signal output
rlabel metal2 s 150714 0 150770 800 6 o_din0[19]
port 278 nsew signal output
rlabel metal2 s 110234 165721 110290 166521 6 o_din0[1]
port 279 nsew signal output
rlabel metal3 s 0 91536 800 91656 6 o_din0[20]
port 280 nsew signal output
rlabel metal3 s 0 94392 800 94512 6 o_din0[21]
port 281 nsew signal output
rlabel metal2 s 157338 0 157394 800 6 o_din0[22]
port 282 nsew signal output
rlabel metal3 s 0 105680 800 105800 6 o_din0[23]
port 283 nsew signal output
rlabel metal3 s 163577 141448 164377 141568 6 o_din0[24]
port 284 nsew signal output
rlabel metal3 s 163577 148112 164377 148232 6 o_din0[25]
port 285 nsew signal output
rlabel metal3 s 0 125400 800 125520 6 o_din0[26]
port 286 nsew signal output
rlabel metal3 s 163577 154776 164377 154896 6 o_din0[27]
port 287 nsew signal output
rlabel metal3 s 0 136688 800 136808 6 o_din0[28]
port 288 nsew signal output
rlabel metal3 s 0 145256 800 145376 6 o_din0[29]
port 289 nsew signal output
rlabel metal2 s 113178 0 113234 800 6 o_din0[2]
port 290 nsew signal output
rlabel metal3 s 163577 164704 164377 164824 6 o_din0[30]
port 291 nsew signal output
rlabel metal3 s 0 164976 800 165096 6 o_din0[31]
port 292 nsew signal output
rlabel metal2 s 114742 165721 114798 166521 6 o_din0[3]
port 293 nsew signal output
rlabel metal2 s 120722 0 120778 800 6 o_din0[4]
port 294 nsew signal output
rlabel metal2 s 121182 165721 121238 166521 6 o_din0[5]
port 295 nsew signal output
rlabel metal3 s 0 43664 800 43784 6 o_din0[6]
port 296 nsew signal output
rlabel metal2 s 125690 165721 125746 166521 6 o_din0[7]
port 297 nsew signal output
rlabel metal2 s 127530 165721 127586 166521 6 o_din0[8]
port 298 nsew signal output
rlabel metal2 s 131946 0 132002 800 6 o_din0[9]
port 299 nsew signal output
rlabel metal3 s 0 6944 800 7064 6 o_din0_1[0]
port 300 nsew signal output
rlabel metal3 s 163577 94800 164377 94920 6 o_din0_1[10]
port 301 nsew signal output
rlabel metal2 s 135718 0 135774 800 6 o_din0_1[11]
port 302 nsew signal output
rlabel metal2 s 138570 0 138626 800 6 o_din0_1[12]
port 303 nsew signal output
rlabel metal2 s 142250 0 142306 800 6 o_din0_1[13]
port 304 nsew signal output
rlabel metal2 s 138386 165721 138442 166521 6 o_din0_1[14]
port 305 nsew signal output
rlabel metal2 s 139306 165721 139362 166521 6 o_din0_1[15]
port 306 nsew signal output
rlabel metal3 s 163577 114792 164377 114912 6 o_din0_1[16]
port 307 nsew signal output
rlabel metal2 s 144734 165721 144790 166521 6 o_din0_1[17]
port 308 nsew signal output
rlabel metal2 s 148874 0 148930 800 6 o_din0_1[18]
port 309 nsew signal output
rlabel metal3 s 0 83104 800 83224 6 o_din0_1[19]
port 310 nsew signal output
rlabel metal3 s 163577 28160 164377 28280 6 o_din0_1[1]
port 311 nsew signal output
rlabel metal2 s 152646 0 152702 800 6 o_din0_1[20]
port 312 nsew signal output
rlabel metal2 s 156418 0 156474 800 6 o_din0_1[21]
port 313 nsew signal output
rlabel metal3 s 163577 134784 164377 134904 6 o_din0_1[22]
port 314 nsew signal output
rlabel metal3 s 0 102824 800 102944 6 o_din0_1[23]
port 315 nsew signal output
rlabel metal3 s 0 111392 800 111512 6 o_din0_1[24]
port 316 nsew signal output
rlabel metal3 s 0 116968 800 117088 6 o_din0_1[25]
port 317 nsew signal output
rlabel metal3 s 0 122680 800 122800 6 o_din0_1[26]
port 318 nsew signal output
rlabel metal3 s 163577 151376 164377 151496 6 o_din0_1[27]
port 319 nsew signal output
rlabel metal2 s 162950 0 163006 800 6 o_din0_1[28]
port 320 nsew signal output
rlabel metal3 s 0 142400 800 142520 6 o_din0_1[29]
port 321 nsew signal output
rlabel metal2 s 112258 0 112314 800 6 o_din0_1[2]
port 322 nsew signal output
rlabel metal2 s 162950 165721 163006 166521 6 o_din0_1[30]
port 323 nsew signal output
rlabel metal3 s 0 162120 800 162240 6 o_din0_1[31]
port 324 nsew signal output
rlabel metal3 s 0 23808 800 23928 6 o_din0_1[3]
port 325 nsew signal output
rlabel metal2 s 117502 165721 117558 166521 6 o_din0_1[4]
port 326 nsew signal output
rlabel metal2 s 120262 165721 120318 166521 6 o_din0_1[5]
port 327 nsew signal output
rlabel metal2 s 122930 165721 122986 166521 6 o_din0_1[6]
port 328 nsew signal output
rlabel metal2 s 124770 165721 124826 166521 6 o_din0_1[7]
port 329 nsew signal output
rlabel metal2 s 126610 165721 126666 166521 6 o_din0_1[8]
port 330 nsew signal output
rlabel metal2 s 131026 0 131082 800 6 o_din0_1[9]
port 331 nsew signal output
rlabel metal3 s 0 9800 800 9920 6 o_waddr0[0]
port 332 nsew signal output
rlabel metal3 s 163577 31560 164377 31680 6 o_waddr0[1]
port 333 nsew signal output
rlabel metal2 s 115018 0 115074 800 6 o_waddr0[2]
port 334 nsew signal output
rlabel metal3 s 0 29520 800 29640 6 o_waddr0[3]
port 335 nsew signal output
rlabel metal3 s 163577 44888 164377 45008 6 o_waddr0[4]
port 336 nsew signal output
rlabel metal2 s 123482 0 123538 800 6 o_waddr0[5]
port 337 nsew signal output
rlabel metal3 s 0 46384 800 46504 6 o_waddr0[6]
port 338 nsew signal output
rlabel metal3 s 163577 78208 164377 78328 6 o_waddr0[7]
port 339 nsew signal output
rlabel metal2 s 128450 165721 128506 166521 6 o_waddr0[8]
port 340 nsew signal output
rlabel metal2 s 104714 0 104770 800 6 o_waddr0_1[0]
port 341 nsew signal output
rlabel metal2 s 111154 165721 111210 166521 6 o_waddr0_1[1]
port 342 nsew signal output
rlabel metal2 s 114098 0 114154 800 6 o_waddr0_1[2]
port 343 nsew signal output
rlabel metal3 s 0 26664 800 26784 6 o_waddr0_1[3]
port 344 nsew signal output
rlabel metal3 s 0 37952 800 38072 6 o_waddr0_1[4]
port 345 nsew signal output
rlabel metal3 s 0 40808 800 40928 6 o_waddr0_1[5]
port 346 nsew signal output
rlabel metal3 s 163577 64880 164377 65000 6 o_waddr0_1[6]
port 347 nsew signal output
rlabel metal3 s 163577 74808 164377 74928 6 o_waddr0_1[7]
port 348 nsew signal output
rlabel metal3 s 163577 88136 164377 88256 6 o_waddr0_1[8]
port 349 nsew signal output
rlabel metal3 s 0 4088 800 4208 6 o_web0
port 350 nsew signal output
rlabel metal2 s 102874 0 102930 800 6 o_web0_1
port 351 nsew signal output
rlabel metal2 s 107566 165721 107622 166521 6 o_wmask0[0]
port 352 nsew signal output
rlabel metal2 s 107566 0 107622 800 6 o_wmask0[1]
port 353 nsew signal output
rlabel metal2 s 112074 165721 112130 166521 6 o_wmask0[2]
port 354 nsew signal output
rlabel metal2 s 117870 0 117926 800 6 o_wmask0[3]
port 355 nsew signal output
rlabel metal3 s 163577 18232 164377 18352 6 o_wmask0_1[0]
port 356 nsew signal output
rlabel metal2 s 106554 0 106610 800 6 o_wmask0_1[1]
port 357 nsew signal output
rlabel metal3 s 0 21088 800 21208 6 o_wmask0_1[2]
port 358 nsew signal output
rlabel metal3 s 0 32376 800 32496 6 o_wmask0_1[3]
port 359 nsew signal output
rlabel metal4 s 4208 2128 4528 164336 6 vccd1
port 360 nsew power input
rlabel metal4 s 34928 2128 35248 164336 6 vccd1
port 360 nsew power input
rlabel metal4 s 65648 2128 65968 164336 6 vccd1
port 360 nsew power input
rlabel metal4 s 96368 2128 96688 164336 6 vccd1
port 360 nsew power input
rlabel metal4 s 127088 2128 127408 164336 6 vccd1
port 360 nsew power input
rlabel metal4 s 157808 2128 158128 164336 6 vccd1
port 360 nsew power input
rlabel metal4 s 19568 2128 19888 164336 6 vssd1
port 361 nsew ground input
rlabel metal4 s 50288 2128 50608 164336 6 vssd1
port 361 nsew ground input
rlabel metal4 s 81008 2128 81328 164336 6 vssd1
port 361 nsew ground input
rlabel metal4 s 111728 2128 112048 164336 6 vssd1
port 361 nsew ground input
rlabel metal4 s 142448 2128 142768 164336 6 vssd1
port 361 nsew ground input
rlabel metal2 s 478 0 534 800 6 wb_clk_i
port 362 nsew signal input
rlabel metal2 s 1398 0 1454 800 6 wb_rst_i
port 363 nsew signal input
rlabel metal2 s 2318 0 2374 800 6 wbs_ack_o
port 364 nsew signal output
rlabel metal2 s 6090 0 6146 800 6 wbs_adr_i[0]
port 365 nsew signal input
rlabel metal2 s 38014 0 38070 800 6 wbs_adr_i[10]
port 366 nsew signal input
rlabel metal2 s 40866 0 40922 800 6 wbs_adr_i[11]
port 367 nsew signal input
rlabel metal2 s 43626 0 43682 800 6 wbs_adr_i[12]
port 368 nsew signal input
rlabel metal2 s 46478 0 46534 800 6 wbs_adr_i[13]
port 369 nsew signal input
rlabel metal2 s 49238 0 49294 800 6 wbs_adr_i[14]
port 370 nsew signal input
rlabel metal2 s 52090 0 52146 800 6 wbs_adr_i[15]
port 371 nsew signal input
rlabel metal2 s 54942 0 54998 800 6 wbs_adr_i[16]
port 372 nsew signal input
rlabel metal2 s 57702 0 57758 800 6 wbs_adr_i[17]
port 373 nsew signal input
rlabel metal2 s 60554 0 60610 800 6 wbs_adr_i[18]
port 374 nsew signal input
rlabel metal2 s 63406 0 63462 800 6 wbs_adr_i[19]
port 375 nsew signal input
rlabel metal2 s 9862 0 9918 800 6 wbs_adr_i[1]
port 376 nsew signal input
rlabel metal2 s 66166 0 66222 800 6 wbs_adr_i[20]
port 377 nsew signal input
rlabel metal2 s 69018 0 69074 800 6 wbs_adr_i[21]
port 378 nsew signal input
rlabel metal2 s 71870 0 71926 800 6 wbs_adr_i[22]
port 379 nsew signal input
rlabel metal2 s 74630 0 74686 800 6 wbs_adr_i[23]
port 380 nsew signal input
rlabel metal2 s 77482 0 77538 800 6 wbs_adr_i[24]
port 381 nsew signal input
rlabel metal2 s 80242 0 80298 800 6 wbs_adr_i[25]
port 382 nsew signal input
rlabel metal2 s 83094 0 83150 800 6 wbs_adr_i[26]
port 383 nsew signal input
rlabel metal2 s 85946 0 86002 800 6 wbs_adr_i[27]
port 384 nsew signal input
rlabel metal2 s 88706 0 88762 800 6 wbs_adr_i[28]
port 385 nsew signal input
rlabel metal2 s 91558 0 91614 800 6 wbs_adr_i[29]
port 386 nsew signal input
rlabel metal2 s 13542 0 13598 800 6 wbs_adr_i[2]
port 387 nsew signal input
rlabel metal2 s 94410 0 94466 800 6 wbs_adr_i[30]
port 388 nsew signal input
rlabel metal2 s 97170 0 97226 800 6 wbs_adr_i[31]
port 389 nsew signal input
rlabel metal2 s 17314 0 17370 800 6 wbs_adr_i[3]
port 390 nsew signal input
rlabel metal2 s 21086 0 21142 800 6 wbs_adr_i[4]
port 391 nsew signal input
rlabel metal2 s 23938 0 23994 800 6 wbs_adr_i[5]
port 392 nsew signal input
rlabel metal2 s 26698 0 26754 800 6 wbs_adr_i[6]
port 393 nsew signal input
rlabel metal2 s 29550 0 29606 800 6 wbs_adr_i[7]
port 394 nsew signal input
rlabel metal2 s 32402 0 32458 800 6 wbs_adr_i[8]
port 395 nsew signal input
rlabel metal2 s 35162 0 35218 800 6 wbs_adr_i[9]
port 396 nsew signal input
rlabel metal2 s 3238 0 3294 800 6 wbs_cyc_i
port 397 nsew signal input
rlabel metal2 s 7010 0 7066 800 6 wbs_dat_i[0]
port 398 nsew signal input
rlabel metal2 s 38934 0 38990 800 6 wbs_dat_i[10]
port 399 nsew signal input
rlabel metal2 s 41786 0 41842 800 6 wbs_dat_i[11]
port 400 nsew signal input
rlabel metal2 s 44546 0 44602 800 6 wbs_dat_i[12]
port 401 nsew signal input
rlabel metal2 s 47398 0 47454 800 6 wbs_dat_i[13]
port 402 nsew signal input
rlabel metal2 s 50250 0 50306 800 6 wbs_dat_i[14]
port 403 nsew signal input
rlabel metal2 s 53010 0 53066 800 6 wbs_dat_i[15]
port 404 nsew signal input
rlabel metal2 s 55862 0 55918 800 6 wbs_dat_i[16]
port 405 nsew signal input
rlabel metal2 s 58714 0 58770 800 6 wbs_dat_i[17]
port 406 nsew signal input
rlabel metal2 s 61474 0 61530 800 6 wbs_dat_i[18]
port 407 nsew signal input
rlabel metal2 s 64326 0 64382 800 6 wbs_dat_i[19]
port 408 nsew signal input
rlabel metal2 s 10782 0 10838 800 6 wbs_dat_i[1]
port 409 nsew signal input
rlabel metal2 s 67178 0 67234 800 6 wbs_dat_i[20]
port 410 nsew signal input
rlabel metal2 s 69938 0 69994 800 6 wbs_dat_i[21]
port 411 nsew signal input
rlabel metal2 s 72790 0 72846 800 6 wbs_dat_i[22]
port 412 nsew signal input
rlabel metal2 s 75550 0 75606 800 6 wbs_dat_i[23]
port 413 nsew signal input
rlabel metal2 s 78402 0 78458 800 6 wbs_dat_i[24]
port 414 nsew signal input
rlabel metal2 s 81254 0 81310 800 6 wbs_dat_i[25]
port 415 nsew signal input
rlabel metal2 s 84014 0 84070 800 6 wbs_dat_i[26]
port 416 nsew signal input
rlabel metal2 s 86866 0 86922 800 6 wbs_dat_i[27]
port 417 nsew signal input
rlabel metal2 s 89718 0 89774 800 6 wbs_dat_i[28]
port 418 nsew signal input
rlabel metal2 s 92478 0 92534 800 6 wbs_dat_i[29]
port 419 nsew signal input
rlabel metal2 s 14554 0 14610 800 6 wbs_dat_i[2]
port 420 nsew signal input
rlabel metal2 s 95330 0 95386 800 6 wbs_dat_i[30]
port 421 nsew signal input
rlabel metal2 s 98090 0 98146 800 6 wbs_dat_i[31]
port 422 nsew signal input
rlabel metal2 s 18326 0 18382 800 6 wbs_dat_i[3]
port 423 nsew signal input
rlabel metal2 s 22006 0 22062 800 6 wbs_dat_i[4]
port 424 nsew signal input
rlabel metal2 s 24858 0 24914 800 6 wbs_dat_i[5]
port 425 nsew signal input
rlabel metal2 s 27710 0 27766 800 6 wbs_dat_i[6]
port 426 nsew signal input
rlabel metal2 s 30470 0 30526 800 6 wbs_dat_i[7]
port 427 nsew signal input
rlabel metal2 s 33322 0 33378 800 6 wbs_dat_i[8]
port 428 nsew signal input
rlabel metal2 s 36174 0 36230 800 6 wbs_dat_i[9]
port 429 nsew signal input
rlabel metal2 s 7930 0 7986 800 6 wbs_dat_o[0]
port 430 nsew signal output
rlabel metal2 s 39854 0 39910 800 6 wbs_dat_o[10]
port 431 nsew signal output
rlabel metal2 s 42706 0 42762 800 6 wbs_dat_o[11]
port 432 nsew signal output
rlabel metal2 s 45558 0 45614 800 6 wbs_dat_o[12]
port 433 nsew signal output
rlabel metal2 s 48318 0 48374 800 6 wbs_dat_o[13]
port 434 nsew signal output
rlabel metal2 s 51170 0 51226 800 6 wbs_dat_o[14]
port 435 nsew signal output
rlabel metal2 s 54022 0 54078 800 6 wbs_dat_o[15]
port 436 nsew signal output
rlabel metal2 s 56782 0 56838 800 6 wbs_dat_o[16]
port 437 nsew signal output
rlabel metal2 s 59634 0 59690 800 6 wbs_dat_o[17]
port 438 nsew signal output
rlabel metal2 s 62394 0 62450 800 6 wbs_dat_o[18]
port 439 nsew signal output
rlabel metal2 s 65246 0 65302 800 6 wbs_dat_o[19]
port 440 nsew signal output
rlabel metal2 s 11702 0 11758 800 6 wbs_dat_o[1]
port 441 nsew signal output
rlabel metal2 s 68098 0 68154 800 6 wbs_dat_o[20]
port 442 nsew signal output
rlabel metal2 s 70858 0 70914 800 6 wbs_dat_o[21]
port 443 nsew signal output
rlabel metal2 s 73710 0 73766 800 6 wbs_dat_o[22]
port 444 nsew signal output
rlabel metal2 s 76562 0 76618 800 6 wbs_dat_o[23]
port 445 nsew signal output
rlabel metal2 s 79322 0 79378 800 6 wbs_dat_o[24]
port 446 nsew signal output
rlabel metal2 s 82174 0 82230 800 6 wbs_dat_o[25]
port 447 nsew signal output
rlabel metal2 s 85026 0 85082 800 6 wbs_dat_o[26]
port 448 nsew signal output
rlabel metal2 s 87786 0 87842 800 6 wbs_dat_o[27]
port 449 nsew signal output
rlabel metal2 s 90638 0 90694 800 6 wbs_dat_o[28]
port 450 nsew signal output
rlabel metal2 s 93398 0 93454 800 6 wbs_dat_o[29]
port 451 nsew signal output
rlabel metal2 s 15474 0 15530 800 6 wbs_dat_o[2]
port 452 nsew signal output
rlabel metal2 s 96250 0 96306 800 6 wbs_dat_o[30]
port 453 nsew signal output
rlabel metal2 s 99102 0 99158 800 6 wbs_dat_o[31]
port 454 nsew signal output
rlabel metal2 s 19246 0 19302 800 6 wbs_dat_o[3]
port 455 nsew signal output
rlabel metal2 s 23018 0 23074 800 6 wbs_dat_o[4]
port 456 nsew signal output
rlabel metal2 s 25778 0 25834 800 6 wbs_dat_o[5]
port 457 nsew signal output
rlabel metal2 s 28630 0 28686 800 6 wbs_dat_o[6]
port 458 nsew signal output
rlabel metal2 s 31390 0 31446 800 6 wbs_dat_o[7]
port 459 nsew signal output
rlabel metal2 s 34242 0 34298 800 6 wbs_dat_o[8]
port 460 nsew signal output
rlabel metal2 s 37094 0 37150 800 6 wbs_dat_o[9]
port 461 nsew signal output
rlabel metal2 s 8850 0 8906 800 6 wbs_sel_i[0]
port 462 nsew signal input
rlabel metal2 s 12622 0 12678 800 6 wbs_sel_i[1]
port 463 nsew signal input
rlabel metal2 s 16394 0 16450 800 6 wbs_sel_i[2]
port 464 nsew signal input
rlabel metal2 s 20166 0 20222 800 6 wbs_sel_i[3]
port 465 nsew signal input
rlabel metal2 s 4158 0 4214 800 6 wbs_stb_i
port 466 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 wbs_we_i
port 467 nsew signal input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 164377 166521
string LEFview TRUE
string GDS_FILE /local/caravel_user_project/openlane/user_proj/runs/user_proj/results/magic/user_proj.gds
string GDS_END 78792886
string GDS_START 1347634
<< end >>

