magic
tech sky130A
magscale 1 2
timestamp 1640767669
<< obsli1 >>
rect 1409 1581 165295 167059
<< obsm1 >>
rect 566 552 165307 167544
<< metal2 >>
rect 478 166914 534 167714
rect 1490 166914 1546 167714
rect 2594 166914 2650 167714
rect 3606 166914 3662 167714
rect 4710 166914 4766 167714
rect 5814 166914 5870 167714
rect 6826 166914 6882 167714
rect 7930 166914 7986 167714
rect 8942 166914 8998 167714
rect 10046 166914 10102 167714
rect 11150 166914 11206 167714
rect 12162 166914 12218 167714
rect 13266 166914 13322 167714
rect 14278 166914 14334 167714
rect 15382 166914 15438 167714
rect 16486 166914 16542 167714
rect 17498 166914 17554 167714
rect 18602 166914 18658 167714
rect 19706 166914 19762 167714
rect 20718 166914 20774 167714
rect 21822 166914 21878 167714
rect 22834 166914 22890 167714
rect 23938 166914 23994 167714
rect 25042 166914 25098 167714
rect 26054 166914 26110 167714
rect 27158 166914 27214 167714
rect 28170 166914 28226 167714
rect 29274 166914 29330 167714
rect 30378 166914 30434 167714
rect 31390 166914 31446 167714
rect 32494 166914 32550 167714
rect 33598 166914 33654 167714
rect 34610 166914 34666 167714
rect 35714 166914 35770 167714
rect 36726 166914 36782 167714
rect 37830 166914 37886 167714
rect 38934 166914 38990 167714
rect 39946 166914 40002 167714
rect 41050 166914 41106 167714
rect 42062 166914 42118 167714
rect 43166 166914 43222 167714
rect 44270 166914 44326 167714
rect 45282 166914 45338 167714
rect 46386 166914 46442 167714
rect 47398 166914 47454 167714
rect 48502 166914 48558 167714
rect 49606 166914 49662 167714
rect 50618 166914 50674 167714
rect 51722 166914 51778 167714
rect 52826 166914 52882 167714
rect 53838 166914 53894 167714
rect 54942 166914 54998 167714
rect 55954 166914 56010 167714
rect 57058 166914 57114 167714
rect 58162 166914 58218 167714
rect 59174 166914 59230 167714
rect 60278 166914 60334 167714
rect 61290 166914 61346 167714
rect 62394 166914 62450 167714
rect 63498 166914 63554 167714
rect 64510 166914 64566 167714
rect 65614 166914 65670 167714
rect 66718 166914 66774 167714
rect 67730 166914 67786 167714
rect 68834 166914 68890 167714
rect 69846 166914 69902 167714
rect 70950 166914 71006 167714
rect 72054 166914 72110 167714
rect 73066 166914 73122 167714
rect 74170 166914 74226 167714
rect 75182 166914 75238 167714
rect 76286 166914 76342 167714
rect 77390 166914 77446 167714
rect 78402 166914 78458 167714
rect 79506 166914 79562 167714
rect 80518 166914 80574 167714
rect 81622 166914 81678 167714
rect 82726 166914 82782 167714
rect 83738 166914 83794 167714
rect 84842 166914 84898 167714
rect 85946 166914 86002 167714
rect 86958 166914 87014 167714
rect 88062 166914 88118 167714
rect 89074 166914 89130 167714
rect 90178 166914 90234 167714
rect 91282 166914 91338 167714
rect 92294 166914 92350 167714
rect 93398 166914 93454 167714
rect 94410 166914 94466 167714
rect 95514 166914 95570 167714
rect 96618 166914 96674 167714
rect 97630 166914 97686 167714
rect 98734 166914 98790 167714
rect 99838 166914 99894 167714
rect 100850 166914 100906 167714
rect 101954 166914 102010 167714
rect 102966 166914 103022 167714
rect 104070 166914 104126 167714
rect 105174 166914 105230 167714
rect 106186 166914 106242 167714
rect 107290 166914 107346 167714
rect 108302 166914 108358 167714
rect 109406 166914 109462 167714
rect 110510 166914 110566 167714
rect 111522 166914 111578 167714
rect 112626 166914 112682 167714
rect 113638 166914 113694 167714
rect 114742 166914 114798 167714
rect 115846 166914 115902 167714
rect 116858 166914 116914 167714
rect 117962 166914 118018 167714
rect 119066 166914 119122 167714
rect 120078 166914 120134 167714
rect 121182 166914 121238 167714
rect 122194 166914 122250 167714
rect 123298 166914 123354 167714
rect 124402 166914 124458 167714
rect 125414 166914 125470 167714
rect 126518 166914 126574 167714
rect 127530 166914 127586 167714
rect 128634 166914 128690 167714
rect 129738 166914 129794 167714
rect 130750 166914 130806 167714
rect 131854 166914 131910 167714
rect 132958 166914 133014 167714
rect 133970 166914 134026 167714
rect 135074 166914 135130 167714
rect 136086 166914 136142 167714
rect 137190 166914 137246 167714
rect 138294 166914 138350 167714
rect 139306 166914 139362 167714
rect 140410 166914 140466 167714
rect 141422 166914 141478 167714
rect 142526 166914 142582 167714
rect 143630 166914 143686 167714
rect 144642 166914 144698 167714
rect 145746 166914 145802 167714
rect 146758 166914 146814 167714
rect 147862 166914 147918 167714
rect 148966 166914 149022 167714
rect 149978 166914 150034 167714
rect 151082 166914 151138 167714
rect 152186 166914 152242 167714
rect 153198 166914 153254 167714
rect 154302 166914 154358 167714
rect 155314 166914 155370 167714
rect 156418 166914 156474 167714
rect 157522 166914 157578 167714
rect 158534 166914 158590 167714
rect 159638 166914 159694 167714
rect 160650 166914 160706 167714
rect 161754 166914 161810 167714
rect 162858 166914 162914 167714
rect 163870 166914 163926 167714
rect 164974 166914 165030 167714
rect 570 0 626 800
rect 1674 0 1730 800
rect 2778 0 2834 800
rect 3974 0 4030 800
rect 5078 0 5134 800
rect 6274 0 6330 800
rect 7378 0 7434 800
rect 8482 0 8538 800
rect 9678 0 9734 800
rect 10782 0 10838 800
rect 11978 0 12034 800
rect 13082 0 13138 800
rect 14186 0 14242 800
rect 15382 0 15438 800
rect 16486 0 16542 800
rect 17682 0 17738 800
rect 18786 0 18842 800
rect 19982 0 20038 800
rect 21086 0 21142 800
rect 22190 0 22246 800
rect 23386 0 23442 800
rect 24490 0 24546 800
rect 25686 0 25742 800
rect 26790 0 26846 800
rect 27894 0 27950 800
rect 29090 0 29146 800
rect 30194 0 30250 800
rect 31390 0 31446 800
rect 32494 0 32550 800
rect 33690 0 33746 800
rect 34794 0 34850 800
rect 35898 0 35954 800
rect 37094 0 37150 800
rect 38198 0 38254 800
rect 39394 0 39450 800
rect 40498 0 40554 800
rect 41602 0 41658 800
rect 42798 0 42854 800
rect 43902 0 43958 800
rect 45098 0 45154 800
rect 46202 0 46258 800
rect 47306 0 47362 800
rect 48502 0 48558 800
rect 49606 0 49662 800
rect 50802 0 50858 800
rect 51906 0 51962 800
rect 53102 0 53158 800
rect 54206 0 54262 800
rect 55310 0 55366 800
rect 56506 0 56562 800
rect 57610 0 57666 800
rect 58806 0 58862 800
rect 59910 0 59966 800
rect 61014 0 61070 800
rect 62210 0 62266 800
rect 63314 0 63370 800
rect 64510 0 64566 800
rect 65614 0 65670 800
rect 66810 0 66866 800
rect 67914 0 67970 800
rect 69018 0 69074 800
rect 70214 0 70270 800
rect 71318 0 71374 800
rect 72514 0 72570 800
rect 73618 0 73674 800
rect 74722 0 74778 800
rect 75918 0 75974 800
rect 77022 0 77078 800
rect 78218 0 78274 800
rect 79322 0 79378 800
rect 80426 0 80482 800
rect 81622 0 81678 800
rect 82726 0 82782 800
rect 83922 0 83978 800
rect 85026 0 85082 800
rect 86222 0 86278 800
rect 87326 0 87382 800
rect 88430 0 88486 800
rect 89626 0 89682 800
rect 90730 0 90786 800
rect 91926 0 91982 800
rect 93030 0 93086 800
rect 94134 0 94190 800
rect 95330 0 95386 800
rect 96434 0 96490 800
rect 97630 0 97686 800
rect 98734 0 98790 800
rect 99930 0 99986 800
rect 101034 0 101090 800
rect 102138 0 102194 800
rect 103334 0 103390 800
rect 104438 0 104494 800
rect 105634 0 105690 800
rect 106738 0 106794 800
rect 107842 0 107898 800
rect 109038 0 109094 800
rect 110142 0 110198 800
rect 111338 0 111394 800
rect 112442 0 112498 800
rect 113546 0 113602 800
rect 114742 0 114798 800
rect 115846 0 115902 800
rect 117042 0 117098 800
rect 118146 0 118202 800
rect 119342 0 119398 800
rect 120446 0 120502 800
rect 121550 0 121606 800
rect 122746 0 122802 800
rect 123850 0 123906 800
rect 125046 0 125102 800
rect 126150 0 126206 800
rect 127254 0 127310 800
rect 128450 0 128506 800
rect 129554 0 129610 800
rect 130750 0 130806 800
rect 131854 0 131910 800
rect 133050 0 133106 800
rect 134154 0 134210 800
rect 135258 0 135314 800
rect 136454 0 136510 800
rect 137558 0 137614 800
rect 138754 0 138810 800
rect 139858 0 139914 800
rect 140962 0 141018 800
rect 142158 0 142214 800
rect 143262 0 143318 800
rect 144458 0 144514 800
rect 145562 0 145618 800
rect 146666 0 146722 800
rect 147862 0 147918 800
rect 148966 0 149022 800
rect 150162 0 150218 800
rect 151266 0 151322 800
rect 152462 0 152518 800
rect 153566 0 153622 800
rect 154670 0 154726 800
rect 155866 0 155922 800
rect 156970 0 157026 800
rect 158166 0 158222 800
rect 159270 0 159326 800
rect 160374 0 160430 800
rect 161570 0 161626 800
rect 162674 0 162730 800
rect 163870 0 163926 800
rect 164974 0 165030 800
<< obsm2 >>
rect 590 166858 1434 167550
rect 1602 166858 2538 167550
rect 2706 166858 3550 167550
rect 3718 166858 4654 167550
rect 4822 166858 5758 167550
rect 5926 166858 6770 167550
rect 6938 166858 7874 167550
rect 8042 166858 8886 167550
rect 9054 166858 9990 167550
rect 10158 166858 11094 167550
rect 11262 166858 12106 167550
rect 12274 166858 13210 167550
rect 13378 166858 14222 167550
rect 14390 166858 15326 167550
rect 15494 166858 16430 167550
rect 16598 166858 17442 167550
rect 17610 166858 18546 167550
rect 18714 166858 19650 167550
rect 19818 166858 20662 167550
rect 20830 166858 21766 167550
rect 21934 166858 22778 167550
rect 22946 166858 23882 167550
rect 24050 166858 24986 167550
rect 25154 166858 25998 167550
rect 26166 166858 27102 167550
rect 27270 166858 28114 167550
rect 28282 166858 29218 167550
rect 29386 166858 30322 167550
rect 30490 166858 31334 167550
rect 31502 166858 32438 167550
rect 32606 166858 33542 167550
rect 33710 166858 34554 167550
rect 34722 166858 35658 167550
rect 35826 166858 36670 167550
rect 36838 166858 37774 167550
rect 37942 166858 38878 167550
rect 39046 166858 39890 167550
rect 40058 166858 40994 167550
rect 41162 166858 42006 167550
rect 42174 166858 43110 167550
rect 43278 166858 44214 167550
rect 44382 166858 45226 167550
rect 45394 166858 46330 167550
rect 46498 166858 47342 167550
rect 47510 166858 48446 167550
rect 48614 166858 49550 167550
rect 49718 166858 50562 167550
rect 50730 166858 51666 167550
rect 51834 166858 52770 167550
rect 52938 166858 53782 167550
rect 53950 166858 54886 167550
rect 55054 166858 55898 167550
rect 56066 166858 57002 167550
rect 57170 166858 58106 167550
rect 58274 166858 59118 167550
rect 59286 166858 60222 167550
rect 60390 166858 61234 167550
rect 61402 166858 62338 167550
rect 62506 166858 63442 167550
rect 63610 166858 64454 167550
rect 64622 166858 65558 167550
rect 65726 166858 66662 167550
rect 66830 166858 67674 167550
rect 67842 166858 68778 167550
rect 68946 166858 69790 167550
rect 69958 166858 70894 167550
rect 71062 166858 71998 167550
rect 72166 166858 73010 167550
rect 73178 166858 74114 167550
rect 74282 166858 75126 167550
rect 75294 166858 76230 167550
rect 76398 166858 77334 167550
rect 77502 166858 78346 167550
rect 78514 166858 79450 167550
rect 79618 166858 80462 167550
rect 80630 166858 81566 167550
rect 81734 166858 82670 167550
rect 82838 166858 83682 167550
rect 83850 166858 84786 167550
rect 84954 166858 85890 167550
rect 86058 166858 86902 167550
rect 87070 166858 88006 167550
rect 88174 166858 89018 167550
rect 89186 166858 90122 167550
rect 90290 166858 91226 167550
rect 91394 166858 92238 167550
rect 92406 166858 93342 167550
rect 93510 166858 94354 167550
rect 94522 166858 95458 167550
rect 95626 166858 96562 167550
rect 96730 166858 97574 167550
rect 97742 166858 98678 167550
rect 98846 166858 99782 167550
rect 99950 166858 100794 167550
rect 100962 166858 101898 167550
rect 102066 166858 102910 167550
rect 103078 166858 104014 167550
rect 104182 166858 105118 167550
rect 105286 166858 106130 167550
rect 106298 166858 107234 167550
rect 107402 166858 108246 167550
rect 108414 166858 109350 167550
rect 109518 166858 110454 167550
rect 110622 166858 111466 167550
rect 111634 166858 112570 167550
rect 112738 166858 113582 167550
rect 113750 166858 114686 167550
rect 114854 166858 115790 167550
rect 115958 166858 116802 167550
rect 116970 166858 117906 167550
rect 118074 166858 119010 167550
rect 119178 166858 120022 167550
rect 120190 166858 121126 167550
rect 121294 166858 122138 167550
rect 122306 166858 123242 167550
rect 123410 166858 124346 167550
rect 124514 166858 125358 167550
rect 125526 166858 126462 167550
rect 126630 166858 127474 167550
rect 127642 166858 128578 167550
rect 128746 166858 129682 167550
rect 129850 166858 130694 167550
rect 130862 166858 131798 167550
rect 131966 166858 132902 167550
rect 133070 166858 133914 167550
rect 134082 166858 135018 167550
rect 135186 166858 136030 167550
rect 136198 166858 137134 167550
rect 137302 166858 138238 167550
rect 138406 166858 139250 167550
rect 139418 166858 140354 167550
rect 140522 166858 141366 167550
rect 141534 166858 142470 167550
rect 142638 166858 143574 167550
rect 143742 166858 144586 167550
rect 144754 166858 145690 167550
rect 145858 166858 146702 167550
rect 146870 166858 147806 167550
rect 147974 166858 148910 167550
rect 149078 166858 149922 167550
rect 150090 166858 151026 167550
rect 151194 166858 152130 167550
rect 152298 166858 153142 167550
rect 153310 166858 154246 167550
rect 154414 166858 155258 167550
rect 155426 166858 156362 167550
rect 156530 166858 157466 167550
rect 157634 166858 158478 167550
rect 158646 166858 159582 167550
rect 159750 166858 160594 167550
rect 160762 166858 161698 167550
rect 161866 166858 162802 167550
rect 162970 166858 163814 167550
rect 163982 166858 164918 167550
rect 570 856 165028 166858
rect 682 546 1618 856
rect 1786 546 2722 856
rect 2890 546 3918 856
rect 4086 546 5022 856
rect 5190 546 6218 856
rect 6386 546 7322 856
rect 7490 546 8426 856
rect 8594 546 9622 856
rect 9790 546 10726 856
rect 10894 546 11922 856
rect 12090 546 13026 856
rect 13194 546 14130 856
rect 14298 546 15326 856
rect 15494 546 16430 856
rect 16598 546 17626 856
rect 17794 546 18730 856
rect 18898 546 19926 856
rect 20094 546 21030 856
rect 21198 546 22134 856
rect 22302 546 23330 856
rect 23498 546 24434 856
rect 24602 546 25630 856
rect 25798 546 26734 856
rect 26902 546 27838 856
rect 28006 546 29034 856
rect 29202 546 30138 856
rect 30306 546 31334 856
rect 31502 546 32438 856
rect 32606 546 33634 856
rect 33802 546 34738 856
rect 34906 546 35842 856
rect 36010 546 37038 856
rect 37206 546 38142 856
rect 38310 546 39338 856
rect 39506 546 40442 856
rect 40610 546 41546 856
rect 41714 546 42742 856
rect 42910 546 43846 856
rect 44014 546 45042 856
rect 45210 546 46146 856
rect 46314 546 47250 856
rect 47418 546 48446 856
rect 48614 546 49550 856
rect 49718 546 50746 856
rect 50914 546 51850 856
rect 52018 546 53046 856
rect 53214 546 54150 856
rect 54318 546 55254 856
rect 55422 546 56450 856
rect 56618 546 57554 856
rect 57722 546 58750 856
rect 58918 546 59854 856
rect 60022 546 60958 856
rect 61126 546 62154 856
rect 62322 546 63258 856
rect 63426 546 64454 856
rect 64622 546 65558 856
rect 65726 546 66754 856
rect 66922 546 67858 856
rect 68026 546 68962 856
rect 69130 546 70158 856
rect 70326 546 71262 856
rect 71430 546 72458 856
rect 72626 546 73562 856
rect 73730 546 74666 856
rect 74834 546 75862 856
rect 76030 546 76966 856
rect 77134 546 78162 856
rect 78330 546 79266 856
rect 79434 546 80370 856
rect 80538 546 81566 856
rect 81734 546 82670 856
rect 82838 546 83866 856
rect 84034 546 84970 856
rect 85138 546 86166 856
rect 86334 546 87270 856
rect 87438 546 88374 856
rect 88542 546 89570 856
rect 89738 546 90674 856
rect 90842 546 91870 856
rect 92038 546 92974 856
rect 93142 546 94078 856
rect 94246 546 95274 856
rect 95442 546 96378 856
rect 96546 546 97574 856
rect 97742 546 98678 856
rect 98846 546 99874 856
rect 100042 546 100978 856
rect 101146 546 102082 856
rect 102250 546 103278 856
rect 103446 546 104382 856
rect 104550 546 105578 856
rect 105746 546 106682 856
rect 106850 546 107786 856
rect 107954 546 108982 856
rect 109150 546 110086 856
rect 110254 546 111282 856
rect 111450 546 112386 856
rect 112554 546 113490 856
rect 113658 546 114686 856
rect 114854 546 115790 856
rect 115958 546 116986 856
rect 117154 546 118090 856
rect 118258 546 119286 856
rect 119454 546 120390 856
rect 120558 546 121494 856
rect 121662 546 122690 856
rect 122858 546 123794 856
rect 123962 546 124990 856
rect 125158 546 126094 856
rect 126262 546 127198 856
rect 127366 546 128394 856
rect 128562 546 129498 856
rect 129666 546 130694 856
rect 130862 546 131798 856
rect 131966 546 132994 856
rect 133162 546 134098 856
rect 134266 546 135202 856
rect 135370 546 136398 856
rect 136566 546 137502 856
rect 137670 546 138698 856
rect 138866 546 139802 856
rect 139970 546 140906 856
rect 141074 546 142102 856
rect 142270 546 143206 856
rect 143374 546 144402 856
rect 144570 546 145506 856
rect 145674 546 146610 856
rect 146778 546 147806 856
rect 147974 546 148910 856
rect 149078 546 150106 856
rect 150274 546 151210 856
rect 151378 546 152406 856
rect 152574 546 153510 856
rect 153678 546 154614 856
rect 154782 546 155810 856
rect 155978 546 156914 856
rect 157082 546 158110 856
rect 158278 546 159214 856
rect 159382 546 160318 856
rect 160486 546 161514 856
rect 161682 546 162618 856
rect 162786 546 163814 856
rect 163982 546 164918 856
<< metal3 >>
rect 164770 165928 165570 166048
rect 0 164976 800 165096
rect 164770 162664 165570 162784
rect 0 159672 800 159792
rect 164770 159400 165570 159520
rect 164770 156136 165570 156256
rect 0 154504 800 154624
rect 164770 152872 165570 152992
rect 164770 149472 165570 149592
rect 0 149200 800 149320
rect 164770 146208 165570 146328
rect 0 144032 800 144152
rect 164770 142944 165570 143064
rect 164770 139680 165570 139800
rect 0 138728 800 138848
rect 164770 136416 165570 136536
rect 0 133560 800 133680
rect 164770 133152 165570 133272
rect 164770 129752 165570 129872
rect 0 128256 800 128376
rect 164770 126488 165570 126608
rect 0 123088 800 123208
rect 164770 123224 165570 123344
rect 164770 119960 165570 120080
rect 0 117784 800 117904
rect 164770 116696 165570 116816
rect 164770 113432 165570 113552
rect 0 112616 800 112736
rect 164770 110032 165570 110152
rect 0 107312 800 107432
rect 164770 106768 165570 106888
rect 164770 103504 165570 103624
rect 0 102144 800 102264
rect 164770 100240 165570 100360
rect 0 96840 800 96960
rect 164770 96976 165570 97096
rect 164770 93576 165570 93696
rect 0 91672 800 91792
rect 164770 90312 165570 90432
rect 164770 87048 165570 87168
rect 0 86368 800 86488
rect 164770 83784 165570 83904
rect 0 81064 800 81184
rect 164770 80520 165570 80640
rect 164770 77256 165570 77376
rect 0 75896 800 76016
rect 164770 73856 165570 73976
rect 0 70592 800 70712
rect 164770 70592 165570 70712
rect 164770 67328 165570 67448
rect 0 65424 800 65544
rect 164770 64064 165570 64184
rect 164770 60800 165570 60920
rect 0 60120 800 60240
rect 164770 57536 165570 57656
rect 0 54952 800 55072
rect 164770 54136 165570 54256
rect 164770 50872 165570 50992
rect 0 49648 800 49768
rect 164770 47608 165570 47728
rect 0 44480 800 44600
rect 164770 44344 165570 44464
rect 164770 41080 165570 41200
rect 0 39176 800 39296
rect 164770 37680 165570 37800
rect 164770 34416 165570 34536
rect 0 34008 800 34128
rect 164770 31152 165570 31272
rect 0 28704 800 28824
rect 164770 27888 165570 28008
rect 164770 24624 165570 24744
rect 0 23536 800 23656
rect 164770 21360 165570 21480
rect 0 18232 800 18352
rect 164770 17960 165570 18080
rect 164770 14696 165570 14816
rect 0 13064 800 13184
rect 164770 11432 165570 11552
rect 164770 8168 165570 8288
rect 0 7760 800 7880
rect 164770 4904 165570 5024
rect 0 2592 800 2712
rect 164770 1640 165570 1760
<< obsm3 >>
rect 565 166128 164943 167245
rect 565 165848 164690 166128
rect 565 165176 164943 165848
rect 880 164896 164943 165176
rect 565 162864 164943 164896
rect 565 162584 164690 162864
rect 565 159872 164943 162584
rect 880 159600 164943 159872
rect 880 159592 164690 159600
rect 565 159320 164690 159592
rect 565 156336 164943 159320
rect 565 156056 164690 156336
rect 565 154704 164943 156056
rect 880 154424 164943 154704
rect 565 153072 164943 154424
rect 565 152792 164690 153072
rect 565 149672 164943 152792
rect 565 149400 164690 149672
rect 880 149392 164690 149400
rect 880 149120 164943 149392
rect 565 146408 164943 149120
rect 565 146128 164690 146408
rect 565 144232 164943 146128
rect 880 143952 164943 144232
rect 565 143144 164943 143952
rect 565 142864 164690 143144
rect 565 139880 164943 142864
rect 565 139600 164690 139880
rect 565 138928 164943 139600
rect 880 138648 164943 138928
rect 565 136616 164943 138648
rect 565 136336 164690 136616
rect 565 133760 164943 136336
rect 880 133480 164943 133760
rect 565 133352 164943 133480
rect 565 133072 164690 133352
rect 565 129952 164943 133072
rect 565 129672 164690 129952
rect 565 128456 164943 129672
rect 880 128176 164943 128456
rect 565 126688 164943 128176
rect 565 126408 164690 126688
rect 565 123424 164943 126408
rect 565 123288 164690 123424
rect 880 123144 164690 123288
rect 880 123008 164943 123144
rect 565 120160 164943 123008
rect 565 119880 164690 120160
rect 565 117984 164943 119880
rect 880 117704 164943 117984
rect 565 116896 164943 117704
rect 565 116616 164690 116896
rect 565 113632 164943 116616
rect 565 113352 164690 113632
rect 565 112816 164943 113352
rect 880 112536 164943 112816
rect 565 110232 164943 112536
rect 565 109952 164690 110232
rect 565 107512 164943 109952
rect 880 107232 164943 107512
rect 565 106968 164943 107232
rect 565 106688 164690 106968
rect 565 103704 164943 106688
rect 565 103424 164690 103704
rect 565 102344 164943 103424
rect 880 102064 164943 102344
rect 565 100440 164943 102064
rect 565 100160 164690 100440
rect 565 97176 164943 100160
rect 565 97040 164690 97176
rect 880 96896 164690 97040
rect 880 96760 164943 96896
rect 565 93776 164943 96760
rect 565 93496 164690 93776
rect 565 91872 164943 93496
rect 880 91592 164943 91872
rect 565 90512 164943 91592
rect 565 90232 164690 90512
rect 565 87248 164943 90232
rect 565 86968 164690 87248
rect 565 86568 164943 86968
rect 880 86288 164943 86568
rect 565 83984 164943 86288
rect 565 83704 164690 83984
rect 565 81264 164943 83704
rect 880 80984 164943 81264
rect 565 80720 164943 80984
rect 565 80440 164690 80720
rect 565 77456 164943 80440
rect 565 77176 164690 77456
rect 565 76096 164943 77176
rect 880 75816 164943 76096
rect 565 74056 164943 75816
rect 565 73776 164690 74056
rect 565 70792 164943 73776
rect 880 70512 164690 70792
rect 565 67528 164943 70512
rect 565 67248 164690 67528
rect 565 65624 164943 67248
rect 880 65344 164943 65624
rect 565 64264 164943 65344
rect 565 63984 164690 64264
rect 565 61000 164943 63984
rect 565 60720 164690 61000
rect 565 60320 164943 60720
rect 880 60040 164943 60320
rect 565 57736 164943 60040
rect 565 57456 164690 57736
rect 565 55152 164943 57456
rect 880 54872 164943 55152
rect 565 54336 164943 54872
rect 565 54056 164690 54336
rect 565 51072 164943 54056
rect 565 50792 164690 51072
rect 565 49848 164943 50792
rect 880 49568 164943 49848
rect 565 47808 164943 49568
rect 565 47528 164690 47808
rect 565 44680 164943 47528
rect 880 44544 164943 44680
rect 880 44400 164690 44544
rect 565 44264 164690 44400
rect 565 41280 164943 44264
rect 565 41000 164690 41280
rect 565 39376 164943 41000
rect 880 39096 164943 39376
rect 565 37880 164943 39096
rect 565 37600 164690 37880
rect 565 34616 164943 37600
rect 565 34336 164690 34616
rect 565 34208 164943 34336
rect 880 33928 164943 34208
rect 565 31352 164943 33928
rect 565 31072 164690 31352
rect 565 28904 164943 31072
rect 880 28624 164943 28904
rect 565 28088 164943 28624
rect 565 27808 164690 28088
rect 565 24824 164943 27808
rect 565 24544 164690 24824
rect 565 23736 164943 24544
rect 880 23456 164943 23736
rect 565 21560 164943 23456
rect 565 21280 164690 21560
rect 565 18432 164943 21280
rect 880 18160 164943 18432
rect 880 18152 164690 18160
rect 565 17880 164690 18152
rect 565 14896 164943 17880
rect 565 14616 164690 14896
rect 565 13264 164943 14616
rect 880 12984 164943 13264
rect 565 11632 164943 12984
rect 565 11352 164690 11632
rect 565 8368 164943 11352
rect 565 8088 164690 8368
rect 565 7960 164943 8088
rect 880 7680 164943 7960
rect 565 5104 164943 7680
rect 565 4824 164690 5104
rect 565 2792 164943 4824
rect 880 2512 164943 2792
rect 565 1840 164943 2512
rect 565 1560 164690 1840
rect 565 1259 164943 1560
<< metal4 >>
rect 4208 2128 4528 165424
rect 19568 2128 19888 165424
rect 34928 2128 35248 165424
rect 50288 2128 50608 165424
rect 65648 2128 65968 165424
rect 81008 2128 81328 165424
rect 96368 2128 96688 165424
rect 111728 2128 112048 165424
rect 127088 2128 127408 165424
rect 142448 2128 142768 165424
rect 157808 2128 158128 165424
<< obsm4 >>
rect 3371 165504 162781 167245
rect 3371 2048 4128 165504
rect 4608 2048 19488 165504
rect 19968 2048 34848 165504
rect 35328 2048 50208 165504
rect 50688 2048 65568 165504
rect 66048 2048 80928 165504
rect 81408 2048 96288 165504
rect 96768 2048 111648 165504
rect 112128 2048 127008 165504
rect 127488 2048 142368 165504
rect 142848 2048 157728 165504
rect 158208 2048 162781 165504
rect 3371 1259 162781 2048
<< labels >>
rlabel metal2 s 122194 166914 122250 167714 6 clk_i
port 1 nsew signal input
rlabel metal2 s 126150 0 126206 800 6 i_dout0[0]
port 2 nsew signal input
rlabel metal3 s 164770 87048 165570 87168 6 i_dout0[10]
port 3 nsew signal input
rlabel metal2 s 143630 166914 143686 167714 6 i_dout0[11]
port 4 nsew signal input
rlabel metal3 s 164770 96976 165570 97096 6 i_dout0[12]
port 5 nsew signal input
rlabel metal2 s 145562 0 145618 800 6 i_dout0[13]
port 6 nsew signal input
rlabel metal2 s 148966 166914 149022 167714 6 i_dout0[14]
port 7 nsew signal input
rlabel metal3 s 164770 100240 165570 100360 6 i_dout0[15]
port 8 nsew signal input
rlabel metal2 s 151082 166914 151138 167714 6 i_dout0[16]
port 9 nsew signal input
rlabel metal2 s 151266 0 151322 800 6 i_dout0[17]
port 10 nsew signal input
rlabel metal2 s 152186 166914 152242 167714 6 i_dout0[18]
port 11 nsew signal input
rlabel metal3 s 0 96840 800 96960 6 i_dout0[19]
port 12 nsew signal input
rlabel metal2 s 126518 166914 126574 167714 6 i_dout0[1]
port 13 nsew signal input
rlabel metal3 s 0 102144 800 102264 6 i_dout0[20]
port 14 nsew signal input
rlabel metal3 s 164770 123224 165570 123344 6 i_dout0[21]
port 15 nsew signal input
rlabel metal3 s 164770 129752 165570 129872 6 i_dout0[22]
port 16 nsew signal input
rlabel metal2 s 158166 0 158222 800 6 i_dout0[23]
port 17 nsew signal input
rlabel metal3 s 164770 136416 165570 136536 6 i_dout0[24]
port 18 nsew signal input
rlabel metal3 s 0 133560 800 133680 6 i_dout0[25]
port 19 nsew signal input
rlabel metal3 s 0 144032 800 144152 6 i_dout0[26]
port 20 nsew signal input
rlabel metal2 s 158534 166914 158590 167714 6 i_dout0[27]
port 21 nsew signal input
rlabel metal2 s 159638 166914 159694 167714 6 i_dout0[28]
port 22 nsew signal input
rlabel metal2 s 160650 166914 160706 167714 6 i_dout0[29]
port 23 nsew signal input
rlabel metal3 s 164770 27888 165570 28008 6 i_dout0[2]
port 24 nsew signal input
rlabel metal3 s 164770 156136 165570 156256 6 i_dout0[30]
port 25 nsew signal input
rlabel metal3 s 0 164976 800 165096 6 i_dout0[31]
port 26 nsew signal input
rlabel metal2 s 130750 166914 130806 167714 6 i_dout0[3]
port 27 nsew signal input
rlabel metal2 s 131854 166914 131910 167714 6 i_dout0[4]
port 28 nsew signal input
rlabel metal2 s 132958 166914 133014 167714 6 i_dout0[5]
port 29 nsew signal input
rlabel metal3 s 0 44480 800 44600 6 i_dout0[6]
port 30 nsew signal input
rlabel metal2 s 142158 0 142214 800 6 i_dout0[7]
port 31 nsew signal input
rlabel metal2 s 143262 0 143318 800 6 i_dout0[8]
port 32 nsew signal input
rlabel metal3 s 164770 77256 165570 77376 6 i_dout0[9]
port 33 nsew signal input
rlabel metal2 s 127254 0 127310 800 6 i_dout0_1[0]
port 34 nsew signal input
rlabel metal3 s 164770 83784 165570 83904 6 i_dout0_1[10]
port 35 nsew signal input
rlabel metal3 s 0 60120 800 60240 6 i_dout0_1[11]
port 36 nsew signal input
rlabel metal2 s 144642 166914 144698 167714 6 i_dout0_1[12]
port 37 nsew signal input
rlabel metal2 s 146758 166914 146814 167714 6 i_dout0_1[13]
port 38 nsew signal input
rlabel metal3 s 0 70592 800 70712 6 i_dout0_1[14]
port 39 nsew signal input
rlabel metal3 s 0 75896 800 76016 6 i_dout0_1[15]
port 40 nsew signal input
rlabel metal3 s 0 81064 800 81184 6 i_dout0_1[16]
port 41 nsew signal input
rlabel metal2 s 150162 0 150218 800 6 i_dout0_1[17]
port 42 nsew signal input
rlabel metal2 s 152462 0 152518 800 6 i_dout0_1[18]
port 43 nsew signal input
rlabel metal3 s 164770 113432 165570 113552 6 i_dout0_1[19]
port 44 nsew signal input
rlabel metal2 s 125414 166914 125470 167714 6 i_dout0_1[1]
port 45 nsew signal input
rlabel metal3 s 164770 119960 165570 120080 6 i_dout0_1[20]
port 46 nsew signal input
rlabel metal2 s 154302 166914 154358 167714 6 i_dout0_1[21]
port 47 nsew signal input
rlabel metal2 s 156970 0 157026 800 6 i_dout0_1[22]
port 48 nsew signal input
rlabel metal2 s 156418 166914 156474 167714 6 i_dout0_1[23]
port 49 nsew signal input
rlabel metal3 s 164770 133152 165570 133272 6 i_dout0_1[24]
port 50 nsew signal input
rlabel metal3 s 164770 146208 165570 146328 6 i_dout0_1[25]
port 51 nsew signal input
rlabel metal2 s 159270 0 159326 800 6 i_dout0_1[26]
port 52 nsew signal input
rlabel metal2 s 161570 0 161626 800 6 i_dout0_1[27]
port 53 nsew signal input
rlabel metal2 s 163870 0 163926 800 6 i_dout0_1[28]
port 54 nsew signal input
rlabel metal3 s 0 159672 800 159792 6 i_dout0_1[29]
port 55 nsew signal input
rlabel metal3 s 164770 24624 165570 24744 6 i_dout0_1[2]
port 56 nsew signal input
rlabel metal2 s 162858 166914 162914 167714 6 i_dout0_1[30]
port 57 nsew signal input
rlabel metal2 s 163870 166914 163926 167714 6 i_dout0_1[31]
port 58 nsew signal input
rlabel metal2 s 131854 0 131910 800 6 i_dout0_1[3]
port 59 nsew signal input
rlabel metal3 s 0 34008 800 34128 6 i_dout0_1[4]
port 60 nsew signal input
rlabel metal3 s 164770 50872 165570 50992 6 i_dout0_1[5]
port 61 nsew signal input
rlabel metal2 s 138754 0 138810 800 6 i_dout0_1[6]
port 62 nsew signal input
rlabel metal3 s 164770 60800 165570 60920 6 i_dout0_1[7]
port 63 nsew signal input
rlabel metal2 s 138294 166914 138350 167714 6 i_dout0_1[8]
port 64 nsew signal input
rlabel metal2 s 140410 166914 140466 167714 6 i_dout0_1[9]
port 65 nsew signal input
rlabel metal2 s 478 166914 534 167714 6 io_in[0]
port 66 nsew signal input
rlabel metal2 s 32494 166914 32550 167714 6 io_in[10]
port 67 nsew signal input
rlabel metal2 s 35714 166914 35770 167714 6 io_in[11]
port 68 nsew signal input
rlabel metal2 s 38934 166914 38990 167714 6 io_in[12]
port 69 nsew signal input
rlabel metal2 s 42062 166914 42118 167714 6 io_in[13]
port 70 nsew signal input
rlabel metal2 s 45282 166914 45338 167714 6 io_in[14]
port 71 nsew signal input
rlabel metal2 s 48502 166914 48558 167714 6 io_in[15]
port 72 nsew signal input
rlabel metal2 s 51722 166914 51778 167714 6 io_in[16]
port 73 nsew signal input
rlabel metal2 s 54942 166914 54998 167714 6 io_in[17]
port 74 nsew signal input
rlabel metal2 s 58162 166914 58218 167714 6 io_in[18]
port 75 nsew signal input
rlabel metal2 s 61290 166914 61346 167714 6 io_in[19]
port 76 nsew signal input
rlabel metal2 s 3606 166914 3662 167714 6 io_in[1]
port 77 nsew signal input
rlabel metal2 s 64510 166914 64566 167714 6 io_in[20]
port 78 nsew signal input
rlabel metal2 s 67730 166914 67786 167714 6 io_in[21]
port 79 nsew signal input
rlabel metal2 s 70950 166914 71006 167714 6 io_in[22]
port 80 nsew signal input
rlabel metal2 s 74170 166914 74226 167714 6 io_in[23]
port 81 nsew signal input
rlabel metal2 s 77390 166914 77446 167714 6 io_in[24]
port 82 nsew signal input
rlabel metal2 s 80518 166914 80574 167714 6 io_in[25]
port 83 nsew signal input
rlabel metal2 s 83738 166914 83794 167714 6 io_in[26]
port 84 nsew signal input
rlabel metal2 s 86958 166914 87014 167714 6 io_in[27]
port 85 nsew signal input
rlabel metal2 s 90178 166914 90234 167714 6 io_in[28]
port 86 nsew signal input
rlabel metal2 s 93398 166914 93454 167714 6 io_in[29]
port 87 nsew signal input
rlabel metal2 s 6826 166914 6882 167714 6 io_in[2]
port 88 nsew signal input
rlabel metal2 s 96618 166914 96674 167714 6 io_in[30]
port 89 nsew signal input
rlabel metal2 s 99838 166914 99894 167714 6 io_in[31]
port 90 nsew signal input
rlabel metal2 s 102966 166914 103022 167714 6 io_in[32]
port 91 nsew signal input
rlabel metal2 s 106186 166914 106242 167714 6 io_in[33]
port 92 nsew signal input
rlabel metal2 s 109406 166914 109462 167714 6 io_in[34]
port 93 nsew signal input
rlabel metal2 s 112626 166914 112682 167714 6 io_in[35]
port 94 nsew signal input
rlabel metal2 s 115846 166914 115902 167714 6 io_in[36]
port 95 nsew signal input
rlabel metal2 s 119066 166914 119122 167714 6 io_in[37]
port 96 nsew signal input
rlabel metal2 s 10046 166914 10102 167714 6 io_in[3]
port 97 nsew signal input
rlabel metal2 s 13266 166914 13322 167714 6 io_in[4]
port 98 nsew signal input
rlabel metal2 s 16486 166914 16542 167714 6 io_in[5]
port 99 nsew signal input
rlabel metal2 s 19706 166914 19762 167714 6 io_in[6]
port 100 nsew signal input
rlabel metal2 s 22834 166914 22890 167714 6 io_in[7]
port 101 nsew signal input
rlabel metal2 s 26054 166914 26110 167714 6 io_in[8]
port 102 nsew signal input
rlabel metal2 s 29274 166914 29330 167714 6 io_in[9]
port 103 nsew signal input
rlabel metal2 s 1490 166914 1546 167714 6 io_oeb[0]
port 104 nsew signal output
rlabel metal2 s 33598 166914 33654 167714 6 io_oeb[10]
port 105 nsew signal output
rlabel metal2 s 36726 166914 36782 167714 6 io_oeb[11]
port 106 nsew signal output
rlabel metal2 s 39946 166914 40002 167714 6 io_oeb[12]
port 107 nsew signal output
rlabel metal2 s 43166 166914 43222 167714 6 io_oeb[13]
port 108 nsew signal output
rlabel metal2 s 46386 166914 46442 167714 6 io_oeb[14]
port 109 nsew signal output
rlabel metal2 s 49606 166914 49662 167714 6 io_oeb[15]
port 110 nsew signal output
rlabel metal2 s 52826 166914 52882 167714 6 io_oeb[16]
port 111 nsew signal output
rlabel metal2 s 55954 166914 56010 167714 6 io_oeb[17]
port 112 nsew signal output
rlabel metal2 s 59174 166914 59230 167714 6 io_oeb[18]
port 113 nsew signal output
rlabel metal2 s 62394 166914 62450 167714 6 io_oeb[19]
port 114 nsew signal output
rlabel metal2 s 4710 166914 4766 167714 6 io_oeb[1]
port 115 nsew signal output
rlabel metal2 s 65614 166914 65670 167714 6 io_oeb[20]
port 116 nsew signal output
rlabel metal2 s 68834 166914 68890 167714 6 io_oeb[21]
port 117 nsew signal output
rlabel metal2 s 72054 166914 72110 167714 6 io_oeb[22]
port 118 nsew signal output
rlabel metal2 s 75182 166914 75238 167714 6 io_oeb[23]
port 119 nsew signal output
rlabel metal2 s 78402 166914 78458 167714 6 io_oeb[24]
port 120 nsew signal output
rlabel metal2 s 81622 166914 81678 167714 6 io_oeb[25]
port 121 nsew signal output
rlabel metal2 s 84842 166914 84898 167714 6 io_oeb[26]
port 122 nsew signal output
rlabel metal2 s 88062 166914 88118 167714 6 io_oeb[27]
port 123 nsew signal output
rlabel metal2 s 91282 166914 91338 167714 6 io_oeb[28]
port 124 nsew signal output
rlabel metal2 s 94410 166914 94466 167714 6 io_oeb[29]
port 125 nsew signal output
rlabel metal2 s 7930 166914 7986 167714 6 io_oeb[2]
port 126 nsew signal output
rlabel metal2 s 97630 166914 97686 167714 6 io_oeb[30]
port 127 nsew signal output
rlabel metal2 s 100850 166914 100906 167714 6 io_oeb[31]
port 128 nsew signal output
rlabel metal2 s 104070 166914 104126 167714 6 io_oeb[32]
port 129 nsew signal output
rlabel metal2 s 107290 166914 107346 167714 6 io_oeb[33]
port 130 nsew signal output
rlabel metal2 s 110510 166914 110566 167714 6 io_oeb[34]
port 131 nsew signal output
rlabel metal2 s 113638 166914 113694 167714 6 io_oeb[35]
port 132 nsew signal output
rlabel metal2 s 116858 166914 116914 167714 6 io_oeb[36]
port 133 nsew signal output
rlabel metal2 s 120078 166914 120134 167714 6 io_oeb[37]
port 134 nsew signal output
rlabel metal2 s 11150 166914 11206 167714 6 io_oeb[3]
port 135 nsew signal output
rlabel metal2 s 14278 166914 14334 167714 6 io_oeb[4]
port 136 nsew signal output
rlabel metal2 s 17498 166914 17554 167714 6 io_oeb[5]
port 137 nsew signal output
rlabel metal2 s 20718 166914 20774 167714 6 io_oeb[6]
port 138 nsew signal output
rlabel metal2 s 23938 166914 23994 167714 6 io_oeb[7]
port 139 nsew signal output
rlabel metal2 s 27158 166914 27214 167714 6 io_oeb[8]
port 140 nsew signal output
rlabel metal2 s 30378 166914 30434 167714 6 io_oeb[9]
port 141 nsew signal output
rlabel metal2 s 2594 166914 2650 167714 6 io_out[0]
port 142 nsew signal output
rlabel metal2 s 34610 166914 34666 167714 6 io_out[10]
port 143 nsew signal output
rlabel metal2 s 37830 166914 37886 167714 6 io_out[11]
port 144 nsew signal output
rlabel metal2 s 41050 166914 41106 167714 6 io_out[12]
port 145 nsew signal output
rlabel metal2 s 44270 166914 44326 167714 6 io_out[13]
port 146 nsew signal output
rlabel metal2 s 47398 166914 47454 167714 6 io_out[14]
port 147 nsew signal output
rlabel metal2 s 50618 166914 50674 167714 6 io_out[15]
port 148 nsew signal output
rlabel metal2 s 53838 166914 53894 167714 6 io_out[16]
port 149 nsew signal output
rlabel metal2 s 57058 166914 57114 167714 6 io_out[17]
port 150 nsew signal output
rlabel metal2 s 60278 166914 60334 167714 6 io_out[18]
port 151 nsew signal output
rlabel metal2 s 63498 166914 63554 167714 6 io_out[19]
port 152 nsew signal output
rlabel metal2 s 5814 166914 5870 167714 6 io_out[1]
port 153 nsew signal output
rlabel metal2 s 66718 166914 66774 167714 6 io_out[20]
port 154 nsew signal output
rlabel metal2 s 69846 166914 69902 167714 6 io_out[21]
port 155 nsew signal output
rlabel metal2 s 73066 166914 73122 167714 6 io_out[22]
port 156 nsew signal output
rlabel metal2 s 76286 166914 76342 167714 6 io_out[23]
port 157 nsew signal output
rlabel metal2 s 79506 166914 79562 167714 6 io_out[24]
port 158 nsew signal output
rlabel metal2 s 82726 166914 82782 167714 6 io_out[25]
port 159 nsew signal output
rlabel metal2 s 85946 166914 86002 167714 6 io_out[26]
port 160 nsew signal output
rlabel metal2 s 89074 166914 89130 167714 6 io_out[27]
port 161 nsew signal output
rlabel metal2 s 92294 166914 92350 167714 6 io_out[28]
port 162 nsew signal output
rlabel metal2 s 95514 166914 95570 167714 6 io_out[29]
port 163 nsew signal output
rlabel metal2 s 8942 166914 8998 167714 6 io_out[2]
port 164 nsew signal output
rlabel metal2 s 98734 166914 98790 167714 6 io_out[30]
port 165 nsew signal output
rlabel metal2 s 101954 166914 102010 167714 6 io_out[31]
port 166 nsew signal output
rlabel metal2 s 105174 166914 105230 167714 6 io_out[32]
port 167 nsew signal output
rlabel metal2 s 108302 166914 108358 167714 6 io_out[33]
port 168 nsew signal output
rlabel metal2 s 111522 166914 111578 167714 6 io_out[34]
port 169 nsew signal output
rlabel metal2 s 114742 166914 114798 167714 6 io_out[35]
port 170 nsew signal output
rlabel metal2 s 117962 166914 118018 167714 6 io_out[36]
port 171 nsew signal output
rlabel metal2 s 121182 166914 121238 167714 6 io_out[37]
port 172 nsew signal output
rlabel metal2 s 12162 166914 12218 167714 6 io_out[3]
port 173 nsew signal output
rlabel metal2 s 15382 166914 15438 167714 6 io_out[4]
port 174 nsew signal output
rlabel metal2 s 18602 166914 18658 167714 6 io_out[5]
port 175 nsew signal output
rlabel metal2 s 21822 166914 21878 167714 6 io_out[6]
port 176 nsew signal output
rlabel metal2 s 25042 166914 25098 167714 6 io_out[7]
port 177 nsew signal output
rlabel metal2 s 28170 166914 28226 167714 6 io_out[8]
port 178 nsew signal output
rlabel metal2 s 31390 166914 31446 167714 6 io_out[9]
port 179 nsew signal output
rlabel metal2 s 121550 0 121606 800 6 irq[0]
port 180 nsew signal output
rlabel metal2 s 122746 0 122802 800 6 irq[1]
port 181 nsew signal output
rlabel metal2 s 123850 0 123906 800 6 irq[2]
port 182 nsew signal output
rlabel metal2 s 123298 166914 123354 167714 6 o_csb0
port 183 nsew signal output
rlabel metal3 s 164770 1640 165570 1760 6 o_csb0_1
port 184 nsew signal output
rlabel metal3 s 164770 8168 165570 8288 6 o_din0[0]
port 185 nsew signal output
rlabel metal3 s 164770 90312 165570 90432 6 o_din0[10]
port 186 nsew signal output
rlabel metal3 s 164770 93576 165570 93696 6 o_din0[11]
port 187 nsew signal output
rlabel metal2 s 145746 166914 145802 167714 6 o_din0[12]
port 188 nsew signal output
rlabel metal2 s 147862 166914 147918 167714 6 o_din0[13]
port 189 nsew signal output
rlabel metal2 s 149978 166914 150034 167714 6 o_din0[14]
port 190 nsew signal output
rlabel metal3 s 164770 103504 165570 103624 6 o_din0[15]
port 191 nsew signal output
rlabel metal3 s 164770 106768 165570 106888 6 o_din0[16]
port 192 nsew signal output
rlabel metal3 s 164770 110032 165570 110152 6 o_din0[17]
port 193 nsew signal output
rlabel metal2 s 154670 0 154726 800 6 o_din0[18]
port 194 nsew signal output
rlabel metal2 s 155866 0 155922 800 6 o_din0[19]
port 195 nsew signal output
rlabel metal2 s 127530 166914 127586 167714 6 o_din0[1]
port 196 nsew signal output
rlabel metal2 s 153198 166914 153254 167714 6 o_din0[20]
port 197 nsew signal output
rlabel metal3 s 0 112616 800 112736 6 o_din0[21]
port 198 nsew signal output
rlabel metal2 s 155314 166914 155370 167714 6 o_din0[22]
port 199 nsew signal output
rlabel metal3 s 0 128256 800 128376 6 o_din0[23]
port 200 nsew signal output
rlabel metal3 s 164770 142944 165570 143064 6 o_din0[24]
port 201 nsew signal output
rlabel metal3 s 0 138728 800 138848 6 o_din0[25]
port 202 nsew signal output
rlabel metal2 s 157522 166914 157578 167714 6 o_din0[26]
port 203 nsew signal output
rlabel metal2 s 162674 0 162730 800 6 o_din0[27]
port 204 nsew signal output
rlabel metal2 s 164974 0 165030 800 6 o_din0[28]
port 205 nsew signal output
rlabel metal3 s 164770 152872 165570 152992 6 o_din0[29]
port 206 nsew signal output
rlabel metal3 s 0 23536 800 23656 6 o_din0[2]
port 207 nsew signal output
rlabel metal3 s 164770 162664 165570 162784 6 o_din0[30]
port 208 nsew signal output
rlabel metal2 s 164974 166914 165030 167714 6 o_din0[31]
port 209 nsew signal output
rlabel metal2 s 133050 0 133106 800 6 o_din0[3]
port 210 nsew signal output
rlabel metal2 s 136454 0 136510 800 6 o_din0[4]
port 211 nsew signal output
rlabel metal2 s 137558 0 137614 800 6 o_din0[5]
port 212 nsew signal output
rlabel metal3 s 164770 57536 165570 57656 6 o_din0[6]
port 213 nsew signal output
rlabel metal2 s 137190 166914 137246 167714 6 o_din0[7]
port 214 nsew signal output
rlabel metal3 s 164770 70592 165570 70712 6 o_din0[8]
port 215 nsew signal output
rlabel metal2 s 141422 166914 141478 167714 6 o_din0[9]
port 216 nsew signal output
rlabel metal3 s 164770 11432 165570 11552 6 o_din0_1[0]
port 217 nsew signal output
rlabel metal2 s 142526 166914 142582 167714 6 o_din0_1[10]
port 218 nsew signal output
rlabel metal3 s 0 65424 800 65544 6 o_din0_1[11]
port 219 nsew signal output
rlabel metal2 s 144458 0 144514 800 6 o_din0_1[12]
port 220 nsew signal output
rlabel metal2 s 146666 0 146722 800 6 o_din0_1[13]
port 221 nsew signal output
rlabel metal2 s 147862 0 147918 800 6 o_din0_1[14]
port 222 nsew signal output
rlabel metal2 s 148966 0 149022 800 6 o_din0_1[15]
port 223 nsew signal output
rlabel metal3 s 0 86368 800 86488 6 o_din0_1[16]
port 224 nsew signal output
rlabel metal3 s 0 91672 800 91792 6 o_din0_1[17]
port 225 nsew signal output
rlabel metal2 s 153566 0 153622 800 6 o_din0_1[18]
port 226 nsew signal output
rlabel metal3 s 164770 116696 165570 116816 6 o_din0_1[19]
port 227 nsew signal output
rlabel metal3 s 0 2592 800 2712 6 o_din0_1[1]
port 228 nsew signal output
rlabel metal3 s 0 107312 800 107432 6 o_din0_1[20]
port 229 nsew signal output
rlabel metal3 s 164770 126488 165570 126608 6 o_din0_1[21]
port 230 nsew signal output
rlabel metal3 s 0 117784 800 117904 6 o_din0_1[22]
port 231 nsew signal output
rlabel metal3 s 0 123088 800 123208 6 o_din0_1[23]
port 232 nsew signal output
rlabel metal3 s 164770 139680 165570 139800 6 o_din0_1[24]
port 233 nsew signal output
rlabel metal3 s 164770 149472 165570 149592 6 o_din0_1[25]
port 234 nsew signal output
rlabel metal2 s 160374 0 160430 800 6 o_din0_1[26]
port 235 nsew signal output
rlabel metal3 s 0 149200 800 149320 6 o_din0_1[27]
port 236 nsew signal output
rlabel metal3 s 0 154504 800 154624 6 o_din0_1[28]
port 237 nsew signal output
rlabel metal2 s 161754 166914 161810 167714 6 o_din0_1[29]
port 238 nsew signal output
rlabel metal2 s 130750 0 130806 800 6 o_din0_1[2]
port 239 nsew signal output
rlabel metal3 s 164770 159400 165570 159520 6 o_din0_1[30]
port 240 nsew signal output
rlabel metal3 s 164770 165928 165570 166048 6 o_din0_1[31]
port 241 nsew signal output
rlabel metal3 s 164770 34416 165570 34536 6 o_din0_1[3]
port 242 nsew signal output
rlabel metal2 s 135258 0 135314 800 6 o_din0_1[4]
port 243 nsew signal output
rlabel metal2 s 133970 166914 134026 167714 6 o_din0_1[5]
port 244 nsew signal output
rlabel metal3 s 0 49648 800 49768 6 o_din0_1[6]
port 245 nsew signal output
rlabel metal2 s 136086 166914 136142 167714 6 o_din0_1[7]
port 246 nsew signal output
rlabel metal3 s 164770 67328 165570 67448 6 o_din0_1[8]
port 247 nsew signal output
rlabel metal3 s 164770 80520 165570 80640 6 o_din0_1[9]
port 248 nsew signal output
rlabel metal2 s 128450 0 128506 800 6 o_waddr0[0]
port 249 nsew signal output
rlabel metal3 s 0 7760 800 7880 6 o_waddr0[1]
port 250 nsew signal output
rlabel metal2 s 128634 166914 128690 167714 6 o_waddr0[2]
port 251 nsew signal output
rlabel metal3 s 164770 41080 165570 41200 6 o_waddr0[3]
port 252 nsew signal output
rlabel metal3 s 0 39176 800 39296 6 o_waddr0[4]
port 253 nsew signal output
rlabel metal2 s 135074 166914 135130 167714 6 o_waddr0[5]
port 254 nsew signal output
rlabel metal2 s 140962 0 141018 800 6 o_waddr0[6]
port 255 nsew signal output
rlabel metal3 s 0 54952 800 55072 6 o_waddr0[7]
port 256 nsew signal output
rlabel metal3 s 164770 73856 165570 73976 6 o_waddr0[8]
port 257 nsew signal output
rlabel metal3 s 164770 14696 165570 14816 6 o_waddr0_1[0]
port 258 nsew signal output
rlabel metal3 s 164770 21360 165570 21480 6 o_waddr0_1[1]
port 259 nsew signal output
rlabel metal3 s 164770 31152 165570 31272 6 o_waddr0_1[2]
port 260 nsew signal output
rlabel metal3 s 164770 37680 165570 37800 6 o_waddr0_1[3]
port 261 nsew signal output
rlabel metal3 s 164770 47608 165570 47728 6 o_waddr0_1[4]
port 262 nsew signal output
rlabel metal3 s 164770 54136 165570 54256 6 o_waddr0_1[5]
port 263 nsew signal output
rlabel metal2 s 139858 0 139914 800 6 o_waddr0_1[6]
port 264 nsew signal output
rlabel metal3 s 164770 64064 165570 64184 6 o_waddr0_1[7]
port 265 nsew signal output
rlabel metal2 s 139306 166914 139362 167714 6 o_waddr0_1[8]
port 266 nsew signal output
rlabel metal2 s 125046 0 125102 800 6 o_web0
port 267 nsew signal output
rlabel metal2 s 124402 166914 124458 167714 6 o_web0_1
port 268 nsew signal output
rlabel metal3 s 164770 17960 165570 18080 6 o_wmask0[0]
port 269 nsew signal output
rlabel metal3 s 0 18232 800 18352 6 o_wmask0[1]
port 270 nsew signal output
rlabel metal3 s 0 28704 800 28824 6 o_wmask0[2]
port 271 nsew signal output
rlabel metal3 s 164770 44344 165570 44464 6 o_wmask0[3]
port 272 nsew signal output
rlabel metal2 s 129554 0 129610 800 6 o_wmask0_1[0]
port 273 nsew signal output
rlabel metal3 s 0 13064 800 13184 6 o_wmask0_1[1]
port 274 nsew signal output
rlabel metal2 s 129738 166914 129794 167714 6 o_wmask0_1[2]
port 275 nsew signal output
rlabel metal2 s 134154 0 134210 800 6 o_wmask0_1[3]
port 276 nsew signal output
rlabel metal3 s 164770 4904 165570 5024 6 rst_i
port 277 nsew signal input
rlabel metal4 s 4208 2128 4528 165424 6 vccd1
port 278 nsew power input
rlabel metal4 s 34928 2128 35248 165424 6 vccd1
port 278 nsew power input
rlabel metal4 s 65648 2128 65968 165424 6 vccd1
port 278 nsew power input
rlabel metal4 s 96368 2128 96688 165424 6 vccd1
port 278 nsew power input
rlabel metal4 s 127088 2128 127408 165424 6 vccd1
port 278 nsew power input
rlabel metal4 s 157808 2128 158128 165424 6 vccd1
port 278 nsew power input
rlabel metal4 s 19568 2128 19888 165424 6 vssd1
port 279 nsew ground input
rlabel metal4 s 50288 2128 50608 165424 6 vssd1
port 279 nsew ground input
rlabel metal4 s 81008 2128 81328 165424 6 vssd1
port 279 nsew ground input
rlabel metal4 s 111728 2128 112048 165424 6 vssd1
port 279 nsew ground input
rlabel metal4 s 142448 2128 142768 165424 6 vssd1
port 279 nsew ground input
rlabel metal2 s 570 0 626 800 6 wb_clk_i
port 280 nsew signal input
rlabel metal2 s 1674 0 1730 800 6 wb_rst_i
port 281 nsew signal input
rlabel metal2 s 2778 0 2834 800 6 wbs_ack_o
port 282 nsew signal output
rlabel metal2 s 7378 0 7434 800 6 wbs_adr_i[0]
port 283 nsew signal input
rlabel metal2 s 46202 0 46258 800 6 wbs_adr_i[10]
port 284 nsew signal input
rlabel metal2 s 49606 0 49662 800 6 wbs_adr_i[11]
port 285 nsew signal input
rlabel metal2 s 53102 0 53158 800 6 wbs_adr_i[12]
port 286 nsew signal input
rlabel metal2 s 56506 0 56562 800 6 wbs_adr_i[13]
port 287 nsew signal input
rlabel metal2 s 59910 0 59966 800 6 wbs_adr_i[14]
port 288 nsew signal input
rlabel metal2 s 63314 0 63370 800 6 wbs_adr_i[15]
port 289 nsew signal input
rlabel metal2 s 66810 0 66866 800 6 wbs_adr_i[16]
port 290 nsew signal input
rlabel metal2 s 70214 0 70270 800 6 wbs_adr_i[17]
port 291 nsew signal input
rlabel metal2 s 73618 0 73674 800 6 wbs_adr_i[18]
port 292 nsew signal input
rlabel metal2 s 77022 0 77078 800 6 wbs_adr_i[19]
port 293 nsew signal input
rlabel metal2 s 11978 0 12034 800 6 wbs_adr_i[1]
port 294 nsew signal input
rlabel metal2 s 80426 0 80482 800 6 wbs_adr_i[20]
port 295 nsew signal input
rlabel metal2 s 83922 0 83978 800 6 wbs_adr_i[21]
port 296 nsew signal input
rlabel metal2 s 87326 0 87382 800 6 wbs_adr_i[22]
port 297 nsew signal input
rlabel metal2 s 90730 0 90786 800 6 wbs_adr_i[23]
port 298 nsew signal input
rlabel metal2 s 94134 0 94190 800 6 wbs_adr_i[24]
port 299 nsew signal input
rlabel metal2 s 97630 0 97686 800 6 wbs_adr_i[25]
port 300 nsew signal input
rlabel metal2 s 101034 0 101090 800 6 wbs_adr_i[26]
port 301 nsew signal input
rlabel metal2 s 104438 0 104494 800 6 wbs_adr_i[27]
port 302 nsew signal input
rlabel metal2 s 107842 0 107898 800 6 wbs_adr_i[28]
port 303 nsew signal input
rlabel metal2 s 111338 0 111394 800 6 wbs_adr_i[29]
port 304 nsew signal input
rlabel metal2 s 16486 0 16542 800 6 wbs_adr_i[2]
port 305 nsew signal input
rlabel metal2 s 114742 0 114798 800 6 wbs_adr_i[30]
port 306 nsew signal input
rlabel metal2 s 118146 0 118202 800 6 wbs_adr_i[31]
port 307 nsew signal input
rlabel metal2 s 21086 0 21142 800 6 wbs_adr_i[3]
port 308 nsew signal input
rlabel metal2 s 25686 0 25742 800 6 wbs_adr_i[4]
port 309 nsew signal input
rlabel metal2 s 29090 0 29146 800 6 wbs_adr_i[5]
port 310 nsew signal input
rlabel metal2 s 32494 0 32550 800 6 wbs_adr_i[6]
port 311 nsew signal input
rlabel metal2 s 35898 0 35954 800 6 wbs_adr_i[7]
port 312 nsew signal input
rlabel metal2 s 39394 0 39450 800 6 wbs_adr_i[8]
port 313 nsew signal input
rlabel metal2 s 42798 0 42854 800 6 wbs_adr_i[9]
port 314 nsew signal input
rlabel metal2 s 3974 0 4030 800 6 wbs_cyc_i
port 315 nsew signal input
rlabel metal2 s 8482 0 8538 800 6 wbs_dat_i[0]
port 316 nsew signal input
rlabel metal2 s 47306 0 47362 800 6 wbs_dat_i[10]
port 317 nsew signal input
rlabel metal2 s 50802 0 50858 800 6 wbs_dat_i[11]
port 318 nsew signal input
rlabel metal2 s 54206 0 54262 800 6 wbs_dat_i[12]
port 319 nsew signal input
rlabel metal2 s 57610 0 57666 800 6 wbs_dat_i[13]
port 320 nsew signal input
rlabel metal2 s 61014 0 61070 800 6 wbs_dat_i[14]
port 321 nsew signal input
rlabel metal2 s 64510 0 64566 800 6 wbs_dat_i[15]
port 322 nsew signal input
rlabel metal2 s 67914 0 67970 800 6 wbs_dat_i[16]
port 323 nsew signal input
rlabel metal2 s 71318 0 71374 800 6 wbs_dat_i[17]
port 324 nsew signal input
rlabel metal2 s 74722 0 74778 800 6 wbs_dat_i[18]
port 325 nsew signal input
rlabel metal2 s 78218 0 78274 800 6 wbs_dat_i[19]
port 326 nsew signal input
rlabel metal2 s 13082 0 13138 800 6 wbs_dat_i[1]
port 327 nsew signal input
rlabel metal2 s 81622 0 81678 800 6 wbs_dat_i[20]
port 328 nsew signal input
rlabel metal2 s 85026 0 85082 800 6 wbs_dat_i[21]
port 329 nsew signal input
rlabel metal2 s 88430 0 88486 800 6 wbs_dat_i[22]
port 330 nsew signal input
rlabel metal2 s 91926 0 91982 800 6 wbs_dat_i[23]
port 331 nsew signal input
rlabel metal2 s 95330 0 95386 800 6 wbs_dat_i[24]
port 332 nsew signal input
rlabel metal2 s 98734 0 98790 800 6 wbs_dat_i[25]
port 333 nsew signal input
rlabel metal2 s 102138 0 102194 800 6 wbs_dat_i[26]
port 334 nsew signal input
rlabel metal2 s 105634 0 105690 800 6 wbs_dat_i[27]
port 335 nsew signal input
rlabel metal2 s 109038 0 109094 800 6 wbs_dat_i[28]
port 336 nsew signal input
rlabel metal2 s 112442 0 112498 800 6 wbs_dat_i[29]
port 337 nsew signal input
rlabel metal2 s 17682 0 17738 800 6 wbs_dat_i[2]
port 338 nsew signal input
rlabel metal2 s 115846 0 115902 800 6 wbs_dat_i[30]
port 339 nsew signal input
rlabel metal2 s 119342 0 119398 800 6 wbs_dat_i[31]
port 340 nsew signal input
rlabel metal2 s 22190 0 22246 800 6 wbs_dat_i[3]
port 341 nsew signal input
rlabel metal2 s 26790 0 26846 800 6 wbs_dat_i[4]
port 342 nsew signal input
rlabel metal2 s 30194 0 30250 800 6 wbs_dat_i[5]
port 343 nsew signal input
rlabel metal2 s 33690 0 33746 800 6 wbs_dat_i[6]
port 344 nsew signal input
rlabel metal2 s 37094 0 37150 800 6 wbs_dat_i[7]
port 345 nsew signal input
rlabel metal2 s 40498 0 40554 800 6 wbs_dat_i[8]
port 346 nsew signal input
rlabel metal2 s 43902 0 43958 800 6 wbs_dat_i[9]
port 347 nsew signal input
rlabel metal2 s 9678 0 9734 800 6 wbs_dat_o[0]
port 348 nsew signal output
rlabel metal2 s 48502 0 48558 800 6 wbs_dat_o[10]
port 349 nsew signal output
rlabel metal2 s 51906 0 51962 800 6 wbs_dat_o[11]
port 350 nsew signal output
rlabel metal2 s 55310 0 55366 800 6 wbs_dat_o[12]
port 351 nsew signal output
rlabel metal2 s 58806 0 58862 800 6 wbs_dat_o[13]
port 352 nsew signal output
rlabel metal2 s 62210 0 62266 800 6 wbs_dat_o[14]
port 353 nsew signal output
rlabel metal2 s 65614 0 65670 800 6 wbs_dat_o[15]
port 354 nsew signal output
rlabel metal2 s 69018 0 69074 800 6 wbs_dat_o[16]
port 355 nsew signal output
rlabel metal2 s 72514 0 72570 800 6 wbs_dat_o[17]
port 356 nsew signal output
rlabel metal2 s 75918 0 75974 800 6 wbs_dat_o[18]
port 357 nsew signal output
rlabel metal2 s 79322 0 79378 800 6 wbs_dat_o[19]
port 358 nsew signal output
rlabel metal2 s 14186 0 14242 800 6 wbs_dat_o[1]
port 359 nsew signal output
rlabel metal2 s 82726 0 82782 800 6 wbs_dat_o[20]
port 360 nsew signal output
rlabel metal2 s 86222 0 86278 800 6 wbs_dat_o[21]
port 361 nsew signal output
rlabel metal2 s 89626 0 89682 800 6 wbs_dat_o[22]
port 362 nsew signal output
rlabel metal2 s 93030 0 93086 800 6 wbs_dat_o[23]
port 363 nsew signal output
rlabel metal2 s 96434 0 96490 800 6 wbs_dat_o[24]
port 364 nsew signal output
rlabel metal2 s 99930 0 99986 800 6 wbs_dat_o[25]
port 365 nsew signal output
rlabel metal2 s 103334 0 103390 800 6 wbs_dat_o[26]
port 366 nsew signal output
rlabel metal2 s 106738 0 106794 800 6 wbs_dat_o[27]
port 367 nsew signal output
rlabel metal2 s 110142 0 110198 800 6 wbs_dat_o[28]
port 368 nsew signal output
rlabel metal2 s 113546 0 113602 800 6 wbs_dat_o[29]
port 369 nsew signal output
rlabel metal2 s 18786 0 18842 800 6 wbs_dat_o[2]
port 370 nsew signal output
rlabel metal2 s 117042 0 117098 800 6 wbs_dat_o[30]
port 371 nsew signal output
rlabel metal2 s 120446 0 120502 800 6 wbs_dat_o[31]
port 372 nsew signal output
rlabel metal2 s 23386 0 23442 800 6 wbs_dat_o[3]
port 373 nsew signal output
rlabel metal2 s 27894 0 27950 800 6 wbs_dat_o[4]
port 374 nsew signal output
rlabel metal2 s 31390 0 31446 800 6 wbs_dat_o[5]
port 375 nsew signal output
rlabel metal2 s 34794 0 34850 800 6 wbs_dat_o[6]
port 376 nsew signal output
rlabel metal2 s 38198 0 38254 800 6 wbs_dat_o[7]
port 377 nsew signal output
rlabel metal2 s 41602 0 41658 800 6 wbs_dat_o[8]
port 378 nsew signal output
rlabel metal2 s 45098 0 45154 800 6 wbs_dat_o[9]
port 379 nsew signal output
rlabel metal2 s 10782 0 10838 800 6 wbs_sel_i[0]
port 380 nsew signal input
rlabel metal2 s 15382 0 15438 800 6 wbs_sel_i[1]
port 381 nsew signal input
rlabel metal2 s 19982 0 20038 800 6 wbs_sel_i[2]
port 382 nsew signal input
rlabel metal2 s 24490 0 24546 800 6 wbs_sel_i[3]
port 383 nsew signal input
rlabel metal2 s 5078 0 5134 800 6 wbs_stb_i
port 384 nsew signal input
rlabel metal2 s 6274 0 6330 800 6 wbs_we_i
port 385 nsew signal input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 165570 167714
string LEFview TRUE
string GDS_FILE /project/openlane/user_proj/runs/user_proj/results/magic/user_proj.gds
string GDS_END 72892618
string GDS_START 110
<< end >>

