magic
tech sky130A
magscale 1 2
timestamp 1640319329
<< obsli1 >>
rect 1104 1173 164743 165427
<< obsm1 >>
rect 14 484 164758 165436
<< metal2 >>
rect 478 166124 534 166924
rect 1398 166124 1454 166924
rect 2410 166124 2466 166924
rect 3422 166124 3478 166924
rect 4342 166124 4398 166924
rect 5354 166124 5410 166924
rect 6366 166124 6422 166924
rect 7378 166124 7434 166924
rect 8298 166124 8354 166924
rect 9310 166124 9366 166924
rect 10322 166124 10378 166924
rect 11242 166124 11298 166924
rect 12254 166124 12310 166924
rect 13266 166124 13322 166924
rect 14278 166124 14334 166924
rect 15198 166124 15254 166924
rect 16210 166124 16266 166924
rect 17222 166124 17278 166924
rect 18234 166124 18290 166924
rect 19154 166124 19210 166924
rect 20166 166124 20222 166924
rect 21178 166124 21234 166924
rect 22098 166124 22154 166924
rect 23110 166124 23166 166924
rect 24122 166124 24178 166924
rect 25134 166124 25190 166924
rect 26054 166124 26110 166924
rect 27066 166124 27122 166924
rect 28078 166124 28134 166924
rect 29090 166124 29146 166924
rect 30010 166124 30066 166924
rect 31022 166124 31078 166924
rect 32034 166124 32090 166924
rect 32954 166124 33010 166924
rect 33966 166124 34022 166924
rect 34978 166124 35034 166924
rect 35990 166124 36046 166924
rect 36910 166124 36966 166924
rect 37922 166124 37978 166924
rect 38934 166124 38990 166924
rect 39854 166124 39910 166924
rect 40866 166124 40922 166924
rect 41878 166124 41934 166924
rect 42890 166124 42946 166924
rect 43810 166124 43866 166924
rect 44822 166124 44878 166924
rect 45834 166124 45890 166924
rect 46846 166124 46902 166924
rect 47766 166124 47822 166924
rect 48778 166124 48834 166924
rect 49790 166124 49846 166924
rect 50710 166124 50766 166924
rect 51722 166124 51778 166924
rect 52734 166124 52790 166924
rect 53746 166124 53802 166924
rect 54666 166124 54722 166924
rect 55678 166124 55734 166924
rect 56690 166124 56746 166924
rect 57702 166124 57758 166924
rect 58622 166124 58678 166924
rect 59634 166124 59690 166924
rect 60646 166124 60702 166924
rect 61566 166124 61622 166924
rect 62578 166124 62634 166924
rect 63590 166124 63646 166924
rect 64602 166124 64658 166924
rect 65522 166124 65578 166924
rect 66534 166124 66590 166924
rect 67546 166124 67602 166924
rect 68466 166124 68522 166924
rect 69478 166124 69534 166924
rect 70490 166124 70546 166924
rect 71502 166124 71558 166924
rect 72422 166124 72478 166924
rect 73434 166124 73490 166924
rect 74446 166124 74502 166924
rect 75458 166124 75514 166924
rect 76378 166124 76434 166924
rect 77390 166124 77446 166924
rect 78402 166124 78458 166924
rect 79322 166124 79378 166924
rect 80334 166124 80390 166924
rect 81346 166124 81402 166924
rect 82358 166124 82414 166924
rect 83278 166124 83334 166924
rect 84290 166124 84346 166924
rect 85302 166124 85358 166924
rect 86314 166124 86370 166924
rect 87234 166124 87290 166924
rect 88246 166124 88302 166924
rect 89258 166124 89314 166924
rect 90178 166124 90234 166924
rect 91190 166124 91246 166924
rect 92202 166124 92258 166924
rect 93214 166124 93270 166924
rect 94134 166124 94190 166924
rect 95146 166124 95202 166924
rect 96158 166124 96214 166924
rect 97170 166124 97226 166924
rect 98090 166124 98146 166924
rect 99102 166124 99158 166924
rect 100114 166124 100170 166924
rect 101034 166124 101090 166924
rect 102046 166124 102102 166924
rect 103058 166124 103114 166924
rect 104070 166124 104126 166924
rect 104990 166124 105046 166924
rect 106002 166124 106058 166924
rect 107014 166124 107070 166924
rect 107934 166124 107990 166924
rect 108946 166124 109002 166924
rect 109958 166124 110014 166924
rect 110970 166124 111026 166924
rect 111890 166124 111946 166924
rect 112902 166124 112958 166924
rect 113914 166124 113970 166924
rect 114926 166124 114982 166924
rect 115846 166124 115902 166924
rect 116858 166124 116914 166924
rect 117870 166124 117926 166924
rect 118790 166124 118846 166924
rect 119802 166124 119858 166924
rect 120814 166124 120870 166924
rect 121826 166124 121882 166924
rect 122746 166124 122802 166924
rect 123758 166124 123814 166924
rect 124770 166124 124826 166924
rect 125782 166124 125838 166924
rect 126702 166124 126758 166924
rect 127714 166124 127770 166924
rect 128726 166124 128782 166924
rect 129646 166124 129702 166924
rect 130658 166124 130714 166924
rect 131670 166124 131726 166924
rect 132682 166124 132738 166924
rect 133602 166124 133658 166924
rect 134614 166124 134670 166924
rect 135626 166124 135682 166924
rect 136546 166124 136602 166924
rect 137558 166124 137614 166924
rect 138570 166124 138626 166924
rect 139582 166124 139638 166924
rect 140502 166124 140558 166924
rect 141514 166124 141570 166924
rect 142526 166124 142582 166924
rect 143538 166124 143594 166924
rect 144458 166124 144514 166924
rect 145470 166124 145526 166924
rect 146482 166124 146538 166924
rect 147402 166124 147458 166924
rect 148414 166124 148470 166924
rect 149426 166124 149482 166924
rect 150438 166124 150494 166924
rect 151358 166124 151414 166924
rect 152370 166124 152426 166924
rect 153382 166124 153438 166924
rect 154394 166124 154450 166924
rect 155314 166124 155370 166924
rect 156326 166124 156382 166924
rect 157338 166124 157394 166924
rect 158258 166124 158314 166924
rect 159270 166124 159326 166924
rect 160282 166124 160338 166924
rect 161294 166124 161350 166924
rect 162214 166124 162270 166924
rect 163226 166124 163282 166924
rect 164238 166124 164294 166924
rect 110 0 166 800
rect 386 0 442 800
rect 662 0 718 800
rect 938 0 994 800
rect 1214 0 1270 800
rect 1490 0 1546 800
rect 1858 0 1914 800
rect 2134 0 2190 800
rect 2410 0 2466 800
rect 2686 0 2742 800
rect 2962 0 3018 800
rect 3238 0 3294 800
rect 3606 0 3662 800
rect 3882 0 3938 800
rect 4158 0 4214 800
rect 4434 0 4490 800
rect 4710 0 4766 800
rect 4986 0 5042 800
rect 5354 0 5410 800
rect 5630 0 5686 800
rect 5906 0 5962 800
rect 6182 0 6238 800
rect 6458 0 6514 800
rect 6734 0 6790 800
rect 7102 0 7158 800
rect 7378 0 7434 800
rect 7654 0 7710 800
rect 7930 0 7986 800
rect 8206 0 8262 800
rect 8482 0 8538 800
rect 8850 0 8906 800
rect 9126 0 9182 800
rect 9402 0 9458 800
rect 9678 0 9734 800
rect 9954 0 10010 800
rect 10230 0 10286 800
rect 10598 0 10654 800
rect 10874 0 10930 800
rect 11150 0 11206 800
rect 11426 0 11482 800
rect 11702 0 11758 800
rect 11978 0 12034 800
rect 12346 0 12402 800
rect 12622 0 12678 800
rect 12898 0 12954 800
rect 13174 0 13230 800
rect 13450 0 13506 800
rect 13726 0 13782 800
rect 14094 0 14150 800
rect 14370 0 14426 800
rect 14646 0 14702 800
rect 14922 0 14978 800
rect 15198 0 15254 800
rect 15566 0 15622 800
rect 15842 0 15898 800
rect 16118 0 16174 800
rect 16394 0 16450 800
rect 16670 0 16726 800
rect 16946 0 17002 800
rect 17314 0 17370 800
rect 17590 0 17646 800
rect 17866 0 17922 800
rect 18142 0 18198 800
rect 18418 0 18474 800
rect 18694 0 18750 800
rect 19062 0 19118 800
rect 19338 0 19394 800
rect 19614 0 19670 800
rect 19890 0 19946 800
rect 20166 0 20222 800
rect 20442 0 20498 800
rect 20810 0 20866 800
rect 21086 0 21142 800
rect 21362 0 21418 800
rect 21638 0 21694 800
rect 21914 0 21970 800
rect 22190 0 22246 800
rect 22558 0 22614 800
rect 22834 0 22890 800
rect 23110 0 23166 800
rect 23386 0 23442 800
rect 23662 0 23718 800
rect 23938 0 23994 800
rect 24306 0 24362 800
rect 24582 0 24638 800
rect 24858 0 24914 800
rect 25134 0 25190 800
rect 25410 0 25466 800
rect 25686 0 25742 800
rect 26054 0 26110 800
rect 26330 0 26386 800
rect 26606 0 26662 800
rect 26882 0 26938 800
rect 27158 0 27214 800
rect 27434 0 27490 800
rect 27802 0 27858 800
rect 28078 0 28134 800
rect 28354 0 28410 800
rect 28630 0 28686 800
rect 28906 0 28962 800
rect 29182 0 29238 800
rect 29550 0 29606 800
rect 29826 0 29882 800
rect 30102 0 30158 800
rect 30378 0 30434 800
rect 30654 0 30710 800
rect 31022 0 31078 800
rect 31298 0 31354 800
rect 31574 0 31630 800
rect 31850 0 31906 800
rect 32126 0 32182 800
rect 32402 0 32458 800
rect 32770 0 32826 800
rect 33046 0 33102 800
rect 33322 0 33378 800
rect 33598 0 33654 800
rect 33874 0 33930 800
rect 34150 0 34206 800
rect 34518 0 34574 800
rect 34794 0 34850 800
rect 35070 0 35126 800
rect 35346 0 35402 800
rect 35622 0 35678 800
rect 35898 0 35954 800
rect 36266 0 36322 800
rect 36542 0 36598 800
rect 36818 0 36874 800
rect 37094 0 37150 800
rect 37370 0 37426 800
rect 37646 0 37702 800
rect 38014 0 38070 800
rect 38290 0 38346 800
rect 38566 0 38622 800
rect 38842 0 38898 800
rect 39118 0 39174 800
rect 39394 0 39450 800
rect 39762 0 39818 800
rect 40038 0 40094 800
rect 40314 0 40370 800
rect 40590 0 40646 800
rect 40866 0 40922 800
rect 41142 0 41198 800
rect 41510 0 41566 800
rect 41786 0 41842 800
rect 42062 0 42118 800
rect 42338 0 42394 800
rect 42614 0 42670 800
rect 42890 0 42946 800
rect 43258 0 43314 800
rect 43534 0 43590 800
rect 43810 0 43866 800
rect 44086 0 44142 800
rect 44362 0 44418 800
rect 44638 0 44694 800
rect 45006 0 45062 800
rect 45282 0 45338 800
rect 45558 0 45614 800
rect 45834 0 45890 800
rect 46110 0 46166 800
rect 46478 0 46534 800
rect 46754 0 46810 800
rect 47030 0 47086 800
rect 47306 0 47362 800
rect 47582 0 47638 800
rect 47858 0 47914 800
rect 48226 0 48282 800
rect 48502 0 48558 800
rect 48778 0 48834 800
rect 49054 0 49110 800
rect 49330 0 49386 800
rect 49606 0 49662 800
rect 49974 0 50030 800
rect 50250 0 50306 800
rect 50526 0 50582 800
rect 50802 0 50858 800
rect 51078 0 51134 800
rect 51354 0 51410 800
rect 51722 0 51778 800
rect 51998 0 52054 800
rect 52274 0 52330 800
rect 52550 0 52606 800
rect 52826 0 52882 800
rect 53102 0 53158 800
rect 53470 0 53526 800
rect 53746 0 53802 800
rect 54022 0 54078 800
rect 54298 0 54354 800
rect 54574 0 54630 800
rect 54850 0 54906 800
rect 55218 0 55274 800
rect 55494 0 55550 800
rect 55770 0 55826 800
rect 56046 0 56102 800
rect 56322 0 56378 800
rect 56598 0 56654 800
rect 56966 0 57022 800
rect 57242 0 57298 800
rect 57518 0 57574 800
rect 57794 0 57850 800
rect 58070 0 58126 800
rect 58346 0 58402 800
rect 58714 0 58770 800
rect 58990 0 59046 800
rect 59266 0 59322 800
rect 59542 0 59598 800
rect 59818 0 59874 800
rect 60186 0 60242 800
rect 60462 0 60518 800
rect 60738 0 60794 800
rect 61014 0 61070 800
rect 61290 0 61346 800
rect 61566 0 61622 800
rect 61934 0 61990 800
rect 62210 0 62266 800
rect 62486 0 62542 800
rect 62762 0 62818 800
rect 63038 0 63094 800
rect 63314 0 63370 800
rect 63682 0 63738 800
rect 63958 0 64014 800
rect 64234 0 64290 800
rect 64510 0 64566 800
rect 64786 0 64842 800
rect 65062 0 65118 800
rect 65430 0 65486 800
rect 65706 0 65762 800
rect 65982 0 66038 800
rect 66258 0 66314 800
rect 66534 0 66590 800
rect 66810 0 66866 800
rect 67178 0 67234 800
rect 67454 0 67510 800
rect 67730 0 67786 800
rect 68006 0 68062 800
rect 68282 0 68338 800
rect 68558 0 68614 800
rect 68926 0 68982 800
rect 69202 0 69258 800
rect 69478 0 69534 800
rect 69754 0 69810 800
rect 70030 0 70086 800
rect 70306 0 70362 800
rect 70674 0 70730 800
rect 70950 0 71006 800
rect 71226 0 71282 800
rect 71502 0 71558 800
rect 71778 0 71834 800
rect 72054 0 72110 800
rect 72422 0 72478 800
rect 72698 0 72754 800
rect 72974 0 73030 800
rect 73250 0 73306 800
rect 73526 0 73582 800
rect 73802 0 73858 800
rect 74170 0 74226 800
rect 74446 0 74502 800
rect 74722 0 74778 800
rect 74998 0 75054 800
rect 75274 0 75330 800
rect 75642 0 75698 800
rect 75918 0 75974 800
rect 76194 0 76250 800
rect 76470 0 76526 800
rect 76746 0 76802 800
rect 77022 0 77078 800
rect 77390 0 77446 800
rect 77666 0 77722 800
rect 77942 0 77998 800
rect 78218 0 78274 800
rect 78494 0 78550 800
rect 78770 0 78826 800
rect 79138 0 79194 800
rect 79414 0 79470 800
rect 79690 0 79746 800
rect 79966 0 80022 800
rect 80242 0 80298 800
rect 80518 0 80574 800
rect 80886 0 80942 800
rect 81162 0 81218 800
rect 81438 0 81494 800
rect 81714 0 81770 800
rect 81990 0 82046 800
rect 82266 0 82322 800
rect 82634 0 82690 800
rect 82910 0 82966 800
rect 83186 0 83242 800
rect 83462 0 83518 800
rect 83738 0 83794 800
rect 84014 0 84070 800
rect 84382 0 84438 800
rect 84658 0 84714 800
rect 84934 0 84990 800
rect 85210 0 85266 800
rect 85486 0 85542 800
rect 85762 0 85818 800
rect 86130 0 86186 800
rect 86406 0 86462 800
rect 86682 0 86738 800
rect 86958 0 87014 800
rect 87234 0 87290 800
rect 87510 0 87566 800
rect 87878 0 87934 800
rect 88154 0 88210 800
rect 88430 0 88486 800
rect 88706 0 88762 800
rect 88982 0 89038 800
rect 89258 0 89314 800
rect 89626 0 89682 800
rect 89902 0 89958 800
rect 90178 0 90234 800
rect 90454 0 90510 800
rect 90730 0 90786 800
rect 91098 0 91154 800
rect 91374 0 91430 800
rect 91650 0 91706 800
rect 91926 0 91982 800
rect 92202 0 92258 800
rect 92478 0 92534 800
rect 92846 0 92902 800
rect 93122 0 93178 800
rect 93398 0 93454 800
rect 93674 0 93730 800
rect 93950 0 94006 800
rect 94226 0 94282 800
rect 94594 0 94650 800
rect 94870 0 94926 800
rect 95146 0 95202 800
rect 95422 0 95478 800
rect 95698 0 95754 800
rect 95974 0 96030 800
rect 96342 0 96398 800
rect 96618 0 96674 800
rect 96894 0 96950 800
rect 97170 0 97226 800
rect 97446 0 97502 800
rect 97722 0 97778 800
rect 98090 0 98146 800
rect 98366 0 98422 800
rect 98642 0 98698 800
rect 98918 0 98974 800
rect 99194 0 99250 800
rect 99470 0 99526 800
rect 99838 0 99894 800
rect 100114 0 100170 800
rect 100390 0 100446 800
rect 100666 0 100722 800
rect 100942 0 100998 800
rect 101218 0 101274 800
rect 101586 0 101642 800
rect 101862 0 101918 800
rect 102138 0 102194 800
rect 102414 0 102470 800
rect 102690 0 102746 800
rect 102966 0 103022 800
rect 103334 0 103390 800
rect 103610 0 103666 800
rect 103886 0 103942 800
rect 104162 0 104218 800
rect 104438 0 104494 800
rect 104714 0 104770 800
rect 105082 0 105138 800
rect 105358 0 105414 800
rect 105634 0 105690 800
rect 105910 0 105966 800
rect 106186 0 106242 800
rect 106554 0 106610 800
rect 106830 0 106886 800
rect 107106 0 107162 800
rect 107382 0 107438 800
rect 107658 0 107714 800
rect 107934 0 107990 800
rect 108302 0 108358 800
rect 108578 0 108634 800
rect 108854 0 108910 800
rect 109130 0 109186 800
rect 109406 0 109462 800
rect 109682 0 109738 800
rect 110050 0 110106 800
rect 110326 0 110382 800
rect 110602 0 110658 800
rect 110878 0 110934 800
rect 111154 0 111210 800
rect 111430 0 111486 800
rect 111798 0 111854 800
rect 112074 0 112130 800
rect 112350 0 112406 800
rect 112626 0 112682 800
rect 112902 0 112958 800
rect 113178 0 113234 800
rect 113546 0 113602 800
rect 113822 0 113878 800
rect 114098 0 114154 800
rect 114374 0 114430 800
rect 114650 0 114706 800
rect 114926 0 114982 800
rect 115294 0 115350 800
rect 115570 0 115626 800
rect 115846 0 115902 800
rect 116122 0 116178 800
rect 116398 0 116454 800
rect 116674 0 116730 800
rect 117042 0 117098 800
rect 117318 0 117374 800
rect 117594 0 117650 800
rect 117870 0 117926 800
rect 118146 0 118202 800
rect 118422 0 118478 800
rect 118790 0 118846 800
rect 119066 0 119122 800
rect 119342 0 119398 800
rect 119618 0 119674 800
rect 119894 0 119950 800
rect 120262 0 120318 800
rect 120538 0 120594 800
rect 120814 0 120870 800
rect 121090 0 121146 800
rect 121366 0 121422 800
rect 121642 0 121698 800
rect 122010 0 122066 800
rect 122286 0 122342 800
rect 122562 0 122618 800
rect 122838 0 122894 800
rect 123114 0 123170 800
rect 123390 0 123446 800
rect 123758 0 123814 800
rect 124034 0 124090 800
rect 124310 0 124366 800
rect 124586 0 124642 800
rect 124862 0 124918 800
rect 125138 0 125194 800
rect 125506 0 125562 800
rect 125782 0 125838 800
rect 126058 0 126114 800
rect 126334 0 126390 800
rect 126610 0 126666 800
rect 126886 0 126942 800
rect 127254 0 127310 800
rect 127530 0 127586 800
rect 127806 0 127862 800
rect 128082 0 128138 800
rect 128358 0 128414 800
rect 128634 0 128690 800
rect 129002 0 129058 800
rect 129278 0 129334 800
rect 129554 0 129610 800
rect 129830 0 129886 800
rect 130106 0 130162 800
rect 130382 0 130438 800
rect 130750 0 130806 800
rect 131026 0 131082 800
rect 131302 0 131358 800
rect 131578 0 131634 800
rect 131854 0 131910 800
rect 132130 0 132186 800
rect 132498 0 132554 800
rect 132774 0 132830 800
rect 133050 0 133106 800
rect 133326 0 133382 800
rect 133602 0 133658 800
rect 133878 0 133934 800
rect 134246 0 134302 800
rect 134522 0 134578 800
rect 134798 0 134854 800
rect 135074 0 135130 800
rect 135350 0 135406 800
rect 135718 0 135774 800
rect 135994 0 136050 800
rect 136270 0 136326 800
rect 136546 0 136602 800
rect 136822 0 136878 800
rect 137098 0 137154 800
rect 137466 0 137522 800
rect 137742 0 137798 800
rect 138018 0 138074 800
rect 138294 0 138350 800
rect 138570 0 138626 800
rect 138846 0 138902 800
rect 139214 0 139270 800
rect 139490 0 139546 800
rect 139766 0 139822 800
rect 140042 0 140098 800
rect 140318 0 140374 800
rect 140594 0 140650 800
rect 140962 0 141018 800
rect 141238 0 141294 800
rect 141514 0 141570 800
rect 141790 0 141846 800
rect 142066 0 142122 800
rect 142342 0 142398 800
rect 142710 0 142766 800
rect 142986 0 143042 800
rect 143262 0 143318 800
rect 143538 0 143594 800
rect 143814 0 143870 800
rect 144090 0 144146 800
rect 144458 0 144514 800
rect 144734 0 144790 800
rect 145010 0 145066 800
rect 145286 0 145342 800
rect 145562 0 145618 800
rect 145838 0 145894 800
rect 146206 0 146262 800
rect 146482 0 146538 800
rect 146758 0 146814 800
rect 147034 0 147090 800
rect 147310 0 147366 800
rect 147586 0 147642 800
rect 147954 0 148010 800
rect 148230 0 148286 800
rect 148506 0 148562 800
rect 148782 0 148838 800
rect 149058 0 149114 800
rect 149334 0 149390 800
rect 149702 0 149758 800
rect 149978 0 150034 800
rect 150254 0 150310 800
rect 150530 0 150586 800
rect 150806 0 150862 800
rect 151174 0 151230 800
rect 151450 0 151506 800
rect 151726 0 151782 800
rect 152002 0 152058 800
rect 152278 0 152334 800
rect 152554 0 152610 800
rect 152922 0 152978 800
rect 153198 0 153254 800
rect 153474 0 153530 800
rect 153750 0 153806 800
rect 154026 0 154082 800
rect 154302 0 154358 800
rect 154670 0 154726 800
rect 154946 0 155002 800
rect 155222 0 155278 800
rect 155498 0 155554 800
rect 155774 0 155830 800
rect 156050 0 156106 800
rect 156418 0 156474 800
rect 156694 0 156750 800
rect 156970 0 157026 800
rect 157246 0 157302 800
rect 157522 0 157578 800
rect 157798 0 157854 800
rect 158166 0 158222 800
rect 158442 0 158498 800
rect 158718 0 158774 800
rect 158994 0 159050 800
rect 159270 0 159326 800
rect 159546 0 159602 800
rect 159914 0 159970 800
rect 160190 0 160246 800
rect 160466 0 160522 800
rect 160742 0 160798 800
rect 161018 0 161074 800
rect 161294 0 161350 800
rect 161662 0 161718 800
rect 161938 0 161994 800
rect 162214 0 162270 800
rect 162490 0 162546 800
rect 162766 0 162822 800
rect 163042 0 163098 800
rect 163410 0 163466 800
rect 163686 0 163742 800
rect 163962 0 164018 800
rect 164238 0 164294 800
rect 164514 0 164570 800
<< obsm2 >>
rect 20 166068 422 166124
rect 590 166068 1342 166124
rect 1510 166068 2354 166124
rect 2522 166068 3366 166124
rect 3534 166068 4286 166124
rect 4454 166068 5298 166124
rect 5466 166068 6310 166124
rect 6478 166068 7322 166124
rect 7490 166068 8242 166124
rect 8410 166068 9254 166124
rect 9422 166068 10266 166124
rect 10434 166068 11186 166124
rect 11354 166068 12198 166124
rect 12366 166068 13210 166124
rect 13378 166068 14222 166124
rect 14390 166068 15142 166124
rect 15310 166068 16154 166124
rect 16322 166068 17166 166124
rect 17334 166068 18178 166124
rect 18346 166068 19098 166124
rect 19266 166068 20110 166124
rect 20278 166068 21122 166124
rect 21290 166068 22042 166124
rect 22210 166068 23054 166124
rect 23222 166068 24066 166124
rect 24234 166068 25078 166124
rect 25246 166068 25998 166124
rect 26166 166068 27010 166124
rect 27178 166068 28022 166124
rect 28190 166068 29034 166124
rect 29202 166068 29954 166124
rect 30122 166068 30966 166124
rect 31134 166068 31978 166124
rect 32146 166068 32898 166124
rect 33066 166068 33910 166124
rect 34078 166068 34922 166124
rect 35090 166068 35934 166124
rect 36102 166068 36854 166124
rect 37022 166068 37866 166124
rect 38034 166068 38878 166124
rect 39046 166068 39798 166124
rect 39966 166068 40810 166124
rect 40978 166068 41822 166124
rect 41990 166068 42834 166124
rect 43002 166068 43754 166124
rect 43922 166068 44766 166124
rect 44934 166068 45778 166124
rect 45946 166068 46790 166124
rect 46958 166068 47710 166124
rect 47878 166068 48722 166124
rect 48890 166068 49734 166124
rect 49902 166068 50654 166124
rect 50822 166068 51666 166124
rect 51834 166068 52678 166124
rect 52846 166068 53690 166124
rect 53858 166068 54610 166124
rect 54778 166068 55622 166124
rect 55790 166068 56634 166124
rect 56802 166068 57646 166124
rect 57814 166068 58566 166124
rect 58734 166068 59578 166124
rect 59746 166068 60590 166124
rect 60758 166068 61510 166124
rect 61678 166068 62522 166124
rect 62690 166068 63534 166124
rect 63702 166068 64546 166124
rect 64714 166068 65466 166124
rect 65634 166068 66478 166124
rect 66646 166068 67490 166124
rect 67658 166068 68410 166124
rect 68578 166068 69422 166124
rect 69590 166068 70434 166124
rect 70602 166068 71446 166124
rect 71614 166068 72366 166124
rect 72534 166068 73378 166124
rect 73546 166068 74390 166124
rect 74558 166068 75402 166124
rect 75570 166068 76322 166124
rect 76490 166068 77334 166124
rect 77502 166068 78346 166124
rect 78514 166068 79266 166124
rect 79434 166068 80278 166124
rect 80446 166068 81290 166124
rect 81458 166068 82302 166124
rect 82470 166068 83222 166124
rect 83390 166068 84234 166124
rect 84402 166068 85246 166124
rect 85414 166068 86258 166124
rect 86426 166068 87178 166124
rect 87346 166068 88190 166124
rect 88358 166068 89202 166124
rect 89370 166068 90122 166124
rect 90290 166068 91134 166124
rect 91302 166068 92146 166124
rect 92314 166068 93158 166124
rect 93326 166068 94078 166124
rect 94246 166068 95090 166124
rect 95258 166068 96102 166124
rect 96270 166068 97114 166124
rect 97282 166068 98034 166124
rect 98202 166068 99046 166124
rect 99214 166068 100058 166124
rect 100226 166068 100978 166124
rect 101146 166068 101990 166124
rect 102158 166068 103002 166124
rect 103170 166068 104014 166124
rect 104182 166068 104934 166124
rect 105102 166068 105946 166124
rect 106114 166068 106958 166124
rect 107126 166068 107878 166124
rect 108046 166068 108890 166124
rect 109058 166068 109902 166124
rect 110070 166068 110914 166124
rect 111082 166068 111834 166124
rect 112002 166068 112846 166124
rect 113014 166068 113858 166124
rect 114026 166068 114870 166124
rect 115038 166068 115790 166124
rect 115958 166068 116802 166124
rect 116970 166068 117814 166124
rect 117982 166068 118734 166124
rect 118902 166068 119746 166124
rect 119914 166068 120758 166124
rect 120926 166068 121770 166124
rect 121938 166068 122690 166124
rect 122858 166068 123702 166124
rect 123870 166068 124714 166124
rect 124882 166068 125726 166124
rect 125894 166068 126646 166124
rect 126814 166068 127658 166124
rect 127826 166068 128670 166124
rect 128838 166068 129590 166124
rect 129758 166068 130602 166124
rect 130770 166068 131614 166124
rect 131782 166068 132626 166124
rect 132794 166068 133546 166124
rect 133714 166068 134558 166124
rect 134726 166068 135570 166124
rect 135738 166068 136490 166124
rect 136658 166068 137502 166124
rect 137670 166068 138514 166124
rect 138682 166068 139526 166124
rect 139694 166068 140446 166124
rect 140614 166068 141458 166124
rect 141626 166068 142470 166124
rect 142638 166068 143482 166124
rect 143650 166068 144402 166124
rect 144570 166068 145414 166124
rect 145582 166068 146426 166124
rect 146594 166068 147346 166124
rect 147514 166068 148358 166124
rect 148526 166068 149370 166124
rect 149538 166068 150382 166124
rect 150550 166068 151302 166124
rect 151470 166068 152314 166124
rect 152482 166068 153326 166124
rect 153494 166068 154338 166124
rect 154506 166068 155258 166124
rect 155426 166068 156270 166124
rect 156438 166068 157282 166124
rect 157450 166068 158202 166124
rect 158370 166068 159214 166124
rect 159382 166068 160226 166124
rect 160394 166068 161238 166124
rect 161406 166068 162158 166124
rect 162326 166068 163170 166124
rect 163338 166068 164182 166124
rect 164350 166068 164754 166124
rect 20 856 164754 166068
rect 20 478 54 856
rect 222 478 330 856
rect 498 478 606 856
rect 774 478 882 856
rect 1050 478 1158 856
rect 1326 478 1434 856
rect 1602 478 1802 856
rect 1970 478 2078 856
rect 2246 478 2354 856
rect 2522 478 2630 856
rect 2798 478 2906 856
rect 3074 478 3182 856
rect 3350 478 3550 856
rect 3718 478 3826 856
rect 3994 478 4102 856
rect 4270 478 4378 856
rect 4546 478 4654 856
rect 4822 478 4930 856
rect 5098 478 5298 856
rect 5466 478 5574 856
rect 5742 478 5850 856
rect 6018 478 6126 856
rect 6294 478 6402 856
rect 6570 478 6678 856
rect 6846 478 7046 856
rect 7214 478 7322 856
rect 7490 478 7598 856
rect 7766 478 7874 856
rect 8042 478 8150 856
rect 8318 478 8426 856
rect 8594 478 8794 856
rect 8962 478 9070 856
rect 9238 478 9346 856
rect 9514 478 9622 856
rect 9790 478 9898 856
rect 10066 478 10174 856
rect 10342 478 10542 856
rect 10710 478 10818 856
rect 10986 478 11094 856
rect 11262 478 11370 856
rect 11538 478 11646 856
rect 11814 478 11922 856
rect 12090 478 12290 856
rect 12458 478 12566 856
rect 12734 478 12842 856
rect 13010 478 13118 856
rect 13286 478 13394 856
rect 13562 478 13670 856
rect 13838 478 14038 856
rect 14206 478 14314 856
rect 14482 478 14590 856
rect 14758 478 14866 856
rect 15034 478 15142 856
rect 15310 478 15510 856
rect 15678 478 15786 856
rect 15954 478 16062 856
rect 16230 478 16338 856
rect 16506 478 16614 856
rect 16782 478 16890 856
rect 17058 478 17258 856
rect 17426 478 17534 856
rect 17702 478 17810 856
rect 17978 478 18086 856
rect 18254 478 18362 856
rect 18530 478 18638 856
rect 18806 478 19006 856
rect 19174 478 19282 856
rect 19450 478 19558 856
rect 19726 478 19834 856
rect 20002 478 20110 856
rect 20278 478 20386 856
rect 20554 478 20754 856
rect 20922 478 21030 856
rect 21198 478 21306 856
rect 21474 478 21582 856
rect 21750 478 21858 856
rect 22026 478 22134 856
rect 22302 478 22502 856
rect 22670 478 22778 856
rect 22946 478 23054 856
rect 23222 478 23330 856
rect 23498 478 23606 856
rect 23774 478 23882 856
rect 24050 478 24250 856
rect 24418 478 24526 856
rect 24694 478 24802 856
rect 24970 478 25078 856
rect 25246 478 25354 856
rect 25522 478 25630 856
rect 25798 478 25998 856
rect 26166 478 26274 856
rect 26442 478 26550 856
rect 26718 478 26826 856
rect 26994 478 27102 856
rect 27270 478 27378 856
rect 27546 478 27746 856
rect 27914 478 28022 856
rect 28190 478 28298 856
rect 28466 478 28574 856
rect 28742 478 28850 856
rect 29018 478 29126 856
rect 29294 478 29494 856
rect 29662 478 29770 856
rect 29938 478 30046 856
rect 30214 478 30322 856
rect 30490 478 30598 856
rect 30766 478 30966 856
rect 31134 478 31242 856
rect 31410 478 31518 856
rect 31686 478 31794 856
rect 31962 478 32070 856
rect 32238 478 32346 856
rect 32514 478 32714 856
rect 32882 478 32990 856
rect 33158 478 33266 856
rect 33434 478 33542 856
rect 33710 478 33818 856
rect 33986 478 34094 856
rect 34262 478 34462 856
rect 34630 478 34738 856
rect 34906 478 35014 856
rect 35182 478 35290 856
rect 35458 478 35566 856
rect 35734 478 35842 856
rect 36010 478 36210 856
rect 36378 478 36486 856
rect 36654 478 36762 856
rect 36930 478 37038 856
rect 37206 478 37314 856
rect 37482 478 37590 856
rect 37758 478 37958 856
rect 38126 478 38234 856
rect 38402 478 38510 856
rect 38678 478 38786 856
rect 38954 478 39062 856
rect 39230 478 39338 856
rect 39506 478 39706 856
rect 39874 478 39982 856
rect 40150 478 40258 856
rect 40426 478 40534 856
rect 40702 478 40810 856
rect 40978 478 41086 856
rect 41254 478 41454 856
rect 41622 478 41730 856
rect 41898 478 42006 856
rect 42174 478 42282 856
rect 42450 478 42558 856
rect 42726 478 42834 856
rect 43002 478 43202 856
rect 43370 478 43478 856
rect 43646 478 43754 856
rect 43922 478 44030 856
rect 44198 478 44306 856
rect 44474 478 44582 856
rect 44750 478 44950 856
rect 45118 478 45226 856
rect 45394 478 45502 856
rect 45670 478 45778 856
rect 45946 478 46054 856
rect 46222 478 46422 856
rect 46590 478 46698 856
rect 46866 478 46974 856
rect 47142 478 47250 856
rect 47418 478 47526 856
rect 47694 478 47802 856
rect 47970 478 48170 856
rect 48338 478 48446 856
rect 48614 478 48722 856
rect 48890 478 48998 856
rect 49166 478 49274 856
rect 49442 478 49550 856
rect 49718 478 49918 856
rect 50086 478 50194 856
rect 50362 478 50470 856
rect 50638 478 50746 856
rect 50914 478 51022 856
rect 51190 478 51298 856
rect 51466 478 51666 856
rect 51834 478 51942 856
rect 52110 478 52218 856
rect 52386 478 52494 856
rect 52662 478 52770 856
rect 52938 478 53046 856
rect 53214 478 53414 856
rect 53582 478 53690 856
rect 53858 478 53966 856
rect 54134 478 54242 856
rect 54410 478 54518 856
rect 54686 478 54794 856
rect 54962 478 55162 856
rect 55330 478 55438 856
rect 55606 478 55714 856
rect 55882 478 55990 856
rect 56158 478 56266 856
rect 56434 478 56542 856
rect 56710 478 56910 856
rect 57078 478 57186 856
rect 57354 478 57462 856
rect 57630 478 57738 856
rect 57906 478 58014 856
rect 58182 478 58290 856
rect 58458 478 58658 856
rect 58826 478 58934 856
rect 59102 478 59210 856
rect 59378 478 59486 856
rect 59654 478 59762 856
rect 59930 478 60130 856
rect 60298 478 60406 856
rect 60574 478 60682 856
rect 60850 478 60958 856
rect 61126 478 61234 856
rect 61402 478 61510 856
rect 61678 478 61878 856
rect 62046 478 62154 856
rect 62322 478 62430 856
rect 62598 478 62706 856
rect 62874 478 62982 856
rect 63150 478 63258 856
rect 63426 478 63626 856
rect 63794 478 63902 856
rect 64070 478 64178 856
rect 64346 478 64454 856
rect 64622 478 64730 856
rect 64898 478 65006 856
rect 65174 478 65374 856
rect 65542 478 65650 856
rect 65818 478 65926 856
rect 66094 478 66202 856
rect 66370 478 66478 856
rect 66646 478 66754 856
rect 66922 478 67122 856
rect 67290 478 67398 856
rect 67566 478 67674 856
rect 67842 478 67950 856
rect 68118 478 68226 856
rect 68394 478 68502 856
rect 68670 478 68870 856
rect 69038 478 69146 856
rect 69314 478 69422 856
rect 69590 478 69698 856
rect 69866 478 69974 856
rect 70142 478 70250 856
rect 70418 478 70618 856
rect 70786 478 70894 856
rect 71062 478 71170 856
rect 71338 478 71446 856
rect 71614 478 71722 856
rect 71890 478 71998 856
rect 72166 478 72366 856
rect 72534 478 72642 856
rect 72810 478 72918 856
rect 73086 478 73194 856
rect 73362 478 73470 856
rect 73638 478 73746 856
rect 73914 478 74114 856
rect 74282 478 74390 856
rect 74558 478 74666 856
rect 74834 478 74942 856
rect 75110 478 75218 856
rect 75386 478 75586 856
rect 75754 478 75862 856
rect 76030 478 76138 856
rect 76306 478 76414 856
rect 76582 478 76690 856
rect 76858 478 76966 856
rect 77134 478 77334 856
rect 77502 478 77610 856
rect 77778 478 77886 856
rect 78054 478 78162 856
rect 78330 478 78438 856
rect 78606 478 78714 856
rect 78882 478 79082 856
rect 79250 478 79358 856
rect 79526 478 79634 856
rect 79802 478 79910 856
rect 80078 478 80186 856
rect 80354 478 80462 856
rect 80630 478 80830 856
rect 80998 478 81106 856
rect 81274 478 81382 856
rect 81550 478 81658 856
rect 81826 478 81934 856
rect 82102 478 82210 856
rect 82378 478 82578 856
rect 82746 478 82854 856
rect 83022 478 83130 856
rect 83298 478 83406 856
rect 83574 478 83682 856
rect 83850 478 83958 856
rect 84126 478 84326 856
rect 84494 478 84602 856
rect 84770 478 84878 856
rect 85046 478 85154 856
rect 85322 478 85430 856
rect 85598 478 85706 856
rect 85874 478 86074 856
rect 86242 478 86350 856
rect 86518 478 86626 856
rect 86794 478 86902 856
rect 87070 478 87178 856
rect 87346 478 87454 856
rect 87622 478 87822 856
rect 87990 478 88098 856
rect 88266 478 88374 856
rect 88542 478 88650 856
rect 88818 478 88926 856
rect 89094 478 89202 856
rect 89370 478 89570 856
rect 89738 478 89846 856
rect 90014 478 90122 856
rect 90290 478 90398 856
rect 90566 478 90674 856
rect 90842 478 91042 856
rect 91210 478 91318 856
rect 91486 478 91594 856
rect 91762 478 91870 856
rect 92038 478 92146 856
rect 92314 478 92422 856
rect 92590 478 92790 856
rect 92958 478 93066 856
rect 93234 478 93342 856
rect 93510 478 93618 856
rect 93786 478 93894 856
rect 94062 478 94170 856
rect 94338 478 94538 856
rect 94706 478 94814 856
rect 94982 478 95090 856
rect 95258 478 95366 856
rect 95534 478 95642 856
rect 95810 478 95918 856
rect 96086 478 96286 856
rect 96454 478 96562 856
rect 96730 478 96838 856
rect 97006 478 97114 856
rect 97282 478 97390 856
rect 97558 478 97666 856
rect 97834 478 98034 856
rect 98202 478 98310 856
rect 98478 478 98586 856
rect 98754 478 98862 856
rect 99030 478 99138 856
rect 99306 478 99414 856
rect 99582 478 99782 856
rect 99950 478 100058 856
rect 100226 478 100334 856
rect 100502 478 100610 856
rect 100778 478 100886 856
rect 101054 478 101162 856
rect 101330 478 101530 856
rect 101698 478 101806 856
rect 101974 478 102082 856
rect 102250 478 102358 856
rect 102526 478 102634 856
rect 102802 478 102910 856
rect 103078 478 103278 856
rect 103446 478 103554 856
rect 103722 478 103830 856
rect 103998 478 104106 856
rect 104274 478 104382 856
rect 104550 478 104658 856
rect 104826 478 105026 856
rect 105194 478 105302 856
rect 105470 478 105578 856
rect 105746 478 105854 856
rect 106022 478 106130 856
rect 106298 478 106498 856
rect 106666 478 106774 856
rect 106942 478 107050 856
rect 107218 478 107326 856
rect 107494 478 107602 856
rect 107770 478 107878 856
rect 108046 478 108246 856
rect 108414 478 108522 856
rect 108690 478 108798 856
rect 108966 478 109074 856
rect 109242 478 109350 856
rect 109518 478 109626 856
rect 109794 478 109994 856
rect 110162 478 110270 856
rect 110438 478 110546 856
rect 110714 478 110822 856
rect 110990 478 111098 856
rect 111266 478 111374 856
rect 111542 478 111742 856
rect 111910 478 112018 856
rect 112186 478 112294 856
rect 112462 478 112570 856
rect 112738 478 112846 856
rect 113014 478 113122 856
rect 113290 478 113490 856
rect 113658 478 113766 856
rect 113934 478 114042 856
rect 114210 478 114318 856
rect 114486 478 114594 856
rect 114762 478 114870 856
rect 115038 478 115238 856
rect 115406 478 115514 856
rect 115682 478 115790 856
rect 115958 478 116066 856
rect 116234 478 116342 856
rect 116510 478 116618 856
rect 116786 478 116986 856
rect 117154 478 117262 856
rect 117430 478 117538 856
rect 117706 478 117814 856
rect 117982 478 118090 856
rect 118258 478 118366 856
rect 118534 478 118734 856
rect 118902 478 119010 856
rect 119178 478 119286 856
rect 119454 478 119562 856
rect 119730 478 119838 856
rect 120006 478 120206 856
rect 120374 478 120482 856
rect 120650 478 120758 856
rect 120926 478 121034 856
rect 121202 478 121310 856
rect 121478 478 121586 856
rect 121754 478 121954 856
rect 122122 478 122230 856
rect 122398 478 122506 856
rect 122674 478 122782 856
rect 122950 478 123058 856
rect 123226 478 123334 856
rect 123502 478 123702 856
rect 123870 478 123978 856
rect 124146 478 124254 856
rect 124422 478 124530 856
rect 124698 478 124806 856
rect 124974 478 125082 856
rect 125250 478 125450 856
rect 125618 478 125726 856
rect 125894 478 126002 856
rect 126170 478 126278 856
rect 126446 478 126554 856
rect 126722 478 126830 856
rect 126998 478 127198 856
rect 127366 478 127474 856
rect 127642 478 127750 856
rect 127918 478 128026 856
rect 128194 478 128302 856
rect 128470 478 128578 856
rect 128746 478 128946 856
rect 129114 478 129222 856
rect 129390 478 129498 856
rect 129666 478 129774 856
rect 129942 478 130050 856
rect 130218 478 130326 856
rect 130494 478 130694 856
rect 130862 478 130970 856
rect 131138 478 131246 856
rect 131414 478 131522 856
rect 131690 478 131798 856
rect 131966 478 132074 856
rect 132242 478 132442 856
rect 132610 478 132718 856
rect 132886 478 132994 856
rect 133162 478 133270 856
rect 133438 478 133546 856
rect 133714 478 133822 856
rect 133990 478 134190 856
rect 134358 478 134466 856
rect 134634 478 134742 856
rect 134910 478 135018 856
rect 135186 478 135294 856
rect 135462 478 135662 856
rect 135830 478 135938 856
rect 136106 478 136214 856
rect 136382 478 136490 856
rect 136658 478 136766 856
rect 136934 478 137042 856
rect 137210 478 137410 856
rect 137578 478 137686 856
rect 137854 478 137962 856
rect 138130 478 138238 856
rect 138406 478 138514 856
rect 138682 478 138790 856
rect 138958 478 139158 856
rect 139326 478 139434 856
rect 139602 478 139710 856
rect 139878 478 139986 856
rect 140154 478 140262 856
rect 140430 478 140538 856
rect 140706 478 140906 856
rect 141074 478 141182 856
rect 141350 478 141458 856
rect 141626 478 141734 856
rect 141902 478 142010 856
rect 142178 478 142286 856
rect 142454 478 142654 856
rect 142822 478 142930 856
rect 143098 478 143206 856
rect 143374 478 143482 856
rect 143650 478 143758 856
rect 143926 478 144034 856
rect 144202 478 144402 856
rect 144570 478 144678 856
rect 144846 478 144954 856
rect 145122 478 145230 856
rect 145398 478 145506 856
rect 145674 478 145782 856
rect 145950 478 146150 856
rect 146318 478 146426 856
rect 146594 478 146702 856
rect 146870 478 146978 856
rect 147146 478 147254 856
rect 147422 478 147530 856
rect 147698 478 147898 856
rect 148066 478 148174 856
rect 148342 478 148450 856
rect 148618 478 148726 856
rect 148894 478 149002 856
rect 149170 478 149278 856
rect 149446 478 149646 856
rect 149814 478 149922 856
rect 150090 478 150198 856
rect 150366 478 150474 856
rect 150642 478 150750 856
rect 150918 478 151118 856
rect 151286 478 151394 856
rect 151562 478 151670 856
rect 151838 478 151946 856
rect 152114 478 152222 856
rect 152390 478 152498 856
rect 152666 478 152866 856
rect 153034 478 153142 856
rect 153310 478 153418 856
rect 153586 478 153694 856
rect 153862 478 153970 856
rect 154138 478 154246 856
rect 154414 478 154614 856
rect 154782 478 154890 856
rect 155058 478 155166 856
rect 155334 478 155442 856
rect 155610 478 155718 856
rect 155886 478 155994 856
rect 156162 478 156362 856
rect 156530 478 156638 856
rect 156806 478 156914 856
rect 157082 478 157190 856
rect 157358 478 157466 856
rect 157634 478 157742 856
rect 157910 478 158110 856
rect 158278 478 158386 856
rect 158554 478 158662 856
rect 158830 478 158938 856
rect 159106 478 159214 856
rect 159382 478 159490 856
rect 159658 478 159858 856
rect 160026 478 160134 856
rect 160302 478 160410 856
rect 160578 478 160686 856
rect 160854 478 160962 856
rect 161130 478 161238 856
rect 161406 478 161606 856
rect 161774 478 161882 856
rect 162050 478 162158 856
rect 162326 478 162434 856
rect 162602 478 162710 856
rect 162878 478 162986 856
rect 163154 478 163354 856
rect 163522 478 163630 856
rect 163798 478 163906 856
rect 164074 478 164182 856
rect 164350 478 164458 856
rect 164626 478 164754 856
<< metal3 >>
rect 0 165248 800 165368
rect 163980 165384 164780 165504
rect 163980 162664 164780 162784
rect 0 162256 800 162376
rect 163980 159944 164780 160064
rect 0 159264 800 159384
rect 163980 157224 164780 157344
rect 0 156272 800 156392
rect 163980 154504 164780 154624
rect 0 153280 800 153400
rect 163980 151784 164780 151904
rect 0 150288 800 150408
rect 163980 149064 164780 149184
rect 0 147296 800 147416
rect 163980 146344 164780 146464
rect 0 144304 800 144424
rect 163980 143488 164780 143608
rect 0 141312 800 141432
rect 163980 140768 164780 140888
rect 0 138320 800 138440
rect 163980 138048 164780 138168
rect 0 135328 800 135448
rect 163980 135328 164780 135448
rect 0 132472 800 132592
rect 163980 132608 164780 132728
rect 163980 129888 164780 130008
rect 0 129480 800 129600
rect 163980 127168 164780 127288
rect 0 126488 800 126608
rect 163980 124448 164780 124568
rect 0 123496 800 123616
rect 163980 121728 164780 121848
rect 0 120504 800 120624
rect 163980 118872 164780 118992
rect 0 117512 800 117632
rect 163980 116152 164780 116272
rect 0 114520 800 114640
rect 163980 113432 164780 113552
rect 0 111528 800 111648
rect 163980 110712 164780 110832
rect 0 108536 800 108656
rect 163980 107992 164780 108112
rect 0 105544 800 105664
rect 163980 105272 164780 105392
rect 0 102552 800 102672
rect 163980 102552 164780 102672
rect 0 99696 800 99816
rect 163980 99832 164780 99952
rect 163980 97112 164780 97232
rect 0 96704 800 96824
rect 163980 94256 164780 94376
rect 0 93712 800 93832
rect 163980 91536 164780 91656
rect 0 90720 800 90840
rect 163980 88816 164780 88936
rect 0 87728 800 87848
rect 163980 86096 164780 86216
rect 0 84736 800 84856
rect 163980 83376 164780 83496
rect 0 81744 800 81864
rect 163980 80656 164780 80776
rect 0 78752 800 78872
rect 163980 77936 164780 78056
rect 0 75760 800 75880
rect 163980 75216 164780 75336
rect 0 72768 800 72888
rect 163980 72360 164780 72480
rect 0 69776 800 69896
rect 163980 69640 164780 69760
rect 0 66920 800 67040
rect 163980 66920 164780 67040
rect 163980 64200 164780 64320
rect 0 63928 800 64048
rect 163980 61480 164780 61600
rect 0 60936 800 61056
rect 163980 58760 164780 58880
rect 0 57944 800 58064
rect 163980 56040 164780 56160
rect 0 54952 800 55072
rect 163980 53320 164780 53440
rect 0 51960 800 52080
rect 163980 50600 164780 50720
rect 0 48968 800 49088
rect 163980 47744 164780 47864
rect 0 45976 800 46096
rect 163980 45024 164780 45144
rect 0 42984 800 43104
rect 163980 42304 164780 42424
rect 0 39992 800 40112
rect 163980 39584 164780 39704
rect 0 37000 800 37120
rect 163980 36864 164780 36984
rect 0 34144 800 34264
rect 163980 34144 164780 34264
rect 163980 31424 164780 31544
rect 0 31152 800 31272
rect 163980 28704 164780 28824
rect 0 28160 800 28280
rect 163980 25984 164780 26104
rect 0 25168 800 25288
rect 163980 23128 164780 23248
rect 0 22176 800 22296
rect 163980 20408 164780 20528
rect 0 19184 800 19304
rect 163980 17688 164780 17808
rect 0 16192 800 16312
rect 163980 14968 164780 15088
rect 0 13200 800 13320
rect 163980 12248 164780 12368
rect 0 10208 800 10328
rect 163980 9528 164780 9648
rect 0 7216 800 7336
rect 163980 6808 164780 6928
rect 0 4224 800 4344
rect 163980 4088 164780 4208
rect 0 1368 800 1488
rect 163980 1368 164780 1488
<< obsm3 >>
rect 800 165448 163900 165477
rect 880 165304 163900 165448
rect 880 165168 164759 165304
rect 800 162864 164759 165168
rect 800 162584 163900 162864
rect 800 162456 164759 162584
rect 880 162176 164759 162456
rect 800 160144 164759 162176
rect 800 159864 163900 160144
rect 800 159464 164759 159864
rect 880 159184 164759 159464
rect 800 157424 164759 159184
rect 800 157144 163900 157424
rect 800 156472 164759 157144
rect 880 156192 164759 156472
rect 800 154704 164759 156192
rect 800 154424 163900 154704
rect 800 153480 164759 154424
rect 880 153200 164759 153480
rect 800 151984 164759 153200
rect 800 151704 163900 151984
rect 800 150488 164759 151704
rect 880 150208 164759 150488
rect 800 149264 164759 150208
rect 800 148984 163900 149264
rect 800 147496 164759 148984
rect 880 147216 164759 147496
rect 800 146544 164759 147216
rect 800 146264 163900 146544
rect 800 144504 164759 146264
rect 880 144224 164759 144504
rect 800 143688 164759 144224
rect 800 143408 163900 143688
rect 800 141512 164759 143408
rect 880 141232 164759 141512
rect 800 140968 164759 141232
rect 800 140688 163900 140968
rect 800 138520 164759 140688
rect 880 138248 164759 138520
rect 880 138240 163900 138248
rect 800 137968 163900 138240
rect 800 135528 164759 137968
rect 880 135248 163900 135528
rect 800 132808 164759 135248
rect 800 132672 163900 132808
rect 880 132528 163900 132672
rect 880 132392 164759 132528
rect 800 130088 164759 132392
rect 800 129808 163900 130088
rect 800 129680 164759 129808
rect 880 129400 164759 129680
rect 800 127368 164759 129400
rect 800 127088 163900 127368
rect 800 126688 164759 127088
rect 880 126408 164759 126688
rect 800 124648 164759 126408
rect 800 124368 163900 124648
rect 800 123696 164759 124368
rect 880 123416 164759 123696
rect 800 121928 164759 123416
rect 800 121648 163900 121928
rect 800 120704 164759 121648
rect 880 120424 164759 120704
rect 800 119072 164759 120424
rect 800 118792 163900 119072
rect 800 117712 164759 118792
rect 880 117432 164759 117712
rect 800 116352 164759 117432
rect 800 116072 163900 116352
rect 800 114720 164759 116072
rect 880 114440 164759 114720
rect 800 113632 164759 114440
rect 800 113352 163900 113632
rect 800 111728 164759 113352
rect 880 111448 164759 111728
rect 800 110912 164759 111448
rect 800 110632 163900 110912
rect 800 108736 164759 110632
rect 880 108456 164759 108736
rect 800 108192 164759 108456
rect 800 107912 163900 108192
rect 800 105744 164759 107912
rect 880 105472 164759 105744
rect 880 105464 163900 105472
rect 800 105192 163900 105464
rect 800 102752 164759 105192
rect 880 102472 163900 102752
rect 800 100032 164759 102472
rect 800 99896 163900 100032
rect 880 99752 163900 99896
rect 880 99616 164759 99752
rect 800 97312 164759 99616
rect 800 97032 163900 97312
rect 800 96904 164759 97032
rect 880 96624 164759 96904
rect 800 94456 164759 96624
rect 800 94176 163900 94456
rect 800 93912 164759 94176
rect 880 93632 164759 93912
rect 800 91736 164759 93632
rect 800 91456 163900 91736
rect 800 90920 164759 91456
rect 880 90640 164759 90920
rect 800 89016 164759 90640
rect 800 88736 163900 89016
rect 800 87928 164759 88736
rect 880 87648 164759 87928
rect 800 86296 164759 87648
rect 800 86016 163900 86296
rect 800 84936 164759 86016
rect 880 84656 164759 84936
rect 800 83576 164759 84656
rect 800 83296 163900 83576
rect 800 81944 164759 83296
rect 880 81664 164759 81944
rect 800 80856 164759 81664
rect 800 80576 163900 80856
rect 800 78952 164759 80576
rect 880 78672 164759 78952
rect 800 78136 164759 78672
rect 800 77856 163900 78136
rect 800 75960 164759 77856
rect 880 75680 164759 75960
rect 800 75416 164759 75680
rect 800 75136 163900 75416
rect 800 72968 164759 75136
rect 880 72688 164759 72968
rect 800 72560 164759 72688
rect 800 72280 163900 72560
rect 800 69976 164759 72280
rect 880 69840 164759 69976
rect 880 69696 163900 69840
rect 800 69560 163900 69696
rect 800 67120 164759 69560
rect 880 66840 163900 67120
rect 800 64400 164759 66840
rect 800 64128 163900 64400
rect 880 64120 163900 64128
rect 880 63848 164759 64120
rect 800 61680 164759 63848
rect 800 61400 163900 61680
rect 800 61136 164759 61400
rect 880 60856 164759 61136
rect 800 58960 164759 60856
rect 800 58680 163900 58960
rect 800 58144 164759 58680
rect 880 57864 164759 58144
rect 800 56240 164759 57864
rect 800 55960 163900 56240
rect 800 55152 164759 55960
rect 880 54872 164759 55152
rect 800 53520 164759 54872
rect 800 53240 163900 53520
rect 800 52160 164759 53240
rect 880 51880 164759 52160
rect 800 50800 164759 51880
rect 800 50520 163900 50800
rect 800 49168 164759 50520
rect 880 48888 164759 49168
rect 800 47944 164759 48888
rect 800 47664 163900 47944
rect 800 46176 164759 47664
rect 880 45896 164759 46176
rect 800 45224 164759 45896
rect 800 44944 163900 45224
rect 800 43184 164759 44944
rect 880 42904 164759 43184
rect 800 42504 164759 42904
rect 800 42224 163900 42504
rect 800 40192 164759 42224
rect 880 39912 164759 40192
rect 800 39784 164759 39912
rect 800 39504 163900 39784
rect 800 37200 164759 39504
rect 880 37064 164759 37200
rect 880 36920 163900 37064
rect 800 36784 163900 36920
rect 800 34344 164759 36784
rect 880 34064 163900 34344
rect 800 31624 164759 34064
rect 800 31352 163900 31624
rect 880 31344 163900 31352
rect 880 31072 164759 31344
rect 800 28904 164759 31072
rect 800 28624 163900 28904
rect 800 28360 164759 28624
rect 880 28080 164759 28360
rect 800 26184 164759 28080
rect 800 25904 163900 26184
rect 800 25368 164759 25904
rect 880 25088 164759 25368
rect 800 23328 164759 25088
rect 800 23048 163900 23328
rect 800 22376 164759 23048
rect 880 22096 164759 22376
rect 800 20608 164759 22096
rect 800 20328 163900 20608
rect 800 19384 164759 20328
rect 880 19104 164759 19384
rect 800 17888 164759 19104
rect 800 17608 163900 17888
rect 800 16392 164759 17608
rect 880 16112 164759 16392
rect 800 15168 164759 16112
rect 800 14888 163900 15168
rect 800 13400 164759 14888
rect 880 13120 164759 13400
rect 800 12448 164759 13120
rect 800 12168 163900 12448
rect 800 10408 164759 12168
rect 880 10128 164759 10408
rect 800 9728 164759 10128
rect 800 9448 163900 9728
rect 800 7416 164759 9448
rect 880 7136 164759 7416
rect 800 7008 164759 7136
rect 800 6728 163900 7008
rect 800 4424 164759 6728
rect 880 4288 164759 4424
rect 880 4144 163900 4288
rect 800 4008 163900 4144
rect 800 1568 164759 4008
rect 880 1288 163900 1568
rect 800 444 164759 1288
<< metal4 >>
rect 4208 2128 4528 164336
rect 19568 2128 19888 164336
rect 34928 2128 35248 164336
rect 50288 2128 50608 164336
rect 65648 2128 65968 164336
rect 81008 2128 81328 164336
rect 96368 2128 96688 164336
rect 111728 2128 112048 164336
rect 127088 2128 127408 164336
rect 142448 2128 142768 164336
rect 157808 2128 158128 164336
<< obsm4 >>
rect 3187 2048 4128 164117
rect 4608 2048 19488 164117
rect 19968 2048 34848 164117
rect 35328 2048 50208 164117
rect 50688 2048 65568 164117
rect 66048 2048 80928 164117
rect 81408 2048 96288 164117
rect 96768 2048 111648 164117
rect 112128 2048 127008 164117
rect 127488 2048 142368 164117
rect 142848 2048 157728 164117
rect 158208 2048 163149 164117
rect 3187 443 163149 2048
<< labels >>
rlabel metal3 s 163980 4088 164780 4208 6 i_dout0[0]
port 1 nsew signal input
rlabel metal2 s 134614 166124 134670 166924 6 i_dout0[10]
port 2 nsew signal input
rlabel metal3 s 163980 72360 164780 72480 6 i_dout0[11]
port 3 nsew signal input
rlabel metal3 s 0 87728 800 87848 6 i_dout0[12]
port 4 nsew signal input
rlabel metal3 s 163980 83376 164780 83496 6 i_dout0[13]
port 5 nsew signal input
rlabel metal3 s 163980 88816 164780 88936 6 i_dout0[14]
port 6 nsew signal input
rlabel metal2 s 142526 166124 142582 166924 6 i_dout0[15]
port 7 nsew signal input
rlabel metal2 s 146482 166124 146538 166924 6 i_dout0[16]
port 8 nsew signal input
rlabel metal3 s 163980 97112 164780 97232 6 i_dout0[17]
port 9 nsew signal input
rlabel metal2 s 148414 166124 148470 166924 6 i_dout0[18]
port 10 nsew signal input
rlabel metal3 s 163980 102552 164780 102672 6 i_dout0[19]
port 11 nsew signal input
rlabel metal3 s 0 13200 800 13320 6 i_dout0[1]
port 12 nsew signal input
rlabel metal3 s 163980 105272 164780 105392 6 i_dout0[20]
port 13 nsew signal input
rlabel metal3 s 0 117512 800 117632 6 i_dout0[21]
port 14 nsew signal input
rlabel metal2 s 154394 166124 154450 166924 6 i_dout0[22]
port 15 nsew signal input
rlabel metal2 s 161294 0 161350 800 6 i_dout0[23]
port 16 nsew signal input
rlabel metal3 s 0 129480 800 129600 6 i_dout0[24]
port 17 nsew signal input
rlabel metal3 s 0 135328 800 135448 6 i_dout0[25]
port 18 nsew signal input
rlabel metal2 s 163042 0 163098 800 6 i_dout0[26]
port 19 nsew signal input
rlabel metal3 s 0 147296 800 147416 6 i_dout0[27]
port 20 nsew signal input
rlabel metal2 s 163686 0 163742 800 6 i_dout0[28]
port 21 nsew signal input
rlabel metal3 s 163980 149064 164780 149184 6 i_dout0[29]
port 22 nsew signal input
rlabel metal3 s 163980 17688 164780 17808 6 i_dout0[2]
port 23 nsew signal input
rlabel metal2 s 164238 0 164294 800 6 i_dout0[30]
port 24 nsew signal input
rlabel metal3 s 163980 159944 164780 160064 6 i_dout0[31]
port 25 nsew signal input
rlabel metal3 s 163980 28704 164780 28824 6 i_dout0[3]
port 26 nsew signal input
rlabel metal3 s 0 42984 800 43104 6 i_dout0[4]
port 27 nsew signal input
rlabel metal2 s 149702 0 149758 800 6 i_dout0[5]
port 28 nsew signal input
rlabel metal2 s 151174 0 151230 800 6 i_dout0[6]
port 29 nsew signal input
rlabel metal2 s 152278 0 152334 800 6 i_dout0[7]
port 30 nsew signal input
rlabel metal2 s 153474 0 153530 800 6 i_dout0[8]
port 31 nsew signal input
rlabel metal2 s 132682 166124 132738 166924 6 i_dout0[9]
port 32 nsew signal input
rlabel metal2 s 144458 0 144514 800 6 i_dout0_1[0]
port 33 nsew signal input
rlabel metal3 s 163980 64200 164780 64320 6 i_dout0_1[10]
port 34 nsew signal input
rlabel metal2 s 136546 166124 136602 166924 6 i_dout0_1[11]
port 35 nsew signal input
rlabel metal2 s 155498 0 155554 800 6 i_dout0_1[12]
port 36 nsew signal input
rlabel metal3 s 0 90720 800 90840 6 i_dout0_1[13]
port 37 nsew signal input
rlabel metal2 s 139582 166124 139638 166924 6 i_dout0_1[14]
port 38 nsew signal input
rlabel metal2 s 141514 166124 141570 166924 6 i_dout0_1[15]
port 39 nsew signal input
rlabel metal2 s 145470 166124 145526 166924 6 i_dout0_1[16]
port 40 nsew signal input
rlabel metal3 s 0 99696 800 99816 6 i_dout0_1[17]
port 41 nsew signal input
rlabel metal3 s 163980 99832 164780 99952 6 i_dout0_1[18]
port 42 nsew signal input
rlabel metal3 s 0 108536 800 108656 6 i_dout0_1[19]
port 43 nsew signal input
rlabel metal3 s 163980 12248 164780 12368 6 i_dout0_1[1]
port 44 nsew signal input
rlabel metal2 s 159914 0 159970 800 6 i_dout0_1[20]
port 45 nsew signal input
rlabel metal2 s 153382 166124 153438 166924 6 i_dout0_1[21]
port 46 nsew signal input
rlabel metal2 s 160742 0 160798 800 6 i_dout0_1[22]
port 47 nsew signal input
rlabel metal3 s 0 123496 800 123616 6 i_dout0_1[23]
port 48 nsew signal input
rlabel metal2 s 162214 0 162270 800 6 i_dout0_1[24]
port 49 nsew signal input
rlabel metal2 s 157338 166124 157394 166924 6 i_dout0_1[25]
port 50 nsew signal input
rlabel metal2 s 158258 166124 158314 166924 6 i_dout0_1[26]
port 51 nsew signal input
rlabel metal2 s 159270 166124 159326 166924 6 i_dout0_1[27]
port 52 nsew signal input
rlabel metal2 s 161294 166124 161350 166924 6 i_dout0_1[28]
port 53 nsew signal input
rlabel metal3 s 163980 146344 164780 146464 6 i_dout0_1[29]
port 54 nsew signal input
rlabel metal2 s 117870 166124 117926 166924 6 i_dout0_1[2]
port 55 nsew signal input
rlabel metal2 s 163962 0 164018 800 6 i_dout0_1[30]
port 56 nsew signal input
rlabel metal3 s 0 162256 800 162376 6 i_dout0_1[31]
port 57 nsew signal input
rlabel metal3 s 163980 25984 164780 26104 6 i_dout0_1[3]
port 58 nsew signal input
rlabel metal2 s 148782 0 148838 800 6 i_dout0_1[4]
port 59 nsew signal input
rlabel metal3 s 163980 45024 164780 45144 6 i_dout0_1[5]
port 60 nsew signal input
rlabel metal2 s 125782 166124 125838 166924 6 i_dout0_1[6]
port 61 nsew signal input
rlabel metal2 s 152002 0 152058 800 6 i_dout0_1[7]
port 62 nsew signal input
rlabel metal2 s 153198 0 153254 800 6 i_dout0_1[8]
port 63 nsew signal input
rlabel metal3 s 163980 61480 164780 61600 6 i_dout0_1[9]
port 64 nsew signal input
rlabel metal2 s 144734 0 144790 800 6 i_dout1[0]
port 65 nsew signal input
rlabel metal3 s 163980 66920 164780 67040 6 i_dout1[10]
port 66 nsew signal input
rlabel metal3 s 163980 75216 164780 75336 6 i_dout1[11]
port 67 nsew signal input
rlabel metal3 s 163980 77936 164780 78056 6 i_dout1[12]
port 68 nsew signal input
rlabel metal2 s 156050 0 156106 800 6 i_dout1[13]
port 69 nsew signal input
rlabel metal3 s 163980 91536 164780 91656 6 i_dout1[14]
port 70 nsew signal input
rlabel metal2 s 143538 166124 143594 166924 6 i_dout1[15]
port 71 nsew signal input
rlabel metal2 s 157246 0 157302 800 6 i_dout1[16]
port 72 nsew signal input
rlabel metal3 s 0 102552 800 102672 6 i_dout1[17]
port 73 nsew signal input
rlabel metal2 s 158994 0 159050 800 6 i_dout1[18]
port 74 nsew signal input
rlabel metal2 s 150438 166124 150494 166924 6 i_dout1[19]
port 75 nsew signal input
rlabel metal3 s 163980 14968 164780 15088 6 i_dout1[1]
port 76 nsew signal input
rlabel metal3 s 163980 107992 164780 108112 6 i_dout1[20]
port 77 nsew signal input
rlabel metal2 s 160466 0 160522 800 6 i_dout1[21]
port 78 nsew signal input
rlabel metal3 s 163980 116152 164780 116272 6 i_dout1[22]
port 79 nsew signal input
rlabel metal3 s 0 126488 800 126608 6 i_dout1[23]
port 80 nsew signal input
rlabel metal2 s 162490 0 162546 800 6 i_dout1[24]
port 81 nsew signal input
rlabel metal3 s 163980 127168 164780 127288 6 i_dout1[25]
port 82 nsew signal input
rlabel metal2 s 163410 0 163466 800 6 i_dout1[26]
port 83 nsew signal input
rlabel metal3 s 0 150288 800 150408 6 i_dout1[27]
port 84 nsew signal input
rlabel metal3 s 163980 140768 164780 140888 6 i_dout1[28]
port 85 nsew signal input
rlabel metal3 s 0 153280 800 153400 6 i_dout1[29]
port 86 nsew signal input
rlabel metal3 s 0 19184 800 19304 6 i_dout1[2]
port 87 nsew signal input
rlabel metal3 s 0 156272 800 156392 6 i_dout1[30]
port 88 nsew signal input
rlabel metal3 s 163980 162664 164780 162784 6 i_dout1[31]
port 89 nsew signal input
rlabel metal2 s 119802 166124 119858 166924 6 i_dout1[3]
port 90 nsew signal input
rlabel metal2 s 123758 166124 123814 166924 6 i_dout1[4]
port 91 nsew signal input
rlabel metal2 s 149978 0 150034 800 6 i_dout1[5]
port 92 nsew signal input
rlabel metal2 s 151450 0 151506 800 6 i_dout1[6]
port 93 nsew signal input
rlabel metal3 s 163980 53320 164780 53440 6 i_dout1[7]
port 94 nsew signal input
rlabel metal2 s 153750 0 153806 800 6 i_dout1[8]
port 95 nsew signal input
rlabel metal3 s 0 75760 800 75880 6 i_dout1[9]
port 96 nsew signal input
rlabel metal3 s 163980 6808 164780 6928 6 i_dout1_1[0]
port 97 nsew signal input
rlabel metal2 s 154946 0 155002 800 6 i_dout1_1[10]
port 98 nsew signal input
rlabel metal3 s 0 81744 800 81864 6 i_dout1_1[11]
port 99 nsew signal input
rlabel metal3 s 0 84736 800 84856 6 i_dout1_1[12]
port 100 nsew signal input
rlabel metal2 s 155774 0 155830 800 6 i_dout1_1[13]
port 101 nsew signal input
rlabel metal3 s 163980 86096 164780 86216 6 i_dout1_1[14]
port 102 nsew signal input
rlabel metal2 s 156970 0 157026 800 6 i_dout1_1[15]
port 103 nsew signal input
rlabel metal3 s 163980 94256 164780 94376 6 i_dout1_1[16]
port 104 nsew signal input
rlabel metal2 s 158166 0 158222 800 6 i_dout1_1[17]
port 105 nsew signal input
rlabel metal2 s 158718 0 158774 800 6 i_dout1_1[18]
port 106 nsew signal input
rlabel metal2 s 159270 0 159326 800 6 i_dout1_1[19]
port 107 nsew signal input
rlabel metal2 s 145838 0 145894 800 6 i_dout1_1[1]
port 108 nsew signal input
rlabel metal2 s 160190 0 160246 800 6 i_dout1_1[20]
port 109 nsew signal input
rlabel metal3 s 0 114520 800 114640 6 i_dout1_1[21]
port 110 nsew signal input
rlabel metal3 s 0 120504 800 120624 6 i_dout1_1[22]
port 111 nsew signal input
rlabel metal3 s 163980 121728 164780 121848 6 i_dout1_1[23]
port 112 nsew signal input
rlabel metal2 s 155314 166124 155370 166924 6 i_dout1_1[24]
port 113 nsew signal input
rlabel metal3 s 0 132472 800 132592 6 i_dout1_1[25]
port 114 nsew signal input
rlabel metal3 s 163980 132608 164780 132728 6 i_dout1_1[26]
port 115 nsew signal input
rlabel metal3 s 0 144304 800 144424 6 i_dout1_1[27]
port 116 nsew signal input
rlabel metal3 s 163980 138048 164780 138168 6 i_dout1_1[28]
port 117 nsew signal input
rlabel metal2 s 163226 166124 163282 166924 6 i_dout1_1[29]
port 118 nsew signal input
rlabel metal2 s 147586 0 147642 800 6 i_dout1_1[2]
port 119 nsew signal input
rlabel metal3 s 163980 154504 164780 154624 6 i_dout1_1[30]
port 120 nsew signal input
rlabel metal2 s 164514 0 164570 800 6 i_dout1_1[31]
port 121 nsew signal input
rlabel metal2 s 148230 0 148286 800 6 i_dout1_1[3]
port 122 nsew signal input
rlabel metal2 s 122746 166124 122802 166924 6 i_dout1_1[4]
port 123 nsew signal input
rlabel metal2 s 124770 166124 124826 166924 6 i_dout1_1[5]
port 124 nsew signal input
rlabel metal2 s 150806 0 150862 800 6 i_dout1_1[6]
port 125 nsew signal input
rlabel metal3 s 0 63928 800 64048 6 i_dout1_1[7]
port 126 nsew signal input
rlabel metal3 s 0 66920 800 67040 6 i_dout1_1[8]
port 127 nsew signal input
rlabel metal2 s 154670 0 154726 800 6 i_dout1_1[9]
port 128 nsew signal input
rlabel metal2 s 478 166124 534 166924 6 io_in[0]
port 129 nsew signal input
rlabel metal2 s 30010 166124 30066 166924 6 io_in[10]
port 130 nsew signal input
rlabel metal2 s 32954 166124 33010 166924 6 io_in[11]
port 131 nsew signal input
rlabel metal2 s 35990 166124 36046 166924 6 io_in[12]
port 132 nsew signal input
rlabel metal2 s 38934 166124 38990 166924 6 io_in[13]
port 133 nsew signal input
rlabel metal2 s 41878 166124 41934 166924 6 io_in[14]
port 134 nsew signal input
rlabel metal2 s 44822 166124 44878 166924 6 io_in[15]
port 135 nsew signal input
rlabel metal2 s 47766 166124 47822 166924 6 io_in[16]
port 136 nsew signal input
rlabel metal2 s 50710 166124 50766 166924 6 io_in[17]
port 137 nsew signal input
rlabel metal2 s 53746 166124 53802 166924 6 io_in[18]
port 138 nsew signal input
rlabel metal2 s 56690 166124 56746 166924 6 io_in[19]
port 139 nsew signal input
rlabel metal2 s 3422 166124 3478 166924 6 io_in[1]
port 140 nsew signal input
rlabel metal2 s 59634 166124 59690 166924 6 io_in[20]
port 141 nsew signal input
rlabel metal2 s 62578 166124 62634 166924 6 io_in[21]
port 142 nsew signal input
rlabel metal2 s 65522 166124 65578 166924 6 io_in[22]
port 143 nsew signal input
rlabel metal2 s 68466 166124 68522 166924 6 io_in[23]
port 144 nsew signal input
rlabel metal2 s 71502 166124 71558 166924 6 io_in[24]
port 145 nsew signal input
rlabel metal2 s 74446 166124 74502 166924 6 io_in[25]
port 146 nsew signal input
rlabel metal2 s 77390 166124 77446 166924 6 io_in[26]
port 147 nsew signal input
rlabel metal2 s 80334 166124 80390 166924 6 io_in[27]
port 148 nsew signal input
rlabel metal2 s 83278 166124 83334 166924 6 io_in[28]
port 149 nsew signal input
rlabel metal2 s 86314 166124 86370 166924 6 io_in[29]
port 150 nsew signal input
rlabel metal2 s 6366 166124 6422 166924 6 io_in[2]
port 151 nsew signal input
rlabel metal2 s 89258 166124 89314 166924 6 io_in[30]
port 152 nsew signal input
rlabel metal2 s 92202 166124 92258 166924 6 io_in[31]
port 153 nsew signal input
rlabel metal2 s 95146 166124 95202 166924 6 io_in[32]
port 154 nsew signal input
rlabel metal2 s 98090 166124 98146 166924 6 io_in[33]
port 155 nsew signal input
rlabel metal2 s 101034 166124 101090 166924 6 io_in[34]
port 156 nsew signal input
rlabel metal2 s 104070 166124 104126 166924 6 io_in[35]
port 157 nsew signal input
rlabel metal2 s 107014 166124 107070 166924 6 io_in[36]
port 158 nsew signal input
rlabel metal2 s 109958 166124 110014 166924 6 io_in[37]
port 159 nsew signal input
rlabel metal2 s 9310 166124 9366 166924 6 io_in[3]
port 160 nsew signal input
rlabel metal2 s 12254 166124 12310 166924 6 io_in[4]
port 161 nsew signal input
rlabel metal2 s 15198 166124 15254 166924 6 io_in[5]
port 162 nsew signal input
rlabel metal2 s 18234 166124 18290 166924 6 io_in[6]
port 163 nsew signal input
rlabel metal2 s 21178 166124 21234 166924 6 io_in[7]
port 164 nsew signal input
rlabel metal2 s 24122 166124 24178 166924 6 io_in[8]
port 165 nsew signal input
rlabel metal2 s 27066 166124 27122 166924 6 io_in[9]
port 166 nsew signal input
rlabel metal2 s 1398 166124 1454 166924 6 io_oeb[0]
port 167 nsew signal output
rlabel metal2 s 31022 166124 31078 166924 6 io_oeb[10]
port 168 nsew signal output
rlabel metal2 s 33966 166124 34022 166924 6 io_oeb[11]
port 169 nsew signal output
rlabel metal2 s 36910 166124 36966 166924 6 io_oeb[12]
port 170 nsew signal output
rlabel metal2 s 39854 166124 39910 166924 6 io_oeb[13]
port 171 nsew signal output
rlabel metal2 s 42890 166124 42946 166924 6 io_oeb[14]
port 172 nsew signal output
rlabel metal2 s 45834 166124 45890 166924 6 io_oeb[15]
port 173 nsew signal output
rlabel metal2 s 48778 166124 48834 166924 6 io_oeb[16]
port 174 nsew signal output
rlabel metal2 s 51722 166124 51778 166924 6 io_oeb[17]
port 175 nsew signal output
rlabel metal2 s 54666 166124 54722 166924 6 io_oeb[18]
port 176 nsew signal output
rlabel metal2 s 57702 166124 57758 166924 6 io_oeb[19]
port 177 nsew signal output
rlabel metal2 s 4342 166124 4398 166924 6 io_oeb[1]
port 178 nsew signal output
rlabel metal2 s 60646 166124 60702 166924 6 io_oeb[20]
port 179 nsew signal output
rlabel metal2 s 63590 166124 63646 166924 6 io_oeb[21]
port 180 nsew signal output
rlabel metal2 s 66534 166124 66590 166924 6 io_oeb[22]
port 181 nsew signal output
rlabel metal2 s 69478 166124 69534 166924 6 io_oeb[23]
port 182 nsew signal output
rlabel metal2 s 72422 166124 72478 166924 6 io_oeb[24]
port 183 nsew signal output
rlabel metal2 s 75458 166124 75514 166924 6 io_oeb[25]
port 184 nsew signal output
rlabel metal2 s 78402 166124 78458 166924 6 io_oeb[26]
port 185 nsew signal output
rlabel metal2 s 81346 166124 81402 166924 6 io_oeb[27]
port 186 nsew signal output
rlabel metal2 s 84290 166124 84346 166924 6 io_oeb[28]
port 187 nsew signal output
rlabel metal2 s 87234 166124 87290 166924 6 io_oeb[29]
port 188 nsew signal output
rlabel metal2 s 7378 166124 7434 166924 6 io_oeb[2]
port 189 nsew signal output
rlabel metal2 s 90178 166124 90234 166924 6 io_oeb[30]
port 190 nsew signal output
rlabel metal2 s 93214 166124 93270 166924 6 io_oeb[31]
port 191 nsew signal output
rlabel metal2 s 96158 166124 96214 166924 6 io_oeb[32]
port 192 nsew signal output
rlabel metal2 s 99102 166124 99158 166924 6 io_oeb[33]
port 193 nsew signal output
rlabel metal2 s 102046 166124 102102 166924 6 io_oeb[34]
port 194 nsew signal output
rlabel metal2 s 104990 166124 105046 166924 6 io_oeb[35]
port 195 nsew signal output
rlabel metal2 s 107934 166124 107990 166924 6 io_oeb[36]
port 196 nsew signal output
rlabel metal2 s 110970 166124 111026 166924 6 io_oeb[37]
port 197 nsew signal output
rlabel metal2 s 10322 166124 10378 166924 6 io_oeb[3]
port 198 nsew signal output
rlabel metal2 s 13266 166124 13322 166924 6 io_oeb[4]
port 199 nsew signal output
rlabel metal2 s 16210 166124 16266 166924 6 io_oeb[5]
port 200 nsew signal output
rlabel metal2 s 19154 166124 19210 166924 6 io_oeb[6]
port 201 nsew signal output
rlabel metal2 s 22098 166124 22154 166924 6 io_oeb[7]
port 202 nsew signal output
rlabel metal2 s 25134 166124 25190 166924 6 io_oeb[8]
port 203 nsew signal output
rlabel metal2 s 28078 166124 28134 166924 6 io_oeb[9]
port 204 nsew signal output
rlabel metal2 s 2410 166124 2466 166924 6 io_out[0]
port 205 nsew signal output
rlabel metal2 s 32034 166124 32090 166924 6 io_out[10]
port 206 nsew signal output
rlabel metal2 s 34978 166124 35034 166924 6 io_out[11]
port 207 nsew signal output
rlabel metal2 s 37922 166124 37978 166924 6 io_out[12]
port 208 nsew signal output
rlabel metal2 s 40866 166124 40922 166924 6 io_out[13]
port 209 nsew signal output
rlabel metal2 s 43810 166124 43866 166924 6 io_out[14]
port 210 nsew signal output
rlabel metal2 s 46846 166124 46902 166924 6 io_out[15]
port 211 nsew signal output
rlabel metal2 s 49790 166124 49846 166924 6 io_out[16]
port 212 nsew signal output
rlabel metal2 s 52734 166124 52790 166924 6 io_out[17]
port 213 nsew signal output
rlabel metal2 s 55678 166124 55734 166924 6 io_out[18]
port 214 nsew signal output
rlabel metal2 s 58622 166124 58678 166924 6 io_out[19]
port 215 nsew signal output
rlabel metal2 s 5354 166124 5410 166924 6 io_out[1]
port 216 nsew signal output
rlabel metal2 s 61566 166124 61622 166924 6 io_out[20]
port 217 nsew signal output
rlabel metal2 s 64602 166124 64658 166924 6 io_out[21]
port 218 nsew signal output
rlabel metal2 s 67546 166124 67602 166924 6 io_out[22]
port 219 nsew signal output
rlabel metal2 s 70490 166124 70546 166924 6 io_out[23]
port 220 nsew signal output
rlabel metal2 s 73434 166124 73490 166924 6 io_out[24]
port 221 nsew signal output
rlabel metal2 s 76378 166124 76434 166924 6 io_out[25]
port 222 nsew signal output
rlabel metal2 s 79322 166124 79378 166924 6 io_out[26]
port 223 nsew signal output
rlabel metal2 s 82358 166124 82414 166924 6 io_out[27]
port 224 nsew signal output
rlabel metal2 s 85302 166124 85358 166924 6 io_out[28]
port 225 nsew signal output
rlabel metal2 s 88246 166124 88302 166924 6 io_out[29]
port 226 nsew signal output
rlabel metal2 s 8298 166124 8354 166924 6 io_out[2]
port 227 nsew signal output
rlabel metal2 s 91190 166124 91246 166924 6 io_out[30]
port 228 nsew signal output
rlabel metal2 s 94134 166124 94190 166924 6 io_out[31]
port 229 nsew signal output
rlabel metal2 s 97170 166124 97226 166924 6 io_out[32]
port 230 nsew signal output
rlabel metal2 s 100114 166124 100170 166924 6 io_out[33]
port 231 nsew signal output
rlabel metal2 s 103058 166124 103114 166924 6 io_out[34]
port 232 nsew signal output
rlabel metal2 s 106002 166124 106058 166924 6 io_out[35]
port 233 nsew signal output
rlabel metal2 s 108946 166124 109002 166924 6 io_out[36]
port 234 nsew signal output
rlabel metal2 s 111890 166124 111946 166924 6 io_out[37]
port 235 nsew signal output
rlabel metal2 s 11242 166124 11298 166924 6 io_out[3]
port 236 nsew signal output
rlabel metal2 s 14278 166124 14334 166924 6 io_out[4]
port 237 nsew signal output
rlabel metal2 s 17222 166124 17278 166924 6 io_out[5]
port 238 nsew signal output
rlabel metal2 s 20166 166124 20222 166924 6 io_out[6]
port 239 nsew signal output
rlabel metal2 s 23110 166124 23166 166924 6 io_out[7]
port 240 nsew signal output
rlabel metal2 s 26054 166124 26110 166924 6 io_out[8]
port 241 nsew signal output
rlabel metal2 s 29090 166124 29146 166924 6 io_out[9]
port 242 nsew signal output
rlabel metal2 s 142986 0 143042 800 6 irq[0]
port 243 nsew signal output
rlabel metal2 s 143262 0 143318 800 6 irq[1]
port 244 nsew signal output
rlabel metal2 s 143538 0 143594 800 6 irq[2]
port 245 nsew signal output
rlabel metal2 s 31022 0 31078 800 6 la_data_in[0]
port 246 nsew signal input
rlabel metal2 s 118422 0 118478 800 6 la_data_in[100]
port 247 nsew signal input
rlabel metal2 s 119342 0 119398 800 6 la_data_in[101]
port 248 nsew signal input
rlabel metal2 s 120262 0 120318 800 6 la_data_in[102]
port 249 nsew signal input
rlabel metal2 s 121090 0 121146 800 6 la_data_in[103]
port 250 nsew signal input
rlabel metal2 s 122010 0 122066 800 6 la_data_in[104]
port 251 nsew signal input
rlabel metal2 s 122838 0 122894 800 6 la_data_in[105]
port 252 nsew signal input
rlabel metal2 s 123758 0 123814 800 6 la_data_in[106]
port 253 nsew signal input
rlabel metal2 s 124586 0 124642 800 6 la_data_in[107]
port 254 nsew signal input
rlabel metal2 s 125506 0 125562 800 6 la_data_in[108]
port 255 nsew signal input
rlabel metal2 s 126334 0 126390 800 6 la_data_in[109]
port 256 nsew signal input
rlabel metal2 s 39762 0 39818 800 6 la_data_in[10]
port 257 nsew signal input
rlabel metal2 s 127254 0 127310 800 6 la_data_in[110]
port 258 nsew signal input
rlabel metal2 s 128082 0 128138 800 6 la_data_in[111]
port 259 nsew signal input
rlabel metal2 s 129002 0 129058 800 6 la_data_in[112]
port 260 nsew signal input
rlabel metal2 s 129830 0 129886 800 6 la_data_in[113]
port 261 nsew signal input
rlabel metal2 s 130750 0 130806 800 6 la_data_in[114]
port 262 nsew signal input
rlabel metal2 s 131578 0 131634 800 6 la_data_in[115]
port 263 nsew signal input
rlabel metal2 s 132498 0 132554 800 6 la_data_in[116]
port 264 nsew signal input
rlabel metal2 s 133326 0 133382 800 6 la_data_in[117]
port 265 nsew signal input
rlabel metal2 s 134246 0 134302 800 6 la_data_in[118]
port 266 nsew signal input
rlabel metal2 s 135074 0 135130 800 6 la_data_in[119]
port 267 nsew signal input
rlabel metal2 s 40590 0 40646 800 6 la_data_in[11]
port 268 nsew signal input
rlabel metal2 s 135994 0 136050 800 6 la_data_in[120]
port 269 nsew signal input
rlabel metal2 s 136822 0 136878 800 6 la_data_in[121]
port 270 nsew signal input
rlabel metal2 s 137742 0 137798 800 6 la_data_in[122]
port 271 nsew signal input
rlabel metal2 s 138570 0 138626 800 6 la_data_in[123]
port 272 nsew signal input
rlabel metal2 s 139490 0 139546 800 6 la_data_in[124]
port 273 nsew signal input
rlabel metal2 s 140318 0 140374 800 6 la_data_in[125]
port 274 nsew signal input
rlabel metal2 s 141238 0 141294 800 6 la_data_in[126]
port 275 nsew signal input
rlabel metal2 s 142066 0 142122 800 6 la_data_in[127]
port 276 nsew signal input
rlabel metal2 s 41510 0 41566 800 6 la_data_in[12]
port 277 nsew signal input
rlabel metal2 s 42338 0 42394 800 6 la_data_in[13]
port 278 nsew signal input
rlabel metal2 s 43258 0 43314 800 6 la_data_in[14]
port 279 nsew signal input
rlabel metal2 s 44086 0 44142 800 6 la_data_in[15]
port 280 nsew signal input
rlabel metal2 s 45006 0 45062 800 6 la_data_in[16]
port 281 nsew signal input
rlabel metal2 s 45834 0 45890 800 6 la_data_in[17]
port 282 nsew signal input
rlabel metal2 s 46754 0 46810 800 6 la_data_in[18]
port 283 nsew signal input
rlabel metal2 s 47582 0 47638 800 6 la_data_in[19]
port 284 nsew signal input
rlabel metal2 s 31850 0 31906 800 6 la_data_in[1]
port 285 nsew signal input
rlabel metal2 s 48502 0 48558 800 6 la_data_in[20]
port 286 nsew signal input
rlabel metal2 s 49330 0 49386 800 6 la_data_in[21]
port 287 nsew signal input
rlabel metal2 s 50250 0 50306 800 6 la_data_in[22]
port 288 nsew signal input
rlabel metal2 s 51078 0 51134 800 6 la_data_in[23]
port 289 nsew signal input
rlabel metal2 s 51998 0 52054 800 6 la_data_in[24]
port 290 nsew signal input
rlabel metal2 s 52826 0 52882 800 6 la_data_in[25]
port 291 nsew signal input
rlabel metal2 s 53746 0 53802 800 6 la_data_in[26]
port 292 nsew signal input
rlabel metal2 s 54574 0 54630 800 6 la_data_in[27]
port 293 nsew signal input
rlabel metal2 s 55494 0 55550 800 6 la_data_in[28]
port 294 nsew signal input
rlabel metal2 s 56322 0 56378 800 6 la_data_in[29]
port 295 nsew signal input
rlabel metal2 s 32770 0 32826 800 6 la_data_in[2]
port 296 nsew signal input
rlabel metal2 s 57242 0 57298 800 6 la_data_in[30]
port 297 nsew signal input
rlabel metal2 s 58070 0 58126 800 6 la_data_in[31]
port 298 nsew signal input
rlabel metal2 s 58990 0 59046 800 6 la_data_in[32]
port 299 nsew signal input
rlabel metal2 s 59818 0 59874 800 6 la_data_in[33]
port 300 nsew signal input
rlabel metal2 s 60738 0 60794 800 6 la_data_in[34]
port 301 nsew signal input
rlabel metal2 s 61566 0 61622 800 6 la_data_in[35]
port 302 nsew signal input
rlabel metal2 s 62486 0 62542 800 6 la_data_in[36]
port 303 nsew signal input
rlabel metal2 s 63314 0 63370 800 6 la_data_in[37]
port 304 nsew signal input
rlabel metal2 s 64234 0 64290 800 6 la_data_in[38]
port 305 nsew signal input
rlabel metal2 s 65062 0 65118 800 6 la_data_in[39]
port 306 nsew signal input
rlabel metal2 s 33598 0 33654 800 6 la_data_in[3]
port 307 nsew signal input
rlabel metal2 s 65982 0 66038 800 6 la_data_in[40]
port 308 nsew signal input
rlabel metal2 s 66810 0 66866 800 6 la_data_in[41]
port 309 nsew signal input
rlabel metal2 s 67730 0 67786 800 6 la_data_in[42]
port 310 nsew signal input
rlabel metal2 s 68558 0 68614 800 6 la_data_in[43]
port 311 nsew signal input
rlabel metal2 s 69478 0 69534 800 6 la_data_in[44]
port 312 nsew signal input
rlabel metal2 s 70306 0 70362 800 6 la_data_in[45]
port 313 nsew signal input
rlabel metal2 s 71226 0 71282 800 6 la_data_in[46]
port 314 nsew signal input
rlabel metal2 s 72054 0 72110 800 6 la_data_in[47]
port 315 nsew signal input
rlabel metal2 s 72974 0 73030 800 6 la_data_in[48]
port 316 nsew signal input
rlabel metal2 s 73802 0 73858 800 6 la_data_in[49]
port 317 nsew signal input
rlabel metal2 s 34518 0 34574 800 6 la_data_in[4]
port 318 nsew signal input
rlabel metal2 s 74722 0 74778 800 6 la_data_in[50]
port 319 nsew signal input
rlabel metal2 s 75642 0 75698 800 6 la_data_in[51]
port 320 nsew signal input
rlabel metal2 s 76470 0 76526 800 6 la_data_in[52]
port 321 nsew signal input
rlabel metal2 s 77390 0 77446 800 6 la_data_in[53]
port 322 nsew signal input
rlabel metal2 s 78218 0 78274 800 6 la_data_in[54]
port 323 nsew signal input
rlabel metal2 s 79138 0 79194 800 6 la_data_in[55]
port 324 nsew signal input
rlabel metal2 s 79966 0 80022 800 6 la_data_in[56]
port 325 nsew signal input
rlabel metal2 s 80886 0 80942 800 6 la_data_in[57]
port 326 nsew signal input
rlabel metal2 s 81714 0 81770 800 6 la_data_in[58]
port 327 nsew signal input
rlabel metal2 s 82634 0 82690 800 6 la_data_in[59]
port 328 nsew signal input
rlabel metal2 s 35346 0 35402 800 6 la_data_in[5]
port 329 nsew signal input
rlabel metal2 s 83462 0 83518 800 6 la_data_in[60]
port 330 nsew signal input
rlabel metal2 s 84382 0 84438 800 6 la_data_in[61]
port 331 nsew signal input
rlabel metal2 s 85210 0 85266 800 6 la_data_in[62]
port 332 nsew signal input
rlabel metal2 s 86130 0 86186 800 6 la_data_in[63]
port 333 nsew signal input
rlabel metal2 s 86958 0 87014 800 6 la_data_in[64]
port 334 nsew signal input
rlabel metal2 s 87878 0 87934 800 6 la_data_in[65]
port 335 nsew signal input
rlabel metal2 s 88706 0 88762 800 6 la_data_in[66]
port 336 nsew signal input
rlabel metal2 s 89626 0 89682 800 6 la_data_in[67]
port 337 nsew signal input
rlabel metal2 s 90454 0 90510 800 6 la_data_in[68]
port 338 nsew signal input
rlabel metal2 s 91374 0 91430 800 6 la_data_in[69]
port 339 nsew signal input
rlabel metal2 s 36266 0 36322 800 6 la_data_in[6]
port 340 nsew signal input
rlabel metal2 s 92202 0 92258 800 6 la_data_in[70]
port 341 nsew signal input
rlabel metal2 s 93122 0 93178 800 6 la_data_in[71]
port 342 nsew signal input
rlabel metal2 s 93950 0 94006 800 6 la_data_in[72]
port 343 nsew signal input
rlabel metal2 s 94870 0 94926 800 6 la_data_in[73]
port 344 nsew signal input
rlabel metal2 s 95698 0 95754 800 6 la_data_in[74]
port 345 nsew signal input
rlabel metal2 s 96618 0 96674 800 6 la_data_in[75]
port 346 nsew signal input
rlabel metal2 s 97446 0 97502 800 6 la_data_in[76]
port 347 nsew signal input
rlabel metal2 s 98366 0 98422 800 6 la_data_in[77]
port 348 nsew signal input
rlabel metal2 s 99194 0 99250 800 6 la_data_in[78]
port 349 nsew signal input
rlabel metal2 s 100114 0 100170 800 6 la_data_in[79]
port 350 nsew signal input
rlabel metal2 s 37094 0 37150 800 6 la_data_in[7]
port 351 nsew signal input
rlabel metal2 s 100942 0 100998 800 6 la_data_in[80]
port 352 nsew signal input
rlabel metal2 s 101862 0 101918 800 6 la_data_in[81]
port 353 nsew signal input
rlabel metal2 s 102690 0 102746 800 6 la_data_in[82]
port 354 nsew signal input
rlabel metal2 s 103610 0 103666 800 6 la_data_in[83]
port 355 nsew signal input
rlabel metal2 s 104438 0 104494 800 6 la_data_in[84]
port 356 nsew signal input
rlabel metal2 s 105358 0 105414 800 6 la_data_in[85]
port 357 nsew signal input
rlabel metal2 s 106186 0 106242 800 6 la_data_in[86]
port 358 nsew signal input
rlabel metal2 s 107106 0 107162 800 6 la_data_in[87]
port 359 nsew signal input
rlabel metal2 s 107934 0 107990 800 6 la_data_in[88]
port 360 nsew signal input
rlabel metal2 s 108854 0 108910 800 6 la_data_in[89]
port 361 nsew signal input
rlabel metal2 s 38014 0 38070 800 6 la_data_in[8]
port 362 nsew signal input
rlabel metal2 s 109682 0 109738 800 6 la_data_in[90]
port 363 nsew signal input
rlabel metal2 s 110602 0 110658 800 6 la_data_in[91]
port 364 nsew signal input
rlabel metal2 s 111430 0 111486 800 6 la_data_in[92]
port 365 nsew signal input
rlabel metal2 s 112350 0 112406 800 6 la_data_in[93]
port 366 nsew signal input
rlabel metal2 s 113178 0 113234 800 6 la_data_in[94]
port 367 nsew signal input
rlabel metal2 s 114098 0 114154 800 6 la_data_in[95]
port 368 nsew signal input
rlabel metal2 s 114926 0 114982 800 6 la_data_in[96]
port 369 nsew signal input
rlabel metal2 s 115846 0 115902 800 6 la_data_in[97]
port 370 nsew signal input
rlabel metal2 s 116674 0 116730 800 6 la_data_in[98]
port 371 nsew signal input
rlabel metal2 s 117594 0 117650 800 6 la_data_in[99]
port 372 nsew signal input
rlabel metal2 s 38842 0 38898 800 6 la_data_in[9]
port 373 nsew signal input
rlabel metal2 s 31298 0 31354 800 6 la_data_out[0]
port 374 nsew signal output
rlabel metal2 s 118790 0 118846 800 6 la_data_out[100]
port 375 nsew signal output
rlabel metal2 s 119618 0 119674 800 6 la_data_out[101]
port 376 nsew signal output
rlabel metal2 s 120538 0 120594 800 6 la_data_out[102]
port 377 nsew signal output
rlabel metal2 s 121366 0 121422 800 6 la_data_out[103]
port 378 nsew signal output
rlabel metal2 s 122286 0 122342 800 6 la_data_out[104]
port 379 nsew signal output
rlabel metal2 s 123114 0 123170 800 6 la_data_out[105]
port 380 nsew signal output
rlabel metal2 s 124034 0 124090 800 6 la_data_out[106]
port 381 nsew signal output
rlabel metal2 s 124862 0 124918 800 6 la_data_out[107]
port 382 nsew signal output
rlabel metal2 s 125782 0 125838 800 6 la_data_out[108]
port 383 nsew signal output
rlabel metal2 s 126610 0 126666 800 6 la_data_out[109]
port 384 nsew signal output
rlabel metal2 s 40038 0 40094 800 6 la_data_out[10]
port 385 nsew signal output
rlabel metal2 s 127530 0 127586 800 6 la_data_out[110]
port 386 nsew signal output
rlabel metal2 s 128358 0 128414 800 6 la_data_out[111]
port 387 nsew signal output
rlabel metal2 s 129278 0 129334 800 6 la_data_out[112]
port 388 nsew signal output
rlabel metal2 s 130106 0 130162 800 6 la_data_out[113]
port 389 nsew signal output
rlabel metal2 s 131026 0 131082 800 6 la_data_out[114]
port 390 nsew signal output
rlabel metal2 s 131854 0 131910 800 6 la_data_out[115]
port 391 nsew signal output
rlabel metal2 s 132774 0 132830 800 6 la_data_out[116]
port 392 nsew signal output
rlabel metal2 s 133602 0 133658 800 6 la_data_out[117]
port 393 nsew signal output
rlabel metal2 s 134522 0 134578 800 6 la_data_out[118]
port 394 nsew signal output
rlabel metal2 s 135350 0 135406 800 6 la_data_out[119]
port 395 nsew signal output
rlabel metal2 s 40866 0 40922 800 6 la_data_out[11]
port 396 nsew signal output
rlabel metal2 s 136270 0 136326 800 6 la_data_out[120]
port 397 nsew signal output
rlabel metal2 s 137098 0 137154 800 6 la_data_out[121]
port 398 nsew signal output
rlabel metal2 s 138018 0 138074 800 6 la_data_out[122]
port 399 nsew signal output
rlabel metal2 s 138846 0 138902 800 6 la_data_out[123]
port 400 nsew signal output
rlabel metal2 s 139766 0 139822 800 6 la_data_out[124]
port 401 nsew signal output
rlabel metal2 s 140594 0 140650 800 6 la_data_out[125]
port 402 nsew signal output
rlabel metal2 s 141514 0 141570 800 6 la_data_out[126]
port 403 nsew signal output
rlabel metal2 s 142342 0 142398 800 6 la_data_out[127]
port 404 nsew signal output
rlabel metal2 s 41786 0 41842 800 6 la_data_out[12]
port 405 nsew signal output
rlabel metal2 s 42614 0 42670 800 6 la_data_out[13]
port 406 nsew signal output
rlabel metal2 s 43534 0 43590 800 6 la_data_out[14]
port 407 nsew signal output
rlabel metal2 s 44362 0 44418 800 6 la_data_out[15]
port 408 nsew signal output
rlabel metal2 s 45282 0 45338 800 6 la_data_out[16]
port 409 nsew signal output
rlabel metal2 s 46110 0 46166 800 6 la_data_out[17]
port 410 nsew signal output
rlabel metal2 s 47030 0 47086 800 6 la_data_out[18]
port 411 nsew signal output
rlabel metal2 s 47858 0 47914 800 6 la_data_out[19]
port 412 nsew signal output
rlabel metal2 s 32126 0 32182 800 6 la_data_out[1]
port 413 nsew signal output
rlabel metal2 s 48778 0 48834 800 6 la_data_out[20]
port 414 nsew signal output
rlabel metal2 s 49606 0 49662 800 6 la_data_out[21]
port 415 nsew signal output
rlabel metal2 s 50526 0 50582 800 6 la_data_out[22]
port 416 nsew signal output
rlabel metal2 s 51354 0 51410 800 6 la_data_out[23]
port 417 nsew signal output
rlabel metal2 s 52274 0 52330 800 6 la_data_out[24]
port 418 nsew signal output
rlabel metal2 s 53102 0 53158 800 6 la_data_out[25]
port 419 nsew signal output
rlabel metal2 s 54022 0 54078 800 6 la_data_out[26]
port 420 nsew signal output
rlabel metal2 s 54850 0 54906 800 6 la_data_out[27]
port 421 nsew signal output
rlabel metal2 s 55770 0 55826 800 6 la_data_out[28]
port 422 nsew signal output
rlabel metal2 s 56598 0 56654 800 6 la_data_out[29]
port 423 nsew signal output
rlabel metal2 s 33046 0 33102 800 6 la_data_out[2]
port 424 nsew signal output
rlabel metal2 s 57518 0 57574 800 6 la_data_out[30]
port 425 nsew signal output
rlabel metal2 s 58346 0 58402 800 6 la_data_out[31]
port 426 nsew signal output
rlabel metal2 s 59266 0 59322 800 6 la_data_out[32]
port 427 nsew signal output
rlabel metal2 s 60186 0 60242 800 6 la_data_out[33]
port 428 nsew signal output
rlabel metal2 s 61014 0 61070 800 6 la_data_out[34]
port 429 nsew signal output
rlabel metal2 s 61934 0 61990 800 6 la_data_out[35]
port 430 nsew signal output
rlabel metal2 s 62762 0 62818 800 6 la_data_out[36]
port 431 nsew signal output
rlabel metal2 s 63682 0 63738 800 6 la_data_out[37]
port 432 nsew signal output
rlabel metal2 s 64510 0 64566 800 6 la_data_out[38]
port 433 nsew signal output
rlabel metal2 s 65430 0 65486 800 6 la_data_out[39]
port 434 nsew signal output
rlabel metal2 s 33874 0 33930 800 6 la_data_out[3]
port 435 nsew signal output
rlabel metal2 s 66258 0 66314 800 6 la_data_out[40]
port 436 nsew signal output
rlabel metal2 s 67178 0 67234 800 6 la_data_out[41]
port 437 nsew signal output
rlabel metal2 s 68006 0 68062 800 6 la_data_out[42]
port 438 nsew signal output
rlabel metal2 s 68926 0 68982 800 6 la_data_out[43]
port 439 nsew signal output
rlabel metal2 s 69754 0 69810 800 6 la_data_out[44]
port 440 nsew signal output
rlabel metal2 s 70674 0 70730 800 6 la_data_out[45]
port 441 nsew signal output
rlabel metal2 s 71502 0 71558 800 6 la_data_out[46]
port 442 nsew signal output
rlabel metal2 s 72422 0 72478 800 6 la_data_out[47]
port 443 nsew signal output
rlabel metal2 s 73250 0 73306 800 6 la_data_out[48]
port 444 nsew signal output
rlabel metal2 s 74170 0 74226 800 6 la_data_out[49]
port 445 nsew signal output
rlabel metal2 s 34794 0 34850 800 6 la_data_out[4]
port 446 nsew signal output
rlabel metal2 s 74998 0 75054 800 6 la_data_out[50]
port 447 nsew signal output
rlabel metal2 s 75918 0 75974 800 6 la_data_out[51]
port 448 nsew signal output
rlabel metal2 s 76746 0 76802 800 6 la_data_out[52]
port 449 nsew signal output
rlabel metal2 s 77666 0 77722 800 6 la_data_out[53]
port 450 nsew signal output
rlabel metal2 s 78494 0 78550 800 6 la_data_out[54]
port 451 nsew signal output
rlabel metal2 s 79414 0 79470 800 6 la_data_out[55]
port 452 nsew signal output
rlabel metal2 s 80242 0 80298 800 6 la_data_out[56]
port 453 nsew signal output
rlabel metal2 s 81162 0 81218 800 6 la_data_out[57]
port 454 nsew signal output
rlabel metal2 s 81990 0 82046 800 6 la_data_out[58]
port 455 nsew signal output
rlabel metal2 s 82910 0 82966 800 6 la_data_out[59]
port 456 nsew signal output
rlabel metal2 s 35622 0 35678 800 6 la_data_out[5]
port 457 nsew signal output
rlabel metal2 s 83738 0 83794 800 6 la_data_out[60]
port 458 nsew signal output
rlabel metal2 s 84658 0 84714 800 6 la_data_out[61]
port 459 nsew signal output
rlabel metal2 s 85486 0 85542 800 6 la_data_out[62]
port 460 nsew signal output
rlabel metal2 s 86406 0 86462 800 6 la_data_out[63]
port 461 nsew signal output
rlabel metal2 s 87234 0 87290 800 6 la_data_out[64]
port 462 nsew signal output
rlabel metal2 s 88154 0 88210 800 6 la_data_out[65]
port 463 nsew signal output
rlabel metal2 s 88982 0 89038 800 6 la_data_out[66]
port 464 nsew signal output
rlabel metal2 s 89902 0 89958 800 6 la_data_out[67]
port 465 nsew signal output
rlabel metal2 s 90730 0 90786 800 6 la_data_out[68]
port 466 nsew signal output
rlabel metal2 s 91650 0 91706 800 6 la_data_out[69]
port 467 nsew signal output
rlabel metal2 s 36542 0 36598 800 6 la_data_out[6]
port 468 nsew signal output
rlabel metal2 s 92478 0 92534 800 6 la_data_out[70]
port 469 nsew signal output
rlabel metal2 s 93398 0 93454 800 6 la_data_out[71]
port 470 nsew signal output
rlabel metal2 s 94226 0 94282 800 6 la_data_out[72]
port 471 nsew signal output
rlabel metal2 s 95146 0 95202 800 6 la_data_out[73]
port 472 nsew signal output
rlabel metal2 s 95974 0 96030 800 6 la_data_out[74]
port 473 nsew signal output
rlabel metal2 s 96894 0 96950 800 6 la_data_out[75]
port 474 nsew signal output
rlabel metal2 s 97722 0 97778 800 6 la_data_out[76]
port 475 nsew signal output
rlabel metal2 s 98642 0 98698 800 6 la_data_out[77]
port 476 nsew signal output
rlabel metal2 s 99470 0 99526 800 6 la_data_out[78]
port 477 nsew signal output
rlabel metal2 s 100390 0 100446 800 6 la_data_out[79]
port 478 nsew signal output
rlabel metal2 s 37370 0 37426 800 6 la_data_out[7]
port 479 nsew signal output
rlabel metal2 s 101218 0 101274 800 6 la_data_out[80]
port 480 nsew signal output
rlabel metal2 s 102138 0 102194 800 6 la_data_out[81]
port 481 nsew signal output
rlabel metal2 s 102966 0 103022 800 6 la_data_out[82]
port 482 nsew signal output
rlabel metal2 s 103886 0 103942 800 6 la_data_out[83]
port 483 nsew signal output
rlabel metal2 s 104714 0 104770 800 6 la_data_out[84]
port 484 nsew signal output
rlabel metal2 s 105634 0 105690 800 6 la_data_out[85]
port 485 nsew signal output
rlabel metal2 s 106554 0 106610 800 6 la_data_out[86]
port 486 nsew signal output
rlabel metal2 s 107382 0 107438 800 6 la_data_out[87]
port 487 nsew signal output
rlabel metal2 s 108302 0 108358 800 6 la_data_out[88]
port 488 nsew signal output
rlabel metal2 s 109130 0 109186 800 6 la_data_out[89]
port 489 nsew signal output
rlabel metal2 s 38290 0 38346 800 6 la_data_out[8]
port 490 nsew signal output
rlabel metal2 s 110050 0 110106 800 6 la_data_out[90]
port 491 nsew signal output
rlabel metal2 s 110878 0 110934 800 6 la_data_out[91]
port 492 nsew signal output
rlabel metal2 s 111798 0 111854 800 6 la_data_out[92]
port 493 nsew signal output
rlabel metal2 s 112626 0 112682 800 6 la_data_out[93]
port 494 nsew signal output
rlabel metal2 s 113546 0 113602 800 6 la_data_out[94]
port 495 nsew signal output
rlabel metal2 s 114374 0 114430 800 6 la_data_out[95]
port 496 nsew signal output
rlabel metal2 s 115294 0 115350 800 6 la_data_out[96]
port 497 nsew signal output
rlabel metal2 s 116122 0 116178 800 6 la_data_out[97]
port 498 nsew signal output
rlabel metal2 s 117042 0 117098 800 6 la_data_out[98]
port 499 nsew signal output
rlabel metal2 s 117870 0 117926 800 6 la_data_out[99]
port 500 nsew signal output
rlabel metal2 s 39118 0 39174 800 6 la_data_out[9]
port 501 nsew signal output
rlabel metal2 s 31574 0 31630 800 6 la_oenb[0]
port 502 nsew signal input
rlabel metal2 s 119066 0 119122 800 6 la_oenb[100]
port 503 nsew signal input
rlabel metal2 s 119894 0 119950 800 6 la_oenb[101]
port 504 nsew signal input
rlabel metal2 s 120814 0 120870 800 6 la_oenb[102]
port 505 nsew signal input
rlabel metal2 s 121642 0 121698 800 6 la_oenb[103]
port 506 nsew signal input
rlabel metal2 s 122562 0 122618 800 6 la_oenb[104]
port 507 nsew signal input
rlabel metal2 s 123390 0 123446 800 6 la_oenb[105]
port 508 nsew signal input
rlabel metal2 s 124310 0 124366 800 6 la_oenb[106]
port 509 nsew signal input
rlabel metal2 s 125138 0 125194 800 6 la_oenb[107]
port 510 nsew signal input
rlabel metal2 s 126058 0 126114 800 6 la_oenb[108]
port 511 nsew signal input
rlabel metal2 s 126886 0 126942 800 6 la_oenb[109]
port 512 nsew signal input
rlabel metal2 s 40314 0 40370 800 6 la_oenb[10]
port 513 nsew signal input
rlabel metal2 s 127806 0 127862 800 6 la_oenb[110]
port 514 nsew signal input
rlabel metal2 s 128634 0 128690 800 6 la_oenb[111]
port 515 nsew signal input
rlabel metal2 s 129554 0 129610 800 6 la_oenb[112]
port 516 nsew signal input
rlabel metal2 s 130382 0 130438 800 6 la_oenb[113]
port 517 nsew signal input
rlabel metal2 s 131302 0 131358 800 6 la_oenb[114]
port 518 nsew signal input
rlabel metal2 s 132130 0 132186 800 6 la_oenb[115]
port 519 nsew signal input
rlabel metal2 s 133050 0 133106 800 6 la_oenb[116]
port 520 nsew signal input
rlabel metal2 s 133878 0 133934 800 6 la_oenb[117]
port 521 nsew signal input
rlabel metal2 s 134798 0 134854 800 6 la_oenb[118]
port 522 nsew signal input
rlabel metal2 s 135718 0 135774 800 6 la_oenb[119]
port 523 nsew signal input
rlabel metal2 s 41142 0 41198 800 6 la_oenb[11]
port 524 nsew signal input
rlabel metal2 s 136546 0 136602 800 6 la_oenb[120]
port 525 nsew signal input
rlabel metal2 s 137466 0 137522 800 6 la_oenb[121]
port 526 nsew signal input
rlabel metal2 s 138294 0 138350 800 6 la_oenb[122]
port 527 nsew signal input
rlabel metal2 s 139214 0 139270 800 6 la_oenb[123]
port 528 nsew signal input
rlabel metal2 s 140042 0 140098 800 6 la_oenb[124]
port 529 nsew signal input
rlabel metal2 s 140962 0 141018 800 6 la_oenb[125]
port 530 nsew signal input
rlabel metal2 s 141790 0 141846 800 6 la_oenb[126]
port 531 nsew signal input
rlabel metal2 s 142710 0 142766 800 6 la_oenb[127]
port 532 nsew signal input
rlabel metal2 s 42062 0 42118 800 6 la_oenb[12]
port 533 nsew signal input
rlabel metal2 s 42890 0 42946 800 6 la_oenb[13]
port 534 nsew signal input
rlabel metal2 s 43810 0 43866 800 6 la_oenb[14]
port 535 nsew signal input
rlabel metal2 s 44638 0 44694 800 6 la_oenb[15]
port 536 nsew signal input
rlabel metal2 s 45558 0 45614 800 6 la_oenb[16]
port 537 nsew signal input
rlabel metal2 s 46478 0 46534 800 6 la_oenb[17]
port 538 nsew signal input
rlabel metal2 s 47306 0 47362 800 6 la_oenb[18]
port 539 nsew signal input
rlabel metal2 s 48226 0 48282 800 6 la_oenb[19]
port 540 nsew signal input
rlabel metal2 s 32402 0 32458 800 6 la_oenb[1]
port 541 nsew signal input
rlabel metal2 s 49054 0 49110 800 6 la_oenb[20]
port 542 nsew signal input
rlabel metal2 s 49974 0 50030 800 6 la_oenb[21]
port 543 nsew signal input
rlabel metal2 s 50802 0 50858 800 6 la_oenb[22]
port 544 nsew signal input
rlabel metal2 s 51722 0 51778 800 6 la_oenb[23]
port 545 nsew signal input
rlabel metal2 s 52550 0 52606 800 6 la_oenb[24]
port 546 nsew signal input
rlabel metal2 s 53470 0 53526 800 6 la_oenb[25]
port 547 nsew signal input
rlabel metal2 s 54298 0 54354 800 6 la_oenb[26]
port 548 nsew signal input
rlabel metal2 s 55218 0 55274 800 6 la_oenb[27]
port 549 nsew signal input
rlabel metal2 s 56046 0 56102 800 6 la_oenb[28]
port 550 nsew signal input
rlabel metal2 s 56966 0 57022 800 6 la_oenb[29]
port 551 nsew signal input
rlabel metal2 s 33322 0 33378 800 6 la_oenb[2]
port 552 nsew signal input
rlabel metal2 s 57794 0 57850 800 6 la_oenb[30]
port 553 nsew signal input
rlabel metal2 s 58714 0 58770 800 6 la_oenb[31]
port 554 nsew signal input
rlabel metal2 s 59542 0 59598 800 6 la_oenb[32]
port 555 nsew signal input
rlabel metal2 s 60462 0 60518 800 6 la_oenb[33]
port 556 nsew signal input
rlabel metal2 s 61290 0 61346 800 6 la_oenb[34]
port 557 nsew signal input
rlabel metal2 s 62210 0 62266 800 6 la_oenb[35]
port 558 nsew signal input
rlabel metal2 s 63038 0 63094 800 6 la_oenb[36]
port 559 nsew signal input
rlabel metal2 s 63958 0 64014 800 6 la_oenb[37]
port 560 nsew signal input
rlabel metal2 s 64786 0 64842 800 6 la_oenb[38]
port 561 nsew signal input
rlabel metal2 s 65706 0 65762 800 6 la_oenb[39]
port 562 nsew signal input
rlabel metal2 s 34150 0 34206 800 6 la_oenb[3]
port 563 nsew signal input
rlabel metal2 s 66534 0 66590 800 6 la_oenb[40]
port 564 nsew signal input
rlabel metal2 s 67454 0 67510 800 6 la_oenb[41]
port 565 nsew signal input
rlabel metal2 s 68282 0 68338 800 6 la_oenb[42]
port 566 nsew signal input
rlabel metal2 s 69202 0 69258 800 6 la_oenb[43]
port 567 nsew signal input
rlabel metal2 s 70030 0 70086 800 6 la_oenb[44]
port 568 nsew signal input
rlabel metal2 s 70950 0 71006 800 6 la_oenb[45]
port 569 nsew signal input
rlabel metal2 s 71778 0 71834 800 6 la_oenb[46]
port 570 nsew signal input
rlabel metal2 s 72698 0 72754 800 6 la_oenb[47]
port 571 nsew signal input
rlabel metal2 s 73526 0 73582 800 6 la_oenb[48]
port 572 nsew signal input
rlabel metal2 s 74446 0 74502 800 6 la_oenb[49]
port 573 nsew signal input
rlabel metal2 s 35070 0 35126 800 6 la_oenb[4]
port 574 nsew signal input
rlabel metal2 s 75274 0 75330 800 6 la_oenb[50]
port 575 nsew signal input
rlabel metal2 s 76194 0 76250 800 6 la_oenb[51]
port 576 nsew signal input
rlabel metal2 s 77022 0 77078 800 6 la_oenb[52]
port 577 nsew signal input
rlabel metal2 s 77942 0 77998 800 6 la_oenb[53]
port 578 nsew signal input
rlabel metal2 s 78770 0 78826 800 6 la_oenb[54]
port 579 nsew signal input
rlabel metal2 s 79690 0 79746 800 6 la_oenb[55]
port 580 nsew signal input
rlabel metal2 s 80518 0 80574 800 6 la_oenb[56]
port 581 nsew signal input
rlabel metal2 s 81438 0 81494 800 6 la_oenb[57]
port 582 nsew signal input
rlabel metal2 s 82266 0 82322 800 6 la_oenb[58]
port 583 nsew signal input
rlabel metal2 s 83186 0 83242 800 6 la_oenb[59]
port 584 nsew signal input
rlabel metal2 s 35898 0 35954 800 6 la_oenb[5]
port 585 nsew signal input
rlabel metal2 s 84014 0 84070 800 6 la_oenb[60]
port 586 nsew signal input
rlabel metal2 s 84934 0 84990 800 6 la_oenb[61]
port 587 nsew signal input
rlabel metal2 s 85762 0 85818 800 6 la_oenb[62]
port 588 nsew signal input
rlabel metal2 s 86682 0 86738 800 6 la_oenb[63]
port 589 nsew signal input
rlabel metal2 s 87510 0 87566 800 6 la_oenb[64]
port 590 nsew signal input
rlabel metal2 s 88430 0 88486 800 6 la_oenb[65]
port 591 nsew signal input
rlabel metal2 s 89258 0 89314 800 6 la_oenb[66]
port 592 nsew signal input
rlabel metal2 s 90178 0 90234 800 6 la_oenb[67]
port 593 nsew signal input
rlabel metal2 s 91098 0 91154 800 6 la_oenb[68]
port 594 nsew signal input
rlabel metal2 s 91926 0 91982 800 6 la_oenb[69]
port 595 nsew signal input
rlabel metal2 s 36818 0 36874 800 6 la_oenb[6]
port 596 nsew signal input
rlabel metal2 s 92846 0 92902 800 6 la_oenb[70]
port 597 nsew signal input
rlabel metal2 s 93674 0 93730 800 6 la_oenb[71]
port 598 nsew signal input
rlabel metal2 s 94594 0 94650 800 6 la_oenb[72]
port 599 nsew signal input
rlabel metal2 s 95422 0 95478 800 6 la_oenb[73]
port 600 nsew signal input
rlabel metal2 s 96342 0 96398 800 6 la_oenb[74]
port 601 nsew signal input
rlabel metal2 s 97170 0 97226 800 6 la_oenb[75]
port 602 nsew signal input
rlabel metal2 s 98090 0 98146 800 6 la_oenb[76]
port 603 nsew signal input
rlabel metal2 s 98918 0 98974 800 6 la_oenb[77]
port 604 nsew signal input
rlabel metal2 s 99838 0 99894 800 6 la_oenb[78]
port 605 nsew signal input
rlabel metal2 s 100666 0 100722 800 6 la_oenb[79]
port 606 nsew signal input
rlabel metal2 s 37646 0 37702 800 6 la_oenb[7]
port 607 nsew signal input
rlabel metal2 s 101586 0 101642 800 6 la_oenb[80]
port 608 nsew signal input
rlabel metal2 s 102414 0 102470 800 6 la_oenb[81]
port 609 nsew signal input
rlabel metal2 s 103334 0 103390 800 6 la_oenb[82]
port 610 nsew signal input
rlabel metal2 s 104162 0 104218 800 6 la_oenb[83]
port 611 nsew signal input
rlabel metal2 s 105082 0 105138 800 6 la_oenb[84]
port 612 nsew signal input
rlabel metal2 s 105910 0 105966 800 6 la_oenb[85]
port 613 nsew signal input
rlabel metal2 s 106830 0 106886 800 6 la_oenb[86]
port 614 nsew signal input
rlabel metal2 s 107658 0 107714 800 6 la_oenb[87]
port 615 nsew signal input
rlabel metal2 s 108578 0 108634 800 6 la_oenb[88]
port 616 nsew signal input
rlabel metal2 s 109406 0 109462 800 6 la_oenb[89]
port 617 nsew signal input
rlabel metal2 s 38566 0 38622 800 6 la_oenb[8]
port 618 nsew signal input
rlabel metal2 s 110326 0 110382 800 6 la_oenb[90]
port 619 nsew signal input
rlabel metal2 s 111154 0 111210 800 6 la_oenb[91]
port 620 nsew signal input
rlabel metal2 s 112074 0 112130 800 6 la_oenb[92]
port 621 nsew signal input
rlabel metal2 s 112902 0 112958 800 6 la_oenb[93]
port 622 nsew signal input
rlabel metal2 s 113822 0 113878 800 6 la_oenb[94]
port 623 nsew signal input
rlabel metal2 s 114650 0 114706 800 6 la_oenb[95]
port 624 nsew signal input
rlabel metal2 s 115570 0 115626 800 6 la_oenb[96]
port 625 nsew signal input
rlabel metal2 s 116398 0 116454 800 6 la_oenb[97]
port 626 nsew signal input
rlabel metal2 s 117318 0 117374 800 6 la_oenb[98]
port 627 nsew signal input
rlabel metal2 s 118146 0 118202 800 6 la_oenb[99]
port 628 nsew signal input
rlabel metal2 s 39394 0 39450 800 6 la_oenb[9]
port 629 nsew signal input
rlabel metal3 s 0 7216 800 7336 6 o_addr1[0]
port 630 nsew signal output
rlabel metal3 s 0 16192 800 16312 6 o_addr1[1]
port 631 nsew signal output
rlabel metal3 s 0 25168 800 25288 6 o_addr1[2]
port 632 nsew signal output
rlabel metal3 s 0 34144 800 34264 6 o_addr1[3]
port 633 nsew signal output
rlabel metal3 s 0 45976 800 46096 6 o_addr1[4]
port 634 nsew signal output
rlabel metal2 s 150254 0 150310 800 6 o_addr1[5]
port 635 nsew signal output
rlabel metal3 s 0 60936 800 61056 6 o_addr1[6]
port 636 nsew signal output
rlabel metal2 s 128726 166124 128782 166924 6 o_addr1[7]
port 637 nsew signal output
rlabel metal2 s 154026 0 154082 800 6 o_addr1[8]
port 638 nsew signal output
rlabel metal3 s 0 4224 800 4344 6 o_addr1_1[0]
port 639 nsew signal output
rlabel metal2 s 146206 0 146262 800 6 o_addr1_1[1]
port 640 nsew signal output
rlabel metal3 s 0 22176 800 22296 6 o_addr1_1[2]
port 641 nsew signal output
rlabel metal3 s 163980 31424 164780 31544 6 o_addr1_1[3]
port 642 nsew signal output
rlabel metal3 s 163980 36864 164780 36984 6 o_addr1_1[4]
port 643 nsew signal output
rlabel metal3 s 0 48968 800 49088 6 o_addr1_1[5]
port 644 nsew signal output
rlabel metal2 s 126702 166124 126758 166924 6 o_addr1_1[6]
port 645 nsew signal output
rlabel metal2 s 152554 0 152610 800 6 o_addr1_1[7]
port 646 nsew signal output
rlabel metal2 s 131670 166124 131726 166924 6 o_addr1_1[8]
port 647 nsew signal output
rlabel metal2 s 143814 0 143870 800 6 o_csb0
port 648 nsew signal output
rlabel metal2 s 144090 0 144146 800 6 o_csb0_1
port 649 nsew signal output
rlabel metal3 s 0 1368 800 1488 6 o_csb1
port 650 nsew signal output
rlabel metal3 s 163980 1368 164780 1488 6 o_csb1_1
port 651 nsew signal output
rlabel metal2 s 145010 0 145066 800 6 o_din0[0]
port 652 nsew signal output
rlabel metal3 s 163980 69640 164780 69760 6 o_din0[10]
port 653 nsew signal output
rlabel metal2 s 137558 166124 137614 166924 6 o_din0[11]
port 654 nsew signal output
rlabel metal2 s 138570 166124 138626 166924 6 o_din0[12]
port 655 nsew signal output
rlabel metal2 s 156418 0 156474 800 6 o_din0[13]
port 656 nsew signal output
rlabel metal2 s 156694 0 156750 800 6 o_din0[14]
port 657 nsew signal output
rlabel metal2 s 144458 166124 144514 166924 6 o_din0[15]
port 658 nsew signal output
rlabel metal2 s 157798 0 157854 800 6 o_din0[16]
port 659 nsew signal output
rlabel metal2 s 147402 166124 147458 166924 6 o_din0[17]
port 660 nsew signal output
rlabel metal3 s 0 105544 800 105664 6 o_din0[18]
port 661 nsew signal output
rlabel metal2 s 159546 0 159602 800 6 o_din0[19]
port 662 nsew signal output
rlabel metal2 s 146758 0 146814 800 6 o_din0[1]
port 663 nsew signal output
rlabel metal2 s 152370 166124 152426 166924 6 o_din0[20]
port 664 nsew signal output
rlabel metal3 s 163980 113432 164780 113552 6 o_din0[21]
port 665 nsew signal output
rlabel metal3 s 163980 118872 164780 118992 6 o_din0[22]
port 666 nsew signal output
rlabel metal2 s 161938 0 161994 800 6 o_din0[23]
port 667 nsew signal output
rlabel metal2 s 156326 166124 156382 166924 6 o_din0[24]
port 668 nsew signal output
rlabel metal3 s 163980 129888 164780 130008 6 o_din0[25]
port 669 nsew signal output
rlabel metal3 s 0 141312 800 141432 6 o_din0[26]
port 670 nsew signal output
rlabel metal2 s 160282 166124 160338 166924 6 o_din0[27]
port 671 nsew signal output
rlabel metal2 s 162214 166124 162270 166924 6 o_din0[28]
port 672 nsew signal output
rlabel metal3 s 163980 151784 164780 151904 6 o_din0[29]
port 673 nsew signal output
rlabel metal3 s 163980 20408 164780 20528 6 o_din0[2]
port 674 nsew signal output
rlabel metal3 s 163980 157224 164780 157344 6 o_din0[30]
port 675 nsew signal output
rlabel metal3 s 163980 165384 164780 165504 6 o_din0[31]
port 676 nsew signal output
rlabel metal3 s 0 37000 800 37120 6 o_din0[3]
port 677 nsew signal output
rlabel metal2 s 149334 0 149390 800 6 o_din0[4]
port 678 nsew signal output
rlabel metal3 s 0 54952 800 55072 6 o_din0[5]
port 679 nsew signal output
rlabel metal3 s 163980 47744 164780 47864 6 o_din0[6]
port 680 nsew signal output
rlabel metal2 s 129646 166124 129702 166924 6 o_din0[7]
port 681 nsew signal output
rlabel metal3 s 0 69776 800 69896 6 o_din0[8]
port 682 nsew signal output
rlabel metal2 s 133602 166124 133658 166924 6 o_din0[9]
port 683 nsew signal output
rlabel metal3 s 0 10208 800 10328 6 o_din0_1[0]
port 684 nsew signal output
rlabel metal2 s 135626 166124 135682 166924 6 o_din0_1[10]
port 685 nsew signal output
rlabel metal2 s 155222 0 155278 800 6 o_din0_1[11]
port 686 nsew signal output
rlabel metal3 s 163980 80656 164780 80776 6 o_din0_1[12]
port 687 nsew signal output
rlabel metal3 s 0 93712 800 93832 6 o_din0_1[13]
port 688 nsew signal output
rlabel metal2 s 140502 166124 140558 166924 6 o_din0_1[14]
port 689 nsew signal output
rlabel metal3 s 0 96704 800 96824 6 o_din0_1[15]
port 690 nsew signal output
rlabel metal2 s 157522 0 157578 800 6 o_din0_1[16]
port 691 nsew signal output
rlabel metal2 s 158442 0 158498 800 6 o_din0_1[17]
port 692 nsew signal output
rlabel metal2 s 149426 166124 149482 166924 6 o_din0_1[18]
port 693 nsew signal output
rlabel metal3 s 0 111528 800 111648 6 o_din0_1[19]
port 694 nsew signal output
rlabel metal2 s 146482 0 146538 800 6 o_din0_1[1]
port 695 nsew signal output
rlabel metal2 s 151358 166124 151414 166924 6 o_din0_1[20]
port 696 nsew signal output
rlabel metal3 s 163980 110712 164780 110832 6 o_din0_1[21]
port 697 nsew signal output
rlabel metal2 s 161018 0 161074 800 6 o_din0_1[22]
port 698 nsew signal output
rlabel metal2 s 161662 0 161718 800 6 o_din0_1[23]
port 699 nsew signal output
rlabel metal3 s 163980 124448 164780 124568 6 o_din0_1[24]
port 700 nsew signal output
rlabel metal2 s 162766 0 162822 800 6 o_din0_1[25]
port 701 nsew signal output
rlabel metal3 s 0 138320 800 138440 6 o_din0_1[26]
port 702 nsew signal output
rlabel metal3 s 163980 135328 164780 135448 6 o_din0_1[27]
port 703 nsew signal output
rlabel metal3 s 163980 143488 164780 143608 6 o_din0_1[28]
port 704 nsew signal output
rlabel metal2 s 164238 166124 164294 166924 6 o_din0_1[29]
port 705 nsew signal output
rlabel metal2 s 118790 166124 118846 166924 6 o_din0_1[2]
port 706 nsew signal output
rlabel metal3 s 0 159264 800 159384 6 o_din0_1[30]
port 707 nsew signal output
rlabel metal3 s 0 165248 800 165368 6 o_din0_1[31]
port 708 nsew signal output
rlabel metal2 s 148506 0 148562 800 6 o_din0_1[3]
port 709 nsew signal output
rlabel metal2 s 149058 0 149114 800 6 o_din0_1[4]
port 710 nsew signal output
rlabel metal3 s 0 51960 800 52080 6 o_din0_1[5]
port 711 nsew signal output
rlabel metal2 s 151726 0 151782 800 6 o_din0_1[6]
port 712 nsew signal output
rlabel metal3 s 163980 56040 164780 56160 6 o_din0_1[7]
port 713 nsew signal output
rlabel metal2 s 154302 0 154358 800 6 o_din0_1[8]
port 714 nsew signal output
rlabel metal3 s 0 78752 800 78872 6 o_din0_1[9]
port 715 nsew signal output
rlabel metal3 s 163980 9528 164780 9648 6 o_waddr0[0]
port 716 nsew signal output
rlabel metal2 s 147034 0 147090 800 6 o_waddr0[1]
port 717 nsew signal output
rlabel metal3 s 163980 23128 164780 23248 6 o_waddr0[2]
port 718 nsew signal output
rlabel metal3 s 0 39992 800 40112 6 o_waddr0[3]
port 719 nsew signal output
rlabel metal3 s 163980 42304 164780 42424 6 o_waddr0[4]
port 720 nsew signal output
rlabel metal2 s 150530 0 150586 800 6 o_waddr0[5]
port 721 nsew signal output
rlabel metal3 s 163980 50600 164780 50720 6 o_waddr0[6]
port 722 nsew signal output
rlabel metal2 s 152922 0 152978 800 6 o_waddr0[7]
port 723 nsew signal output
rlabel metal3 s 0 72768 800 72888 6 o_waddr0[8]
port 724 nsew signal output
rlabel metal2 s 145286 0 145342 800 6 o_waddr0_1[0]
port 725 nsew signal output
rlabel metal2 s 115846 166124 115902 166924 6 o_waddr0_1[1]
port 726 nsew signal output
rlabel metal3 s 0 28160 800 28280 6 o_waddr0_1[2]
port 727 nsew signal output
rlabel metal2 s 120814 166124 120870 166924 6 o_waddr0_1[3]
port 728 nsew signal output
rlabel metal3 s 163980 39584 164780 39704 6 o_waddr0_1[4]
port 729 nsew signal output
rlabel metal3 s 0 57944 800 58064 6 o_waddr0_1[5]
port 730 nsew signal output
rlabel metal2 s 127714 166124 127770 166924 6 o_waddr0_1[6]
port 731 nsew signal output
rlabel metal2 s 130658 166124 130714 166924 6 o_waddr0_1[7]
port 732 nsew signal output
rlabel metal3 s 163980 58760 164780 58880 6 o_waddr0_1[8]
port 733 nsew signal output
rlabel metal2 s 112902 166124 112958 166924 6 o_web0
port 734 nsew signal output
rlabel metal2 s 113914 166124 113970 166924 6 o_web0_1
port 735 nsew signal output
rlabel metal2 s 114926 166124 114982 166924 6 o_wmask0[0]
port 736 nsew signal output
rlabel metal2 s 116858 166124 116914 166924 6 o_wmask0[1]
port 737 nsew signal output
rlabel metal3 s 0 31152 800 31272 6 o_wmask0[2]
port 738 nsew signal output
rlabel metal3 s 163980 34144 164780 34264 6 o_wmask0[3]
port 739 nsew signal output
rlabel metal2 s 145562 0 145618 800 6 o_wmask0_1[0]
port 740 nsew signal output
rlabel metal2 s 147310 0 147366 800 6 o_wmask0_1[1]
port 741 nsew signal output
rlabel metal2 s 147954 0 148010 800 6 o_wmask0_1[2]
port 742 nsew signal output
rlabel metal2 s 121826 166124 121882 166924 6 o_wmask0_1[3]
port 743 nsew signal output
rlabel metal4 s 4208 2128 4528 164336 6 vccd1
port 744 nsew power input
rlabel metal4 s 34928 2128 35248 164336 6 vccd1
port 744 nsew power input
rlabel metal4 s 65648 2128 65968 164336 6 vccd1
port 744 nsew power input
rlabel metal4 s 96368 2128 96688 164336 6 vccd1
port 744 nsew power input
rlabel metal4 s 127088 2128 127408 164336 6 vccd1
port 744 nsew power input
rlabel metal4 s 157808 2128 158128 164336 6 vccd1
port 744 nsew power input
rlabel metal4 s 19568 2128 19888 164336 6 vssd1
port 745 nsew ground input
rlabel metal4 s 50288 2128 50608 164336 6 vssd1
port 745 nsew ground input
rlabel metal4 s 81008 2128 81328 164336 6 vssd1
port 745 nsew ground input
rlabel metal4 s 111728 2128 112048 164336 6 vssd1
port 745 nsew ground input
rlabel metal4 s 142448 2128 142768 164336 6 vssd1
port 745 nsew ground input
rlabel metal2 s 110 0 166 800 6 wb_clk_i
port 746 nsew signal input
rlabel metal2 s 386 0 442 800 6 wb_rst_i
port 747 nsew signal input
rlabel metal2 s 662 0 718 800 6 wbs_ack_o
port 748 nsew signal output
rlabel metal2 s 1858 0 1914 800 6 wbs_adr_i[0]
port 749 nsew signal input
rlabel metal2 s 11702 0 11758 800 6 wbs_adr_i[10]
port 750 nsew signal input
rlabel metal2 s 12622 0 12678 800 6 wbs_adr_i[11]
port 751 nsew signal input
rlabel metal2 s 13450 0 13506 800 6 wbs_adr_i[12]
port 752 nsew signal input
rlabel metal2 s 14370 0 14426 800 6 wbs_adr_i[13]
port 753 nsew signal input
rlabel metal2 s 15198 0 15254 800 6 wbs_adr_i[14]
port 754 nsew signal input
rlabel metal2 s 16118 0 16174 800 6 wbs_adr_i[15]
port 755 nsew signal input
rlabel metal2 s 16946 0 17002 800 6 wbs_adr_i[16]
port 756 nsew signal input
rlabel metal2 s 17866 0 17922 800 6 wbs_adr_i[17]
port 757 nsew signal input
rlabel metal2 s 18694 0 18750 800 6 wbs_adr_i[18]
port 758 nsew signal input
rlabel metal2 s 19614 0 19670 800 6 wbs_adr_i[19]
port 759 nsew signal input
rlabel metal2 s 2962 0 3018 800 6 wbs_adr_i[1]
port 760 nsew signal input
rlabel metal2 s 20442 0 20498 800 6 wbs_adr_i[20]
port 761 nsew signal input
rlabel metal2 s 21362 0 21418 800 6 wbs_adr_i[21]
port 762 nsew signal input
rlabel metal2 s 22190 0 22246 800 6 wbs_adr_i[22]
port 763 nsew signal input
rlabel metal2 s 23110 0 23166 800 6 wbs_adr_i[23]
port 764 nsew signal input
rlabel metal2 s 23938 0 23994 800 6 wbs_adr_i[24]
port 765 nsew signal input
rlabel metal2 s 24858 0 24914 800 6 wbs_adr_i[25]
port 766 nsew signal input
rlabel metal2 s 25686 0 25742 800 6 wbs_adr_i[26]
port 767 nsew signal input
rlabel metal2 s 26606 0 26662 800 6 wbs_adr_i[27]
port 768 nsew signal input
rlabel metal2 s 27434 0 27490 800 6 wbs_adr_i[28]
port 769 nsew signal input
rlabel metal2 s 28354 0 28410 800 6 wbs_adr_i[29]
port 770 nsew signal input
rlabel metal2 s 4158 0 4214 800 6 wbs_adr_i[2]
port 771 nsew signal input
rlabel metal2 s 29182 0 29238 800 6 wbs_adr_i[30]
port 772 nsew signal input
rlabel metal2 s 30102 0 30158 800 6 wbs_adr_i[31]
port 773 nsew signal input
rlabel metal2 s 5354 0 5410 800 6 wbs_adr_i[3]
port 774 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 wbs_adr_i[4]
port 775 nsew signal input
rlabel metal2 s 7378 0 7434 800 6 wbs_adr_i[5]
port 776 nsew signal input
rlabel metal2 s 8206 0 8262 800 6 wbs_adr_i[6]
port 777 nsew signal input
rlabel metal2 s 9126 0 9182 800 6 wbs_adr_i[7]
port 778 nsew signal input
rlabel metal2 s 9954 0 10010 800 6 wbs_adr_i[8]
port 779 nsew signal input
rlabel metal2 s 10874 0 10930 800 6 wbs_adr_i[9]
port 780 nsew signal input
rlabel metal2 s 938 0 994 800 6 wbs_cyc_i
port 781 nsew signal input
rlabel metal2 s 2134 0 2190 800 6 wbs_dat_i[0]
port 782 nsew signal input
rlabel metal2 s 11978 0 12034 800 6 wbs_dat_i[10]
port 783 nsew signal input
rlabel metal2 s 12898 0 12954 800 6 wbs_dat_i[11]
port 784 nsew signal input
rlabel metal2 s 13726 0 13782 800 6 wbs_dat_i[12]
port 785 nsew signal input
rlabel metal2 s 14646 0 14702 800 6 wbs_dat_i[13]
port 786 nsew signal input
rlabel metal2 s 15566 0 15622 800 6 wbs_dat_i[14]
port 787 nsew signal input
rlabel metal2 s 16394 0 16450 800 6 wbs_dat_i[15]
port 788 nsew signal input
rlabel metal2 s 17314 0 17370 800 6 wbs_dat_i[16]
port 789 nsew signal input
rlabel metal2 s 18142 0 18198 800 6 wbs_dat_i[17]
port 790 nsew signal input
rlabel metal2 s 19062 0 19118 800 6 wbs_dat_i[18]
port 791 nsew signal input
rlabel metal2 s 19890 0 19946 800 6 wbs_dat_i[19]
port 792 nsew signal input
rlabel metal2 s 3238 0 3294 800 6 wbs_dat_i[1]
port 793 nsew signal input
rlabel metal2 s 20810 0 20866 800 6 wbs_dat_i[20]
port 794 nsew signal input
rlabel metal2 s 21638 0 21694 800 6 wbs_dat_i[21]
port 795 nsew signal input
rlabel metal2 s 22558 0 22614 800 6 wbs_dat_i[22]
port 796 nsew signal input
rlabel metal2 s 23386 0 23442 800 6 wbs_dat_i[23]
port 797 nsew signal input
rlabel metal2 s 24306 0 24362 800 6 wbs_dat_i[24]
port 798 nsew signal input
rlabel metal2 s 25134 0 25190 800 6 wbs_dat_i[25]
port 799 nsew signal input
rlabel metal2 s 26054 0 26110 800 6 wbs_dat_i[26]
port 800 nsew signal input
rlabel metal2 s 26882 0 26938 800 6 wbs_dat_i[27]
port 801 nsew signal input
rlabel metal2 s 27802 0 27858 800 6 wbs_dat_i[28]
port 802 nsew signal input
rlabel metal2 s 28630 0 28686 800 6 wbs_dat_i[29]
port 803 nsew signal input
rlabel metal2 s 4434 0 4490 800 6 wbs_dat_i[2]
port 804 nsew signal input
rlabel metal2 s 29550 0 29606 800 6 wbs_dat_i[30]
port 805 nsew signal input
rlabel metal2 s 30378 0 30434 800 6 wbs_dat_i[31]
port 806 nsew signal input
rlabel metal2 s 5630 0 5686 800 6 wbs_dat_i[3]
port 807 nsew signal input
rlabel metal2 s 6734 0 6790 800 6 wbs_dat_i[4]
port 808 nsew signal input
rlabel metal2 s 7654 0 7710 800 6 wbs_dat_i[5]
port 809 nsew signal input
rlabel metal2 s 8482 0 8538 800 6 wbs_dat_i[6]
port 810 nsew signal input
rlabel metal2 s 9402 0 9458 800 6 wbs_dat_i[7]
port 811 nsew signal input
rlabel metal2 s 10230 0 10286 800 6 wbs_dat_i[8]
port 812 nsew signal input
rlabel metal2 s 11150 0 11206 800 6 wbs_dat_i[9]
port 813 nsew signal input
rlabel metal2 s 2410 0 2466 800 6 wbs_dat_o[0]
port 814 nsew signal output
rlabel metal2 s 12346 0 12402 800 6 wbs_dat_o[10]
port 815 nsew signal output
rlabel metal2 s 13174 0 13230 800 6 wbs_dat_o[11]
port 816 nsew signal output
rlabel metal2 s 14094 0 14150 800 6 wbs_dat_o[12]
port 817 nsew signal output
rlabel metal2 s 14922 0 14978 800 6 wbs_dat_o[13]
port 818 nsew signal output
rlabel metal2 s 15842 0 15898 800 6 wbs_dat_o[14]
port 819 nsew signal output
rlabel metal2 s 16670 0 16726 800 6 wbs_dat_o[15]
port 820 nsew signal output
rlabel metal2 s 17590 0 17646 800 6 wbs_dat_o[16]
port 821 nsew signal output
rlabel metal2 s 18418 0 18474 800 6 wbs_dat_o[17]
port 822 nsew signal output
rlabel metal2 s 19338 0 19394 800 6 wbs_dat_o[18]
port 823 nsew signal output
rlabel metal2 s 20166 0 20222 800 6 wbs_dat_o[19]
port 824 nsew signal output
rlabel metal2 s 3606 0 3662 800 6 wbs_dat_o[1]
port 825 nsew signal output
rlabel metal2 s 21086 0 21142 800 6 wbs_dat_o[20]
port 826 nsew signal output
rlabel metal2 s 21914 0 21970 800 6 wbs_dat_o[21]
port 827 nsew signal output
rlabel metal2 s 22834 0 22890 800 6 wbs_dat_o[22]
port 828 nsew signal output
rlabel metal2 s 23662 0 23718 800 6 wbs_dat_o[23]
port 829 nsew signal output
rlabel metal2 s 24582 0 24638 800 6 wbs_dat_o[24]
port 830 nsew signal output
rlabel metal2 s 25410 0 25466 800 6 wbs_dat_o[25]
port 831 nsew signal output
rlabel metal2 s 26330 0 26386 800 6 wbs_dat_o[26]
port 832 nsew signal output
rlabel metal2 s 27158 0 27214 800 6 wbs_dat_o[27]
port 833 nsew signal output
rlabel metal2 s 28078 0 28134 800 6 wbs_dat_o[28]
port 834 nsew signal output
rlabel metal2 s 28906 0 28962 800 6 wbs_dat_o[29]
port 835 nsew signal output
rlabel metal2 s 4710 0 4766 800 6 wbs_dat_o[2]
port 836 nsew signal output
rlabel metal2 s 29826 0 29882 800 6 wbs_dat_o[30]
port 837 nsew signal output
rlabel metal2 s 30654 0 30710 800 6 wbs_dat_o[31]
port 838 nsew signal output
rlabel metal2 s 5906 0 5962 800 6 wbs_dat_o[3]
port 839 nsew signal output
rlabel metal2 s 7102 0 7158 800 6 wbs_dat_o[4]
port 840 nsew signal output
rlabel metal2 s 7930 0 7986 800 6 wbs_dat_o[5]
port 841 nsew signal output
rlabel metal2 s 8850 0 8906 800 6 wbs_dat_o[6]
port 842 nsew signal output
rlabel metal2 s 9678 0 9734 800 6 wbs_dat_o[7]
port 843 nsew signal output
rlabel metal2 s 10598 0 10654 800 6 wbs_dat_o[8]
port 844 nsew signal output
rlabel metal2 s 11426 0 11482 800 6 wbs_dat_o[9]
port 845 nsew signal output
rlabel metal2 s 2686 0 2742 800 6 wbs_sel_i[0]
port 846 nsew signal input
rlabel metal2 s 3882 0 3938 800 6 wbs_sel_i[1]
port 847 nsew signal input
rlabel metal2 s 4986 0 5042 800 6 wbs_sel_i[2]
port 848 nsew signal input
rlabel metal2 s 6182 0 6238 800 6 wbs_sel_i[3]
port 849 nsew signal input
rlabel metal2 s 1214 0 1270 800 6 wbs_stb_i
port 850 nsew signal input
rlabel metal2 s 1490 0 1546 800 6 wbs_we_i
port 851 nsew signal input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 164780 166924
string LEFview TRUE
string GDS_FILE /local/caravel_user_project/openlane/user_proj/runs/user_proj/results/magic/user_proj.gds
string GDS_END 79752872
string GDS_START 1315924
<< end >>

