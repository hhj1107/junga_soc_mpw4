VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_proj
  CLASS BLOCK ;
  FOREIGN user_proj ;
  ORIGIN 0.000 0.000 ;
  SIZE 823.065 BY 833.785 ;
  PIN i_dout0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END i_dout0[0]
  PIN i_dout0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 669.850 0.000 670.130 4.000 ;
    END
  END i_dout0[10]
  PIN i_dout0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 449.520 823.065 450.120 ;
    END
  END i_dout0[11]
  PIN i_dout0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 679.050 829.785 679.330 833.785 ;
    END
  END i_dout0[12]
  PIN i_dout0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 503.240 823.065 503.840 ;
    END
  END i_dout0[13]
  PIN i_dout0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 430.480 4.000 431.080 ;
    END
  END i_dout0[14]
  PIN i_dout0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 698.370 829.785 698.650 833.785 ;
    END
  END i_dout0[15]
  PIN i_dout0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 556.960 823.065 557.560 ;
    END
  END i_dout0[16]
  PIN i_dout0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 712.170 0.000 712.450 4.000 ;
    END
  END i_dout0[17]
  PIN i_dout0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 713.090 829.785 713.370 833.785 ;
    END
  END i_dout0[18]
  PIN i_dout0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 722.750 829.785 723.030 833.785 ;
    END
  END i_dout0[19]
  PIN i_dout0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 571.870 829.785 572.150 833.785 ;
    END
  END i_dout0[1]
  PIN i_dout0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 732.410 829.785 732.690 833.785 ;
    END
  END i_dout0[20]
  PIN i_dout0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 599.800 4.000 600.400 ;
    END
  END i_dout0[21]
  PIN i_dout0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 614.080 4.000 614.680 ;
    END
  END i_dout0[22]
  PIN i_dout0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 749.890 0.000 750.170 4.000 ;
    END
  END i_dout0[23]
  PIN i_dout0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 656.240 4.000 656.840 ;
    END
  END i_dout0[24]
  PIN i_dout0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 705.200 823.065 705.800 ;
    END
  END i_dout0[25]
  PIN i_dout0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 768.750 0.000 769.030 4.000 ;
    END
  END i_dout0[26]
  PIN i_dout0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 712.680 4.000 713.280 ;
    END
  END i_dout0[27]
  PIN i_dout0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 787.610 0.000 787.890 4.000 ;
    END
  END i_dout0[28]
  PIN i_dout0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 792.210 0.000 792.490 4.000 ;
    END
  END i_dout0[29]
  PIN i_dout0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 113.600 823.065 114.200 ;
    END
  END i_dout0[2]
  PIN i_dout0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 812.640 823.065 813.240 ;
    END
  END i_dout0[30]
  PIN i_dout0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 811.960 4.000 812.560 ;
    END
  END i_dout0[31]
  PIN i_dout0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 134.000 4.000 134.600 ;
    END
  END i_dout0[3]
  PIN i_dout0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.670 0.000 608.950 4.000 ;
    END
  END i_dout0[4]
  PIN i_dout0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 247.560 823.065 248.160 ;
    END
  END i_dout0[5]
  PIN i_dout0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 641.790 0.000 642.070 4.000 ;
    END
  END i_dout0[6]
  PIN i_dout0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 625.230 829.785 625.510 833.785 ;
    END
  END i_dout0[7]
  PIN i_dout0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 303.320 4.000 303.920 ;
    END
  END i_dout0[8]
  PIN i_dout0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 395.800 823.065 396.400 ;
    END
  END i_dout0[9]
  PIN i_dout0_1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 19.080 823.065 19.680 ;
    END
  END i_dout0_1[0]
  PIN i_dout0_1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 665.250 0.000 665.530 4.000 ;
    END
  END i_dout0_1[10]
  PIN i_dout0_1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 435.920 823.065 436.520 ;
    END
  END i_dout0_1[11]
  PIN i_dout0_1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.990 829.785 674.270 833.785 ;
    END
  END i_dout0_1[12]
  PIN i_dout0_1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 489.640 823.065 490.240 ;
    END
  END i_dout0_1[13]
  PIN i_dout0_1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 693.310 0.000 693.590 4.000 ;
    END
  END i_dout0_1[14]
  PIN i_dout0_1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 458.360 4.000 458.960 ;
    END
  END i_dout0_1[15]
  PIN i_dout0_1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 543.360 823.065 543.960 ;
    END
  END i_dout0_1[16]
  PIN i_dout0_1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 501.200 4.000 501.800 ;
    END
  END i_dout0_1[17]
  PIN i_dout0_1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 529.080 4.000 529.680 ;
    END
  END i_dout0_1[18]
  PIN i_dout0_1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 726.430 0.000 726.710 4.000 ;
    END
  END i_dout0_1[19]
  PIN i_dout0_1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 552.550 0.000 552.830 4.000 ;
    END
  END i_dout0_1[1]
  PIN i_dout0_1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 735.630 0.000 735.910 4.000 ;
    END
  END i_dout0_1[20]
  PIN i_dout0_1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 624.280 823.065 624.880 ;
    END
  END i_dout0_1[21]
  PIN i_dout0_1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 651.480 823.065 652.080 ;
    END
  END i_dout0_1[22]
  PIN i_dout0_1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 745.290 0.000 745.570 4.000 ;
    END
  END i_dout0_1[23]
  PIN i_dout0_1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 776.570 829.785 776.850 833.785 ;
    END
  END i_dout0_1[24]
  PIN i_dout0_1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 691.600 823.065 692.200 ;
    END
  END i_dout0_1[25]
  PIN i_dout0_1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 731.720 823.065 732.320 ;
    END
  END i_dout0_1[26]
  PIN i_dout0_1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 777.950 0.000 778.230 4.000 ;
    END
  END i_dout0_1[27]
  PIN i_dout0_1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 741.240 4.000 741.840 ;
    END
  END i_dout0_1[28]
  PIN i_dout0_1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 810.610 829.785 810.890 833.785 ;
    END
  END i_dout0_1[29]
  PIN i_dout0_1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 100.000 823.065 100.600 ;
    END
  END i_dout0_1[2]
  PIN i_dout0_1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 799.040 823.065 799.640 ;
    END
  END i_dout0_1[30]
  PIN i_dout0_1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 815.670 0.000 815.950 4.000 ;
    END
  END i_dout0_1[31]
  PIN i_dout0_1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.720 4.000 120.320 ;
    END
  END i_dout0_1[3]
  PIN i_dout0_1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 193.840 823.065 194.440 ;
    END
  END i_dout0_1[4]
  PIN i_dout0_1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 601.310 829.785 601.590 833.785 ;
    END
  END i_dout0_1[5]
  PIN i_dout0_1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 610.970 829.785 611.250 833.785 ;
    END
  END i_dout0_1[6]
  PIN i_dout0_1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 328.480 823.065 329.080 ;
    END
  END i_dout0_1[7]
  PIN i_dout0_1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 655.590 0.000 655.870 4.000 ;
    END
  END i_dout0_1[8]
  PIN i_dout0_1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 645.010 829.785 645.290 833.785 ;
    END
  END i_dout0_1[9]
  PIN i_dout1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 562.210 829.785 562.490 833.785 ;
    END
  END i_dout1[0]
  PIN i_dout1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 388.320 4.000 388.920 ;
    END
  END i_dout1[10]
  PIN i_dout1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 463.120 823.065 463.720 ;
    END
  END i_dout1[11]
  PIN i_dout1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 679.510 0.000 679.790 4.000 ;
    END
  END i_dout1[12]
  PIN i_dout1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 684.110 0.000 684.390 4.000 ;
    END
  END i_dout1[13]
  PIN i_dout1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 444.760 4.000 445.360 ;
    END
  END i_dout1[14]
  PIN i_dout1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 703.430 829.785 703.710 833.785 ;
    END
  END i_dout1[15]
  PIN i_dout1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 486.920 4.000 487.520 ;
    END
  END i_dout1[16]
  PIN i_dout1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 716.770 0.000 717.050 4.000 ;
    END
  END i_dout1[17]
  PIN i_dout1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 543.360 4.000 543.960 ;
    END
  END i_dout1[18]
  PIN i_dout1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 731.030 0.000 731.310 4.000 ;
    END
  END i_dout1[19]
  PIN i_dout1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 59.880 823.065 60.480 ;
    END
  END i_dout1[1]
  PIN i_dout1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.470 829.785 737.750 833.785 ;
    END
  END i_dout1[20]
  PIN i_dout1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 740.230 0.000 740.510 4.000 ;
    END
  END i_dout1[21]
  PIN i_dout1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 664.400 823.065 665.000 ;
    END
  END i_dout1[22]
  PIN i_dout1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 642.640 4.000 643.240 ;
    END
  END i_dout1[23]
  PIN i_dout1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 670.520 4.000 671.120 ;
    END
  END i_dout1[24]
  PIN i_dout1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 684.800 4.000 685.400 ;
    END
  END i_dout1[25]
  PIN i_dout1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 790.830 829.785 791.110 833.785 ;
    END
  END i_dout1[26]
  PIN i_dout1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 772.520 823.065 773.120 ;
    END
  END i_dout1[27]
  PIN i_dout1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 755.520 4.000 756.120 ;
    END
  END i_dout1[28]
  PIN i_dout1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 815.210 829.785 815.490 833.785 ;
    END
  END i_dout1[29]
  PIN i_dout1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.880 4.000 77.480 ;
    END
  END i_dout1[2]
  PIN i_dout1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 820.270 829.785 820.550 833.785 ;
    END
  END i_dout1[30]
  PIN i_dout1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 820.270 0.000 820.550 4.000 ;
    END
  END i_dout1[31]
  PIN i_dout1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 594.870 0.000 595.150 4.000 ;
    END
  END i_dout1[3]
  PIN i_dout1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 221.040 823.065 221.640 ;
    END
  END i_dout1[4]
  PIN i_dout1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 261.160 823.065 261.760 ;
    END
  END i_dout1[5]
  PIN i_dout1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 615.570 829.785 615.850 833.785 ;
    END
  END i_dout1[6]
  PIN i_dout1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 630.290 829.785 630.570 833.785 ;
    END
  END i_dout1[7]
  PIN i_dout1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 355.680 823.065 356.280 ;
    END
  END i_dout1[8]
  PIN i_dout1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 654.670 829.785 654.950 833.785 ;
    END
  END i_dout1[9]
  PIN i_dout1_1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END i_dout1_1[0]
  PIN i_dout1_1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 374.040 4.000 374.640 ;
    END
  END i_dout1_1[10]
  PIN i_dout1_1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 664.330 829.785 664.610 833.785 ;
    END
  END i_dout1_1[11]
  PIN i_dout1_1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 674.450 0.000 674.730 4.000 ;
    END
  END i_dout1_1[12]
  PIN i_dout1_1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 684.110 829.785 684.390 833.785 ;
    END
  END i_dout1_1[13]
  PIN i_dout1_1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 516.840 823.065 517.440 ;
    END
  END i_dout1_1[14]
  PIN i_dout1_1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 530.440 823.065 531.040 ;
    END
  END i_dout1_1[15]
  PIN i_dout1_1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 472.640 4.000 473.240 ;
    END
  END i_dout1_1[16]
  PIN i_dout1_1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 515.480 4.000 516.080 ;
    END
  END i_dout1_1[17]
  PIN i_dout1_1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 597.760 823.065 598.360 ;
    END
  END i_dout1_1[18]
  PIN i_dout1_1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 571.920 4.000 572.520 ;
    END
  END i_dout1_1[19]
  PIN i_dout1_1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.000 4.000 49.600 ;
    END
  END i_dout1_1[1]
  PIN i_dout1_1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 585.520 4.000 586.120 ;
    END
  END i_dout1_1[20]
  PIN i_dout1_1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 637.880 823.065 638.480 ;
    END
  END i_dout1_1[21]
  PIN i_dout1_1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 761.850 829.785 762.130 833.785 ;
    END
  END i_dout1_1[22]
  PIN i_dout1_1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 628.360 4.000 628.960 ;
    END
  END i_dout1_1[23]
  PIN i_dout1_1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 678.000 823.065 678.600 ;
    END
  END i_dout1_1[24]
  PIN i_dout1_1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 764.150 0.000 764.430 4.000 ;
    END
  END i_dout1_1[25]
  PIN i_dout1_1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 745.320 823.065 745.920 ;
    END
  END i_dout1_1[26]
  PIN i_dout1_1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 758.920 823.065 759.520 ;
    END
  END i_dout1_1[27]
  PIN i_dout1_1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 800.950 829.785 801.230 833.785 ;
    END
  END i_dout1_1[28]
  PIN i_dout1_1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 785.440 823.065 786.040 ;
    END
  END i_dout1_1[29]
  PIN i_dout1_1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 580.610 0.000 580.890 4.000 ;
    END
  END i_dout1_1[2]
  PIN i_dout1_1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 806.470 0.000 806.750 4.000 ;
    END
  END i_dout1_1[30]
  PIN i_dout1_1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 797.680 4.000 798.280 ;
    END
  END i_dout1_1[31]
  PIN i_dout1_1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 589.810 0.000 590.090 4.000 ;
    END
  END i_dout1_1[3]
  PIN i_dout1_1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 207.440 823.065 208.040 ;
    END
  END i_dout1_1[4]
  PIN i_dout1_1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 190.440 4.000 191.040 ;
    END
  END i_dout1_1[5]
  PIN i_dout1_1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 218.320 4.000 218.920 ;
    END
  END i_dout1_1[6]
  PIN i_dout1_1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 261.160 4.000 261.760 ;
    END
  END i_dout1_1[7]
  PIN i_dout1_1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 660.650 0.000 660.930 4.000 ;
    END
  END i_dout1_1[8]
  PIN i_dout1_1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 649.610 829.785 649.890 833.785 ;
    END
  END i_dout1_1[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.390 829.785 2.670 833.785 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 829.785 148.490 833.785 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.930 829.785 163.210 833.785 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.650 829.785 177.930 833.785 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.910 829.785 192.190 833.785 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.630 829.785 206.910 833.785 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.350 829.785 221.630 833.785 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.070 829.785 236.350 833.785 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.330 829.785 250.610 833.785 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.050 829.785 265.330 833.785 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.770 829.785 280.050 833.785 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.650 829.785 16.930 833.785 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.490 829.785 294.770 833.785 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.750 829.785 309.030 833.785 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.470 829.785 323.750 833.785 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.190 829.785 338.470 833.785 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.910 829.785 353.190 833.785 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.170 829.785 367.450 833.785 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 381.890 829.785 382.170 833.785 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.610 829.785 396.890 833.785 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 411.330 829.785 411.610 833.785 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.590 829.785 425.870 833.785 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.370 829.785 31.650 833.785 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 440.310 829.785 440.590 833.785 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.030 829.785 455.310 833.785 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.750 829.785 470.030 833.785 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.010 829.785 484.290 833.785 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 498.730 829.785 499.010 833.785 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 513.450 829.785 513.730 833.785 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.170 829.785 528.450 833.785 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 542.890 829.785 543.170 833.785 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.090 829.785 46.370 833.785 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.810 829.785 61.090 833.785 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.070 829.785 75.350 833.785 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.790 829.785 90.070 833.785 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.510 829.785 104.790 833.785 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 829.785 119.510 833.785 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.490 829.785 133.770 833.785 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 829.785 7.270 833.785 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.270 829.785 153.550 833.785 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 829.785 167.810 833.785 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.250 829.785 182.530 833.785 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.970 829.785 197.250 833.785 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.690 829.785 211.970 833.785 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.950 829.785 226.230 833.785 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.670 829.785 240.950 833.785 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.390 829.785 255.670 833.785 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.110 829.785 270.390 833.785 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.370 829.785 284.650 833.785 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.710 829.785 21.990 833.785 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.090 829.785 299.370 833.785 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 313.810 829.785 314.090 833.785 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.530 829.785 328.810 833.785 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.250 829.785 343.530 833.785 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.510 829.785 357.790 833.785 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 372.230 829.785 372.510 833.785 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.950 829.785 387.230 833.785 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 401.670 829.785 401.950 833.785 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.930 829.785 416.210 833.785 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 430.650 829.785 430.930 833.785 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.430 829.785 36.710 833.785 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.370 829.785 445.650 833.785 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.090 829.785 460.370 833.785 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 474.350 829.785 474.630 833.785 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.070 829.785 489.350 833.785 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 503.790 829.785 504.070 833.785 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.510 829.785 518.790 833.785 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 532.770 829.785 533.050 833.785 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.490 829.785 547.770 833.785 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.690 829.785 50.970 833.785 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.410 829.785 65.690 833.785 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.130 829.785 80.410 833.785 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.850 829.785 95.130 833.785 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.110 829.785 109.390 833.785 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.830 829.785 124.110 833.785 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 829.785 138.830 833.785 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.050 829.785 12.330 833.785 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 829.785 158.150 833.785 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.590 829.785 172.870 833.785 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.310 829.785 187.590 833.785 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.030 829.785 202.310 833.785 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.290 829.785 216.570 833.785 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.010 829.785 231.290 833.785 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.730 829.785 246.010 833.785 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.450 829.785 260.730 833.785 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.710 829.785 274.990 833.785 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.430 829.785 289.710 833.785 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.310 829.785 26.590 833.785 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.150 829.785 304.430 833.785 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.870 829.785 319.150 833.785 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.130 829.785 333.410 833.785 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.850 829.785 348.130 833.785 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.570 829.785 362.850 833.785 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.290 829.785 377.570 833.785 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.550 829.785 391.830 833.785 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 406.270 829.785 406.550 833.785 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.990 829.785 421.270 833.785 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 435.710 829.785 435.990 833.785 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.030 829.785 41.310 833.785 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.970 829.785 450.250 833.785 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 464.690 829.785 464.970 833.785 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.410 829.785 479.690 833.785 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 494.130 829.785 494.410 833.785 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.390 829.785 508.670 833.785 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 523.110 829.785 523.390 833.785 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.830 829.785 538.110 833.785 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 552.550 829.785 552.830 833.785 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.750 829.785 56.030 833.785 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.470 829.785 70.750 833.785 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.730 829.785 85.010 833.785 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.450 829.785 99.730 833.785 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.170 829.785 114.450 833.785 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 829.785 129.170 833.785 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.150 829.785 143.430 833.785 ;
    END
  END io_out[9]
  PIN irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 500.570 0.000 500.850 4.000 ;
    END
  END irq[0]
  PIN irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.170 0.000 505.450 4.000 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 510.230 0.000 510.510 4.000 ;
    END
  END irq[2]
  PIN o_addr1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 533.690 0.000 533.970 4.000 ;
    END
  END o_addr1[0]
  PIN o_addr1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.150 0.000 557.430 4.000 ;
    END
  END o_addr1[1]
  PIN o_addr1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.160 4.000 91.760 ;
    END
  END o_addr1[2]
  PIN o_addr1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 147.600 4.000 148.200 ;
    END
  END o_addr1[3]
  PIN o_addr1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 613.270 0.000 613.550 4.000 ;
    END
  END o_addr1[4]
  PIN o_addr1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 274.760 823.065 275.360 ;
    END
  END o_addr1[5]
  PIN o_addr1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 301.960 823.065 302.560 ;
    END
  END o_addr1[6]
  PIN o_addr1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 646.390 0.000 646.670 4.000 ;
    END
  END o_addr1[7]
  PIN o_addr1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 317.600 4.000 318.200 ;
    END
  END o_addr1[8]
  PIN o_addr1_1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 566.810 829.785 567.090 833.785 ;
    END
  END o_addr1_1[0]
  PIN o_addr1_1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 72.800 823.065 73.400 ;
    END
  END o_addr1_1[1]
  PIN o_addr1_1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.930 829.785 577.210 833.785 ;
    END
  END o_addr1_1[2]
  PIN o_addr1_1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 591.190 829.785 591.470 833.785 ;
    END
  END o_addr1_1[3]
  PIN o_addr1_1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 596.250 829.785 596.530 833.785 ;
    END
  END o_addr1_1[4]
  PIN o_addr1_1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.040 4.000 204.640 ;
    END
  END o_addr1_1[5]
  PIN o_addr1_1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 288.360 823.065 288.960 ;
    END
  END o_addr1_1[6]
  PIN o_addr1_1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 342.080 823.065 342.680 ;
    END
  END o_addr1_1[7]
  PIN o_addr1_1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 639.950 829.785 640.230 833.785 ;
    END
  END o_addr1_1[8]
  PIN o_csb0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 514.830 0.000 515.110 4.000 ;
    END
  END o_csb0
  PIN o_csb0_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.150 829.785 557.430 833.785 ;
    END
  END o_csb0_1
  PIN o_csb1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 519.430 0.000 519.710 4.000 ;
    END
  END o_csb1
  PIN o_csb1_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 6.160 823.065 6.760 ;
    END
  END o_csb1_1
  PIN o_din0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.720 4.000 35.320 ;
    END
  END o_din0[0]
  PIN o_din0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 659.730 829.785 660.010 833.785 ;
    END
  END o_din0[10]
  PIN o_din0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 669.390 829.785 669.670 833.785 ;
    END
  END o_din0[11]
  PIN o_din0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 416.200 4.000 416.800 ;
    END
  END o_din0[12]
  PIN o_din0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 688.710 829.785 688.990 833.785 ;
    END
  END o_din0[13]
  PIN o_din0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 697.910 0.000 698.190 4.000 ;
    END
  END o_din0[14]
  PIN o_din0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.970 0.000 703.250 4.000 ;
    END
  END o_din0[15]
  PIN o_din0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 570.560 823.065 571.160 ;
    END
  END o_din0[16]
  PIN o_din0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 721.830 0.000 722.110 4.000 ;
    END
  END o_din0[17]
  PIN o_din0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 718.150 829.785 718.430 833.785 ;
    END
  END o_din0[18]
  PIN o_din0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 727.810 829.785 728.090 833.785 ;
    END
  END o_din0[19]
  PIN o_din0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 566.350 0.000 566.630 4.000 ;
    END
  END o_din0[1]
  PIN o_din0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 747.130 829.785 747.410 833.785 ;
    END
  END o_din0[20]
  PIN o_din0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 756.790 829.785 757.070 833.785 ;
    END
  END o_din0[21]
  PIN o_din0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 771.510 829.785 771.790 833.785 ;
    END
  END o_din0[22]
  PIN o_din0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 759.090 0.000 759.370 4.000 ;
    END
  END o_din0[23]
  PIN o_din0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 786.230 829.785 786.510 833.785 ;
    END
  END o_din0[24]
  PIN o_din0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 699.080 4.000 699.680 ;
    END
  END o_din0[25]
  PIN o_din0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 773.350 0.000 773.630 4.000 ;
    END
  END o_din0[26]
  PIN o_din0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 782.550 0.000 782.830 4.000 ;
    END
  END o_din0[27]
  PIN o_din0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 769.800 4.000 770.400 ;
    END
  END o_din0[28]
  PIN o_din0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 801.410 0.000 801.690 4.000 ;
    END
  END o_din0[29]
  PIN o_din0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 4.000 106.040 ;
    END
  END o_din0[2]
  PIN o_din0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 783.400 4.000 784.000 ;
    END
  END o_din0[30]
  PIN o_din0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 826.240 823.065 826.840 ;
    END
  END o_din0[31]
  PIN o_din0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.880 4.000 162.480 ;
    END
  END o_din0[3]
  PIN o_din0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 234.640 823.065 235.240 ;
    END
  END o_din0[4]
  PIN o_din0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.910 829.785 606.190 833.785 ;
    END
  END o_din0[5]
  PIN o_din0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 232.600 4.000 233.200 ;
    END
  END o_din0[6]
  PIN o_din0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 274.760 4.000 275.360 ;
    END
  END o_din0[7]
  PIN o_din0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 345.480 4.000 346.080 ;
    END
  END o_din0[8]
  PIN o_din0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 359.760 4.000 360.360 ;
    END
  END o_din0[9]
  PIN o_din0_1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 538.290 0.000 538.570 4.000 ;
    END
  END o_din0_1[0]
  PIN o_din0_1[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 423.000 823.065 423.600 ;
    END
  END o_din0_1[10]
  PIN o_din0_1[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 476.720 823.065 477.320 ;
    END
  END o_din0_1[11]
  PIN o_din0_1[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 401.920 4.000 402.520 ;
    END
  END o_din0_1[12]
  PIN o_din0_1[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 688.710 0.000 688.990 4.000 ;
    END
  END o_din0_1[13]
  PIN o_din0_1[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 693.770 829.785 694.050 833.785 ;
    END
  END o_din0_1[14]
  PIN o_din0_1[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.030 829.785 708.310 833.785 ;
    END
  END o_din0_1[15]
  PIN o_din0_1[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 707.570 0.000 707.850 4.000 ;
    END
  END o_din0_1[16]
  PIN o_din0_1[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 584.160 823.065 584.760 ;
    END
  END o_din0_1[17]
  PIN o_din0_1[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 557.640 4.000 558.240 ;
    END
  END o_din0_1[18]
  PIN o_din0_1[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 610.680 823.065 611.280 ;
    END
  END o_din0_1[19]
  PIN o_din0_1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 561.750 0.000 562.030 4.000 ;
    END
  END o_din0_1[1]
  PIN o_din0_1[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 742.530 829.785 742.810 833.785 ;
    END
  END o_din0_1[20]
  PIN o_din0_1[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 752.190 829.785 752.470 833.785 ;
    END
  END o_din0_1[21]
  PIN o_din0_1[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 766.450 829.785 766.730 833.785 ;
    END
  END o_din0_1[22]
  PIN o_din0_1[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 754.490 0.000 754.770 4.000 ;
    END
  END o_din0_1[23]
  PIN o_din0_1[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 781.170 829.785 781.450 833.785 ;
    END
  END o_din0_1[24]
  PIN o_din0_1[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 718.800 823.065 719.400 ;
    END
  END o_din0_1[25]
  PIN o_din0_1[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 795.890 829.785 796.170 833.785 ;
    END
  END o_din0_1[26]
  PIN o_din0_1[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 726.960 4.000 727.560 ;
    END
  END o_din0_1[27]
  PIN o_din0_1[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 805.550 829.785 805.830 833.785 ;
    END
  END o_din0_1[28]
  PIN o_din0_1[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 796.810 0.000 797.090 4.000 ;
    END
  END o_din0_1[29]
  PIN o_din0_1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.530 829.785 581.810 833.785 ;
    END
  END o_din0_1[2]
  PIN o_din0_1[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 811.070 0.000 811.350 4.000 ;
    END
  END o_din0_1[30]
  PIN o_din0_1[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 826.240 4.000 826.840 ;
    END
  END o_din0_1[31]
  PIN o_din0_1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.470 0.000 599.750 4.000 ;
    END
  END o_din0_1[3]
  PIN o_din0_1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.160 4.000 176.760 ;
    END
  END o_din0_1[4]
  PIN o_din0_1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.530 0.000 627.810 4.000 ;
    END
  END o_din0_1[5]
  PIN o_din0_1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 620.630 829.785 620.910 833.785 ;
    END
  END o_din0_1[6]
  PIN o_din0_1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 635.350 829.785 635.630 833.785 ;
    END
  END o_din0_1[7]
  PIN o_din0_1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 331.200 4.000 331.800 ;
    END
  END o_din0_1[8]
  PIN o_din0_1[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 409.400 823.065 410.000 ;
    END
  END o_din0_1[9]
  PIN o_waddr0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 32.680 823.065 33.280 ;
    END
  END o_waddr0[0]
  PIN o_waddr0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.280 4.000 63.880 ;
    END
  END o_waddr0[1]
  PIN o_waddr0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 585.210 0.000 585.490 4.000 ;
    END
  END o_waddr0[2]
  PIN o_waddr0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 167.320 823.065 167.920 ;
    END
  END o_waddr0[3]
  PIN o_waddr0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 622.930 0.000 623.210 4.000 ;
    END
  END o_waddr0[4]
  PIN o_waddr0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 637.190 0.000 637.470 4.000 ;
    END
  END o_waddr0[5]
  PIN o_waddr0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 246.880 4.000 247.480 ;
    END
  END o_waddr0[6]
  PIN o_waddr0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 289.040 4.000 289.640 ;
    END
  END o_waddr0[7]
  PIN o_waddr0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 382.200 823.065 382.800 ;
    END
  END o_waddr0[8]
  PIN o_waddr0_1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 542.890 0.000 543.170 4.000 ;
    END
  END o_waddr0_1[0]
  PIN o_waddr0_1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 86.400 823.065 87.000 ;
    END
  END o_waddr0_1[1]
  PIN o_waddr0_1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 126.520 823.065 127.120 ;
    END
  END o_waddr0_1[2]
  PIN o_waddr0_1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 153.720 823.065 154.320 ;
    END
  END o_waddr0_1[3]
  PIN o_waddr0_1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 618.330 0.000 618.610 4.000 ;
    END
  END o_waddr0_1[4]
  PIN o_waddr0_1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 632.130 0.000 632.410 4.000 ;
    END
  END o_waddr0_1[5]
  PIN o_waddr0_1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 314.880 823.065 315.480 ;
    END
  END o_waddr0_1[6]
  PIN o_waddr0_1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.990 0.000 651.270 4.000 ;
    END
  END o_waddr0_1[7]
  PIN o_waddr0_1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 368.600 823.065 369.200 ;
    END
  END o_waddr0_1[8]
  PIN o_web0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.030 0.000 524.310 4.000 ;
    END
  END o_web0
  PIN o_web0_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.630 0.000 528.910 4.000 ;
    END
  END o_web0_1
  PIN o_wmask0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 46.280 823.065 46.880 ;
    END
  END o_wmask0[0]
  PIN o_wmask0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.010 0.000 576.290 4.000 ;
    END
  END o_wmask0[1]
  PIN o_wmask0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 140.120 823.065 140.720 ;
    END
  END o_wmask0[2]
  PIN o_wmask0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 180.920 823.065 181.520 ;
    END
  END o_wmask0[3]
  PIN o_wmask0_1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.490 0.000 547.770 4.000 ;
    END
  END o_wmask0_1[0]
  PIN o_wmask0_1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.950 0.000 571.230 4.000 ;
    END
  END o_wmask0_1[1]
  PIN o_wmask0_1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.590 829.785 586.870 833.785 ;
    END
  END o_wmask0_1[2]
  PIN o_wmask0_1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 604.070 0.000 604.350 4.000 ;
    END
  END o_wmask0_1[3]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 821.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 821.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 821.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 821.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 821.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 821.680 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 821.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 821.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 821.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 821.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 821.680 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.390 0.000 2.670 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 0.000 7.270 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 0.000 11.870 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.450 0.000 30.730 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.070 0.000 190.350 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.330 0.000 204.610 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.590 0.000 218.870 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.390 0.000 232.670 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.650 0.000 246.930 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.910 0.000 261.190 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.710 0.000 274.990 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.970 0.000 289.250 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.230 0.000 303.510 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.030 0.000 317.310 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.310 0.000 49.590 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.290 0.000 331.570 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.550 0.000 345.830 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 359.350 0.000 359.630 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.610 0.000 373.890 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 387.870 0.000 388.150 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 401.670 0.000 401.950 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.930 0.000 416.210 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 430.190 0.000 430.470 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.990 0.000 444.270 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 458.250 0.000 458.530 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.170 0.000 68.450 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.510 0.000 472.790 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 486.310 0.000 486.590 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.430 0.000 105.710 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.690 0.000 119.970 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.950 0.000 134.230 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.750 0.000 148.030 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.010 0.000 162.290 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.270 0.000 176.550 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.050 0.000 35.330 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.130 0.000 195.410 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.930 0.000 209.210 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.190 0.000 223.470 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.450 0.000 237.730 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.250 0.000 251.530 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.510 0.000 265.790 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.770 0.000 280.050 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.570 0.000 293.850 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 307.830 0.000 308.110 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.090 0.000 322.370 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.910 0.000 54.190 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.890 0.000 336.170 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 350.150 0.000 350.430 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.410 0.000 364.690 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.210 0.000 378.490 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.470 0.000 392.750 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 406.730 0.000 407.010 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.530 0.000 420.810 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.790 0.000 435.070 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.050 0.000 449.330 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 462.850 0.000 463.130 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.770 0.000 73.050 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 477.110 0.000 477.390 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 491.370 0.000 491.650 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.630 0.000 91.910 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.490 0.000 110.770 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.290 0.000 124.570 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 0.000 138.830 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.810 0.000 153.090 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.610 0.000 166.890 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.870 0.000 181.150 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.650 0.000 39.930 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.730 0.000 200.010 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.990 0.000 214.270 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.790 0.000 228.070 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.050 0.000 242.330 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.310 0.000 256.590 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.110 0.000 270.390 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.370 0.000 284.650 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.630 0.000 298.910 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.430 0.000 312.710 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.690 0.000 326.970 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.510 0.000 58.790 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.950 0.000 341.230 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.750 0.000 355.030 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.010 0.000 369.290 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.270 0.000 383.550 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.070 0.000 397.350 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 411.330 0.000 411.610 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.590 0.000 425.870 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.390 0.000 439.670 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 453.650 0.000 453.930 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 467.910 0.000 468.190 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 481.710 0.000 481.990 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.970 0.000 496.250 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.230 0.000 96.510 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.090 0.000 115.370 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.350 0.000 129.630 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.150 0.000 143.430 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.410 0.000 157.690 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.670 0.000 171.950 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.470 0.000 185.750 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.710 0.000 44.990 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.110 0.000 63.390 4.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.970 0.000 82.250 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.830 0.000 101.110 4.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 0.000 21.070 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 7.045 11.305 818.655 821.015 ;
      LAYER met1 ;
        RECT 1.450 0.040 818.715 821.680 ;
      LAYER met2 ;
        RECT 1.470 829.505 2.110 830.010 ;
        RECT 2.950 829.505 6.710 830.010 ;
        RECT 7.550 829.505 11.770 830.010 ;
        RECT 12.610 829.505 16.370 830.010 ;
        RECT 17.210 829.505 21.430 830.010 ;
        RECT 22.270 829.505 26.030 830.010 ;
        RECT 26.870 829.505 31.090 830.010 ;
        RECT 31.930 829.505 36.150 830.010 ;
        RECT 36.990 829.505 40.750 830.010 ;
        RECT 41.590 829.505 45.810 830.010 ;
        RECT 46.650 829.505 50.410 830.010 ;
        RECT 51.250 829.505 55.470 830.010 ;
        RECT 56.310 829.505 60.530 830.010 ;
        RECT 61.370 829.505 65.130 830.010 ;
        RECT 65.970 829.505 70.190 830.010 ;
        RECT 71.030 829.505 74.790 830.010 ;
        RECT 75.630 829.505 79.850 830.010 ;
        RECT 80.690 829.505 84.450 830.010 ;
        RECT 85.290 829.505 89.510 830.010 ;
        RECT 90.350 829.505 94.570 830.010 ;
        RECT 95.410 829.505 99.170 830.010 ;
        RECT 100.010 829.505 104.230 830.010 ;
        RECT 105.070 829.505 108.830 830.010 ;
        RECT 109.670 829.505 113.890 830.010 ;
        RECT 114.730 829.505 118.950 830.010 ;
        RECT 119.790 829.505 123.550 830.010 ;
        RECT 124.390 829.505 128.610 830.010 ;
        RECT 129.450 829.505 133.210 830.010 ;
        RECT 134.050 829.505 138.270 830.010 ;
        RECT 139.110 829.505 142.870 830.010 ;
        RECT 143.710 829.505 147.930 830.010 ;
        RECT 148.770 829.505 152.990 830.010 ;
        RECT 153.830 829.505 157.590 830.010 ;
        RECT 158.430 829.505 162.650 830.010 ;
        RECT 163.490 829.505 167.250 830.010 ;
        RECT 168.090 829.505 172.310 830.010 ;
        RECT 173.150 829.505 177.370 830.010 ;
        RECT 178.210 829.505 181.970 830.010 ;
        RECT 182.810 829.505 187.030 830.010 ;
        RECT 187.870 829.505 191.630 830.010 ;
        RECT 192.470 829.505 196.690 830.010 ;
        RECT 197.530 829.505 201.750 830.010 ;
        RECT 202.590 829.505 206.350 830.010 ;
        RECT 207.190 829.505 211.410 830.010 ;
        RECT 212.250 829.505 216.010 830.010 ;
        RECT 216.850 829.505 221.070 830.010 ;
        RECT 221.910 829.505 225.670 830.010 ;
        RECT 226.510 829.505 230.730 830.010 ;
        RECT 231.570 829.505 235.790 830.010 ;
        RECT 236.630 829.505 240.390 830.010 ;
        RECT 241.230 829.505 245.450 830.010 ;
        RECT 246.290 829.505 250.050 830.010 ;
        RECT 250.890 829.505 255.110 830.010 ;
        RECT 255.950 829.505 260.170 830.010 ;
        RECT 261.010 829.505 264.770 830.010 ;
        RECT 265.610 829.505 269.830 830.010 ;
        RECT 270.670 829.505 274.430 830.010 ;
        RECT 275.270 829.505 279.490 830.010 ;
        RECT 280.330 829.505 284.090 830.010 ;
        RECT 284.930 829.505 289.150 830.010 ;
        RECT 289.990 829.505 294.210 830.010 ;
        RECT 295.050 829.505 298.810 830.010 ;
        RECT 299.650 829.505 303.870 830.010 ;
        RECT 304.710 829.505 308.470 830.010 ;
        RECT 309.310 829.505 313.530 830.010 ;
        RECT 314.370 829.505 318.590 830.010 ;
        RECT 319.430 829.505 323.190 830.010 ;
        RECT 324.030 829.505 328.250 830.010 ;
        RECT 329.090 829.505 332.850 830.010 ;
        RECT 333.690 829.505 337.910 830.010 ;
        RECT 338.750 829.505 342.970 830.010 ;
        RECT 343.810 829.505 347.570 830.010 ;
        RECT 348.410 829.505 352.630 830.010 ;
        RECT 353.470 829.505 357.230 830.010 ;
        RECT 358.070 829.505 362.290 830.010 ;
        RECT 363.130 829.505 366.890 830.010 ;
        RECT 367.730 829.505 371.950 830.010 ;
        RECT 372.790 829.505 377.010 830.010 ;
        RECT 377.850 829.505 381.610 830.010 ;
        RECT 382.450 829.505 386.670 830.010 ;
        RECT 387.510 829.505 391.270 830.010 ;
        RECT 392.110 829.505 396.330 830.010 ;
        RECT 397.170 829.505 401.390 830.010 ;
        RECT 402.230 829.505 405.990 830.010 ;
        RECT 406.830 829.505 411.050 830.010 ;
        RECT 411.890 829.505 415.650 830.010 ;
        RECT 416.490 829.505 420.710 830.010 ;
        RECT 421.550 829.505 425.310 830.010 ;
        RECT 426.150 829.505 430.370 830.010 ;
        RECT 431.210 829.505 435.430 830.010 ;
        RECT 436.270 829.505 440.030 830.010 ;
        RECT 440.870 829.505 445.090 830.010 ;
        RECT 445.930 829.505 449.690 830.010 ;
        RECT 450.530 829.505 454.750 830.010 ;
        RECT 455.590 829.505 459.810 830.010 ;
        RECT 460.650 829.505 464.410 830.010 ;
        RECT 465.250 829.505 469.470 830.010 ;
        RECT 470.310 829.505 474.070 830.010 ;
        RECT 474.910 829.505 479.130 830.010 ;
        RECT 479.970 829.505 483.730 830.010 ;
        RECT 484.570 829.505 488.790 830.010 ;
        RECT 489.630 829.505 493.850 830.010 ;
        RECT 494.690 829.505 498.450 830.010 ;
        RECT 499.290 829.505 503.510 830.010 ;
        RECT 504.350 829.505 508.110 830.010 ;
        RECT 508.950 829.505 513.170 830.010 ;
        RECT 514.010 829.505 518.230 830.010 ;
        RECT 519.070 829.505 522.830 830.010 ;
        RECT 523.670 829.505 527.890 830.010 ;
        RECT 528.730 829.505 532.490 830.010 ;
        RECT 533.330 829.505 537.550 830.010 ;
        RECT 538.390 829.505 542.610 830.010 ;
        RECT 543.450 829.505 547.210 830.010 ;
        RECT 548.050 829.505 552.270 830.010 ;
        RECT 553.110 829.505 556.870 830.010 ;
        RECT 557.710 829.505 561.930 830.010 ;
        RECT 562.770 829.505 566.530 830.010 ;
        RECT 567.370 829.505 571.590 830.010 ;
        RECT 572.430 829.505 576.650 830.010 ;
        RECT 577.490 829.505 581.250 830.010 ;
        RECT 582.090 829.505 586.310 830.010 ;
        RECT 587.150 829.505 590.910 830.010 ;
        RECT 591.750 829.505 595.970 830.010 ;
        RECT 596.810 829.505 601.030 830.010 ;
        RECT 601.870 829.505 605.630 830.010 ;
        RECT 606.470 829.505 610.690 830.010 ;
        RECT 611.530 829.505 615.290 830.010 ;
        RECT 616.130 829.505 620.350 830.010 ;
        RECT 621.190 829.505 624.950 830.010 ;
        RECT 625.790 829.505 630.010 830.010 ;
        RECT 630.850 829.505 635.070 830.010 ;
        RECT 635.910 829.505 639.670 830.010 ;
        RECT 640.510 829.505 644.730 830.010 ;
        RECT 645.570 829.505 649.330 830.010 ;
        RECT 650.170 829.505 654.390 830.010 ;
        RECT 655.230 829.505 659.450 830.010 ;
        RECT 660.290 829.505 664.050 830.010 ;
        RECT 664.890 829.505 669.110 830.010 ;
        RECT 669.950 829.505 673.710 830.010 ;
        RECT 674.550 829.505 678.770 830.010 ;
        RECT 679.610 829.505 683.830 830.010 ;
        RECT 684.670 829.505 688.430 830.010 ;
        RECT 689.270 829.505 693.490 830.010 ;
        RECT 694.330 829.505 698.090 830.010 ;
        RECT 698.930 829.505 703.150 830.010 ;
        RECT 703.990 829.505 707.750 830.010 ;
        RECT 708.590 829.505 712.810 830.010 ;
        RECT 713.650 829.505 717.870 830.010 ;
        RECT 718.710 829.505 722.470 830.010 ;
        RECT 723.310 829.505 727.530 830.010 ;
        RECT 728.370 829.505 732.130 830.010 ;
        RECT 732.970 829.505 737.190 830.010 ;
        RECT 738.030 829.505 742.250 830.010 ;
        RECT 743.090 829.505 746.850 830.010 ;
        RECT 747.690 829.505 751.910 830.010 ;
        RECT 752.750 829.505 756.510 830.010 ;
        RECT 757.350 829.505 761.570 830.010 ;
        RECT 762.410 829.505 766.170 830.010 ;
        RECT 767.010 829.505 771.230 830.010 ;
        RECT 772.070 829.505 776.290 830.010 ;
        RECT 777.130 829.505 780.890 830.010 ;
        RECT 781.730 829.505 785.950 830.010 ;
        RECT 786.790 829.505 790.550 830.010 ;
        RECT 791.390 829.505 795.610 830.010 ;
        RECT 796.450 829.505 800.670 830.010 ;
        RECT 801.510 829.505 805.270 830.010 ;
        RECT 806.110 829.505 810.330 830.010 ;
        RECT 811.170 829.505 814.930 830.010 ;
        RECT 1.470 4.280 815.030 829.505 ;
        RECT 1.470 0.010 2.110 4.280 ;
        RECT 2.950 0.010 6.710 4.280 ;
        RECT 7.550 0.010 11.310 4.280 ;
        RECT 12.150 0.010 15.910 4.280 ;
        RECT 16.750 0.010 20.510 4.280 ;
        RECT 21.350 0.010 25.570 4.280 ;
        RECT 26.410 0.010 30.170 4.280 ;
        RECT 31.010 0.010 34.770 4.280 ;
        RECT 35.610 0.010 39.370 4.280 ;
        RECT 40.210 0.010 44.430 4.280 ;
        RECT 45.270 0.010 49.030 4.280 ;
        RECT 49.870 0.010 53.630 4.280 ;
        RECT 54.470 0.010 58.230 4.280 ;
        RECT 59.070 0.010 62.830 4.280 ;
        RECT 63.670 0.010 67.890 4.280 ;
        RECT 68.730 0.010 72.490 4.280 ;
        RECT 73.330 0.010 77.090 4.280 ;
        RECT 77.930 0.010 81.690 4.280 ;
        RECT 82.530 0.010 86.750 4.280 ;
        RECT 87.590 0.010 91.350 4.280 ;
        RECT 92.190 0.010 95.950 4.280 ;
        RECT 96.790 0.010 100.550 4.280 ;
        RECT 101.390 0.010 105.150 4.280 ;
        RECT 105.990 0.010 110.210 4.280 ;
        RECT 111.050 0.010 114.810 4.280 ;
        RECT 115.650 0.010 119.410 4.280 ;
        RECT 120.250 0.010 124.010 4.280 ;
        RECT 124.850 0.010 129.070 4.280 ;
        RECT 129.910 0.010 133.670 4.280 ;
        RECT 134.510 0.010 138.270 4.280 ;
        RECT 139.110 0.010 142.870 4.280 ;
        RECT 143.710 0.010 147.470 4.280 ;
        RECT 148.310 0.010 152.530 4.280 ;
        RECT 153.370 0.010 157.130 4.280 ;
        RECT 157.970 0.010 161.730 4.280 ;
        RECT 162.570 0.010 166.330 4.280 ;
        RECT 167.170 0.010 171.390 4.280 ;
        RECT 172.230 0.010 175.990 4.280 ;
        RECT 176.830 0.010 180.590 4.280 ;
        RECT 181.430 0.010 185.190 4.280 ;
        RECT 186.030 0.010 189.790 4.280 ;
        RECT 190.630 0.010 194.850 4.280 ;
        RECT 195.690 0.010 199.450 4.280 ;
        RECT 200.290 0.010 204.050 4.280 ;
        RECT 204.890 0.010 208.650 4.280 ;
        RECT 209.490 0.010 213.710 4.280 ;
        RECT 214.550 0.010 218.310 4.280 ;
        RECT 219.150 0.010 222.910 4.280 ;
        RECT 223.750 0.010 227.510 4.280 ;
        RECT 228.350 0.010 232.110 4.280 ;
        RECT 232.950 0.010 237.170 4.280 ;
        RECT 238.010 0.010 241.770 4.280 ;
        RECT 242.610 0.010 246.370 4.280 ;
        RECT 247.210 0.010 250.970 4.280 ;
        RECT 251.810 0.010 256.030 4.280 ;
        RECT 256.870 0.010 260.630 4.280 ;
        RECT 261.470 0.010 265.230 4.280 ;
        RECT 266.070 0.010 269.830 4.280 ;
        RECT 270.670 0.010 274.430 4.280 ;
        RECT 275.270 0.010 279.490 4.280 ;
        RECT 280.330 0.010 284.090 4.280 ;
        RECT 284.930 0.010 288.690 4.280 ;
        RECT 289.530 0.010 293.290 4.280 ;
        RECT 294.130 0.010 298.350 4.280 ;
        RECT 299.190 0.010 302.950 4.280 ;
        RECT 303.790 0.010 307.550 4.280 ;
        RECT 308.390 0.010 312.150 4.280 ;
        RECT 312.990 0.010 316.750 4.280 ;
        RECT 317.590 0.010 321.810 4.280 ;
        RECT 322.650 0.010 326.410 4.280 ;
        RECT 327.250 0.010 331.010 4.280 ;
        RECT 331.850 0.010 335.610 4.280 ;
        RECT 336.450 0.010 340.670 4.280 ;
        RECT 341.510 0.010 345.270 4.280 ;
        RECT 346.110 0.010 349.870 4.280 ;
        RECT 350.710 0.010 354.470 4.280 ;
        RECT 355.310 0.010 359.070 4.280 ;
        RECT 359.910 0.010 364.130 4.280 ;
        RECT 364.970 0.010 368.730 4.280 ;
        RECT 369.570 0.010 373.330 4.280 ;
        RECT 374.170 0.010 377.930 4.280 ;
        RECT 378.770 0.010 382.990 4.280 ;
        RECT 383.830 0.010 387.590 4.280 ;
        RECT 388.430 0.010 392.190 4.280 ;
        RECT 393.030 0.010 396.790 4.280 ;
        RECT 397.630 0.010 401.390 4.280 ;
        RECT 402.230 0.010 406.450 4.280 ;
        RECT 407.290 0.010 411.050 4.280 ;
        RECT 411.890 0.010 415.650 4.280 ;
        RECT 416.490 0.010 420.250 4.280 ;
        RECT 421.090 0.010 425.310 4.280 ;
        RECT 426.150 0.010 429.910 4.280 ;
        RECT 430.750 0.010 434.510 4.280 ;
        RECT 435.350 0.010 439.110 4.280 ;
        RECT 439.950 0.010 443.710 4.280 ;
        RECT 444.550 0.010 448.770 4.280 ;
        RECT 449.610 0.010 453.370 4.280 ;
        RECT 454.210 0.010 457.970 4.280 ;
        RECT 458.810 0.010 462.570 4.280 ;
        RECT 463.410 0.010 467.630 4.280 ;
        RECT 468.470 0.010 472.230 4.280 ;
        RECT 473.070 0.010 476.830 4.280 ;
        RECT 477.670 0.010 481.430 4.280 ;
        RECT 482.270 0.010 486.030 4.280 ;
        RECT 486.870 0.010 491.090 4.280 ;
        RECT 491.930 0.010 495.690 4.280 ;
        RECT 496.530 0.010 500.290 4.280 ;
        RECT 501.130 0.010 504.890 4.280 ;
        RECT 505.730 0.010 509.950 4.280 ;
        RECT 510.790 0.010 514.550 4.280 ;
        RECT 515.390 0.010 519.150 4.280 ;
        RECT 519.990 0.010 523.750 4.280 ;
        RECT 524.590 0.010 528.350 4.280 ;
        RECT 529.190 0.010 533.410 4.280 ;
        RECT 534.250 0.010 538.010 4.280 ;
        RECT 538.850 0.010 542.610 4.280 ;
        RECT 543.450 0.010 547.210 4.280 ;
        RECT 548.050 0.010 552.270 4.280 ;
        RECT 553.110 0.010 556.870 4.280 ;
        RECT 557.710 0.010 561.470 4.280 ;
        RECT 562.310 0.010 566.070 4.280 ;
        RECT 566.910 0.010 570.670 4.280 ;
        RECT 571.510 0.010 575.730 4.280 ;
        RECT 576.570 0.010 580.330 4.280 ;
        RECT 581.170 0.010 584.930 4.280 ;
        RECT 585.770 0.010 589.530 4.280 ;
        RECT 590.370 0.010 594.590 4.280 ;
        RECT 595.430 0.010 599.190 4.280 ;
        RECT 600.030 0.010 603.790 4.280 ;
        RECT 604.630 0.010 608.390 4.280 ;
        RECT 609.230 0.010 612.990 4.280 ;
        RECT 613.830 0.010 618.050 4.280 ;
        RECT 618.890 0.010 622.650 4.280 ;
        RECT 623.490 0.010 627.250 4.280 ;
        RECT 628.090 0.010 631.850 4.280 ;
        RECT 632.690 0.010 636.910 4.280 ;
        RECT 637.750 0.010 641.510 4.280 ;
        RECT 642.350 0.010 646.110 4.280 ;
        RECT 646.950 0.010 650.710 4.280 ;
        RECT 651.550 0.010 655.310 4.280 ;
        RECT 656.150 0.010 660.370 4.280 ;
        RECT 661.210 0.010 664.970 4.280 ;
        RECT 665.810 0.010 669.570 4.280 ;
        RECT 670.410 0.010 674.170 4.280 ;
        RECT 675.010 0.010 679.230 4.280 ;
        RECT 680.070 0.010 683.830 4.280 ;
        RECT 684.670 0.010 688.430 4.280 ;
        RECT 689.270 0.010 693.030 4.280 ;
        RECT 693.870 0.010 697.630 4.280 ;
        RECT 698.470 0.010 702.690 4.280 ;
        RECT 703.530 0.010 707.290 4.280 ;
        RECT 708.130 0.010 711.890 4.280 ;
        RECT 712.730 0.010 716.490 4.280 ;
        RECT 717.330 0.010 721.550 4.280 ;
        RECT 722.390 0.010 726.150 4.280 ;
        RECT 726.990 0.010 730.750 4.280 ;
        RECT 731.590 0.010 735.350 4.280 ;
        RECT 736.190 0.010 739.950 4.280 ;
        RECT 740.790 0.010 745.010 4.280 ;
        RECT 745.850 0.010 749.610 4.280 ;
        RECT 750.450 0.010 754.210 4.280 ;
        RECT 755.050 0.010 758.810 4.280 ;
        RECT 759.650 0.010 763.870 4.280 ;
        RECT 764.710 0.010 768.470 4.280 ;
        RECT 769.310 0.010 773.070 4.280 ;
        RECT 773.910 0.010 777.670 4.280 ;
        RECT 778.510 0.010 782.270 4.280 ;
        RECT 783.110 0.010 787.330 4.280 ;
        RECT 788.170 0.010 791.930 4.280 ;
        RECT 792.770 0.010 796.530 4.280 ;
        RECT 797.370 0.010 801.130 4.280 ;
        RECT 801.970 0.010 806.190 4.280 ;
        RECT 807.030 0.010 810.790 4.280 ;
        RECT 811.630 0.010 815.030 4.280 ;
      LAYER met3 ;
        RECT 4.400 825.840 818.665 826.705 ;
        RECT 1.190 813.640 819.065 825.840 ;
        RECT 1.190 812.960 818.665 813.640 ;
        RECT 4.400 812.240 818.665 812.960 ;
        RECT 4.400 811.560 819.065 812.240 ;
        RECT 1.190 800.040 819.065 811.560 ;
        RECT 1.190 798.680 818.665 800.040 ;
        RECT 4.400 798.640 818.665 798.680 ;
        RECT 4.400 797.280 819.065 798.640 ;
        RECT 1.190 786.440 819.065 797.280 ;
        RECT 1.190 785.040 818.665 786.440 ;
        RECT 1.190 784.400 819.065 785.040 ;
        RECT 4.400 783.000 819.065 784.400 ;
        RECT 1.190 773.520 819.065 783.000 ;
        RECT 1.190 772.120 818.665 773.520 ;
        RECT 1.190 770.800 819.065 772.120 ;
        RECT 4.400 769.400 819.065 770.800 ;
        RECT 1.190 759.920 819.065 769.400 ;
        RECT 1.190 758.520 818.665 759.920 ;
        RECT 1.190 756.520 819.065 758.520 ;
        RECT 4.400 755.120 819.065 756.520 ;
        RECT 1.190 746.320 819.065 755.120 ;
        RECT 1.190 744.920 818.665 746.320 ;
        RECT 1.190 742.240 819.065 744.920 ;
        RECT 4.400 740.840 819.065 742.240 ;
        RECT 1.190 732.720 819.065 740.840 ;
        RECT 1.190 731.320 818.665 732.720 ;
        RECT 1.190 727.960 819.065 731.320 ;
        RECT 4.400 726.560 819.065 727.960 ;
        RECT 1.190 719.800 819.065 726.560 ;
        RECT 1.190 718.400 818.665 719.800 ;
        RECT 1.190 713.680 819.065 718.400 ;
        RECT 4.400 712.280 819.065 713.680 ;
        RECT 1.190 706.200 819.065 712.280 ;
        RECT 1.190 704.800 818.665 706.200 ;
        RECT 1.190 700.080 819.065 704.800 ;
        RECT 4.400 698.680 819.065 700.080 ;
        RECT 1.190 692.600 819.065 698.680 ;
        RECT 1.190 691.200 818.665 692.600 ;
        RECT 1.190 685.800 819.065 691.200 ;
        RECT 4.400 684.400 819.065 685.800 ;
        RECT 1.190 679.000 819.065 684.400 ;
        RECT 1.190 677.600 818.665 679.000 ;
        RECT 1.190 671.520 819.065 677.600 ;
        RECT 4.400 670.120 819.065 671.520 ;
        RECT 1.190 665.400 819.065 670.120 ;
        RECT 1.190 664.000 818.665 665.400 ;
        RECT 1.190 657.240 819.065 664.000 ;
        RECT 4.400 655.840 819.065 657.240 ;
        RECT 1.190 652.480 819.065 655.840 ;
        RECT 1.190 651.080 818.665 652.480 ;
        RECT 1.190 643.640 819.065 651.080 ;
        RECT 4.400 642.240 819.065 643.640 ;
        RECT 1.190 638.880 819.065 642.240 ;
        RECT 1.190 637.480 818.665 638.880 ;
        RECT 1.190 629.360 819.065 637.480 ;
        RECT 4.400 627.960 819.065 629.360 ;
        RECT 1.190 625.280 819.065 627.960 ;
        RECT 1.190 623.880 818.665 625.280 ;
        RECT 1.190 615.080 819.065 623.880 ;
        RECT 4.400 613.680 819.065 615.080 ;
        RECT 1.190 611.680 819.065 613.680 ;
        RECT 1.190 610.280 818.665 611.680 ;
        RECT 1.190 600.800 819.065 610.280 ;
        RECT 4.400 599.400 819.065 600.800 ;
        RECT 1.190 598.760 819.065 599.400 ;
        RECT 1.190 597.360 818.665 598.760 ;
        RECT 1.190 586.520 819.065 597.360 ;
        RECT 4.400 585.160 819.065 586.520 ;
        RECT 4.400 585.120 818.665 585.160 ;
        RECT 1.190 583.760 818.665 585.120 ;
        RECT 1.190 572.920 819.065 583.760 ;
        RECT 4.400 571.560 819.065 572.920 ;
        RECT 4.400 571.520 818.665 571.560 ;
        RECT 1.190 570.160 818.665 571.520 ;
        RECT 1.190 558.640 819.065 570.160 ;
        RECT 4.400 557.960 819.065 558.640 ;
        RECT 4.400 557.240 818.665 557.960 ;
        RECT 1.190 556.560 818.665 557.240 ;
        RECT 1.190 544.360 819.065 556.560 ;
        RECT 4.400 542.960 818.665 544.360 ;
        RECT 1.190 531.440 819.065 542.960 ;
        RECT 1.190 530.080 818.665 531.440 ;
        RECT 4.400 530.040 818.665 530.080 ;
        RECT 4.400 528.680 819.065 530.040 ;
        RECT 1.190 517.840 819.065 528.680 ;
        RECT 1.190 516.480 818.665 517.840 ;
        RECT 4.400 516.440 818.665 516.480 ;
        RECT 4.400 515.080 819.065 516.440 ;
        RECT 1.190 504.240 819.065 515.080 ;
        RECT 1.190 502.840 818.665 504.240 ;
        RECT 1.190 502.200 819.065 502.840 ;
        RECT 4.400 500.800 819.065 502.200 ;
        RECT 1.190 490.640 819.065 500.800 ;
        RECT 1.190 489.240 818.665 490.640 ;
        RECT 1.190 487.920 819.065 489.240 ;
        RECT 4.400 486.520 819.065 487.920 ;
        RECT 1.190 477.720 819.065 486.520 ;
        RECT 1.190 476.320 818.665 477.720 ;
        RECT 1.190 473.640 819.065 476.320 ;
        RECT 4.400 472.240 819.065 473.640 ;
        RECT 1.190 464.120 819.065 472.240 ;
        RECT 1.190 462.720 818.665 464.120 ;
        RECT 1.190 459.360 819.065 462.720 ;
        RECT 4.400 457.960 819.065 459.360 ;
        RECT 1.190 450.520 819.065 457.960 ;
        RECT 1.190 449.120 818.665 450.520 ;
        RECT 1.190 445.760 819.065 449.120 ;
        RECT 4.400 444.360 819.065 445.760 ;
        RECT 1.190 436.920 819.065 444.360 ;
        RECT 1.190 435.520 818.665 436.920 ;
        RECT 1.190 431.480 819.065 435.520 ;
        RECT 4.400 430.080 819.065 431.480 ;
        RECT 1.190 424.000 819.065 430.080 ;
        RECT 1.190 422.600 818.665 424.000 ;
        RECT 1.190 417.200 819.065 422.600 ;
        RECT 4.400 415.800 819.065 417.200 ;
        RECT 1.190 410.400 819.065 415.800 ;
        RECT 1.190 409.000 818.665 410.400 ;
        RECT 1.190 402.920 819.065 409.000 ;
        RECT 4.400 401.520 819.065 402.920 ;
        RECT 1.190 396.800 819.065 401.520 ;
        RECT 1.190 395.400 818.665 396.800 ;
        RECT 1.190 389.320 819.065 395.400 ;
        RECT 4.400 387.920 819.065 389.320 ;
        RECT 1.190 383.200 819.065 387.920 ;
        RECT 1.190 381.800 818.665 383.200 ;
        RECT 1.190 375.040 819.065 381.800 ;
        RECT 4.400 373.640 819.065 375.040 ;
        RECT 1.190 369.600 819.065 373.640 ;
        RECT 1.190 368.200 818.665 369.600 ;
        RECT 1.190 360.760 819.065 368.200 ;
        RECT 4.400 359.360 819.065 360.760 ;
        RECT 1.190 356.680 819.065 359.360 ;
        RECT 1.190 355.280 818.665 356.680 ;
        RECT 1.190 346.480 819.065 355.280 ;
        RECT 4.400 345.080 819.065 346.480 ;
        RECT 1.190 343.080 819.065 345.080 ;
        RECT 1.190 341.680 818.665 343.080 ;
        RECT 1.190 332.200 819.065 341.680 ;
        RECT 4.400 330.800 819.065 332.200 ;
        RECT 1.190 329.480 819.065 330.800 ;
        RECT 1.190 328.080 818.665 329.480 ;
        RECT 1.190 318.600 819.065 328.080 ;
        RECT 4.400 317.200 819.065 318.600 ;
        RECT 1.190 315.880 819.065 317.200 ;
        RECT 1.190 314.480 818.665 315.880 ;
        RECT 1.190 304.320 819.065 314.480 ;
        RECT 4.400 302.960 819.065 304.320 ;
        RECT 4.400 302.920 818.665 302.960 ;
        RECT 1.190 301.560 818.665 302.920 ;
        RECT 1.190 290.040 819.065 301.560 ;
        RECT 4.400 289.360 819.065 290.040 ;
        RECT 4.400 288.640 818.665 289.360 ;
        RECT 1.190 287.960 818.665 288.640 ;
        RECT 1.190 275.760 819.065 287.960 ;
        RECT 4.400 274.360 818.665 275.760 ;
        RECT 1.190 262.160 819.065 274.360 ;
        RECT 4.400 260.760 818.665 262.160 ;
        RECT 1.190 248.560 819.065 260.760 ;
        RECT 1.190 247.880 818.665 248.560 ;
        RECT 4.400 247.160 818.665 247.880 ;
        RECT 4.400 246.480 819.065 247.160 ;
        RECT 1.190 235.640 819.065 246.480 ;
        RECT 1.190 234.240 818.665 235.640 ;
        RECT 1.190 233.600 819.065 234.240 ;
        RECT 4.400 232.200 819.065 233.600 ;
        RECT 1.190 222.040 819.065 232.200 ;
        RECT 1.190 220.640 818.665 222.040 ;
        RECT 1.190 219.320 819.065 220.640 ;
        RECT 4.400 217.920 819.065 219.320 ;
        RECT 1.190 208.440 819.065 217.920 ;
        RECT 1.190 207.040 818.665 208.440 ;
        RECT 1.190 205.040 819.065 207.040 ;
        RECT 4.400 203.640 819.065 205.040 ;
        RECT 1.190 194.840 819.065 203.640 ;
        RECT 1.190 193.440 818.665 194.840 ;
        RECT 1.190 191.440 819.065 193.440 ;
        RECT 4.400 190.040 819.065 191.440 ;
        RECT 1.190 181.920 819.065 190.040 ;
        RECT 1.190 180.520 818.665 181.920 ;
        RECT 1.190 177.160 819.065 180.520 ;
        RECT 4.400 175.760 819.065 177.160 ;
        RECT 1.190 168.320 819.065 175.760 ;
        RECT 1.190 166.920 818.665 168.320 ;
        RECT 1.190 162.880 819.065 166.920 ;
        RECT 4.400 161.480 819.065 162.880 ;
        RECT 1.190 154.720 819.065 161.480 ;
        RECT 1.190 153.320 818.665 154.720 ;
        RECT 1.190 148.600 819.065 153.320 ;
        RECT 4.400 147.200 819.065 148.600 ;
        RECT 1.190 141.120 819.065 147.200 ;
        RECT 1.190 139.720 818.665 141.120 ;
        RECT 1.190 135.000 819.065 139.720 ;
        RECT 4.400 133.600 819.065 135.000 ;
        RECT 1.190 127.520 819.065 133.600 ;
        RECT 1.190 126.120 818.665 127.520 ;
        RECT 1.190 120.720 819.065 126.120 ;
        RECT 4.400 119.320 819.065 120.720 ;
        RECT 1.190 114.600 819.065 119.320 ;
        RECT 1.190 113.200 818.665 114.600 ;
        RECT 1.190 106.440 819.065 113.200 ;
        RECT 4.400 105.040 819.065 106.440 ;
        RECT 1.190 101.000 819.065 105.040 ;
        RECT 1.190 99.600 818.665 101.000 ;
        RECT 1.190 92.160 819.065 99.600 ;
        RECT 4.400 90.760 819.065 92.160 ;
        RECT 1.190 87.400 819.065 90.760 ;
        RECT 1.190 86.000 818.665 87.400 ;
        RECT 1.190 77.880 819.065 86.000 ;
        RECT 4.400 76.480 819.065 77.880 ;
        RECT 1.190 73.800 819.065 76.480 ;
        RECT 1.190 72.400 818.665 73.800 ;
        RECT 1.190 64.280 819.065 72.400 ;
        RECT 4.400 62.880 819.065 64.280 ;
        RECT 1.190 60.880 819.065 62.880 ;
        RECT 1.190 59.480 818.665 60.880 ;
        RECT 1.190 50.000 819.065 59.480 ;
        RECT 4.400 48.600 819.065 50.000 ;
        RECT 1.190 47.280 819.065 48.600 ;
        RECT 1.190 45.880 818.665 47.280 ;
        RECT 1.190 35.720 819.065 45.880 ;
        RECT 4.400 34.320 819.065 35.720 ;
        RECT 1.190 33.680 819.065 34.320 ;
        RECT 1.190 32.280 818.665 33.680 ;
        RECT 1.190 21.440 819.065 32.280 ;
        RECT 4.400 20.080 819.065 21.440 ;
        RECT 4.400 20.040 818.665 20.080 ;
        RECT 1.190 18.680 818.665 20.040 ;
        RECT 1.190 7.840 819.065 18.680 ;
        RECT 4.400 7.160 819.065 7.840 ;
        RECT 4.400 6.440 818.665 7.160 ;
        RECT 1.190 5.760 818.665 6.440 ;
        RECT 1.190 0.175 819.065 5.760 ;
      LAYER met4 ;
        RECT 1.215 10.240 20.640 820.585 ;
        RECT 23.040 10.240 97.440 820.585 ;
        RECT 99.840 10.240 174.240 820.585 ;
        RECT 176.640 10.240 251.040 820.585 ;
        RECT 253.440 10.240 327.840 820.585 ;
        RECT 330.240 10.240 404.640 820.585 ;
        RECT 407.040 10.240 481.440 820.585 ;
        RECT 483.840 10.240 558.240 820.585 ;
        RECT 560.640 10.240 635.040 820.585 ;
        RECT 637.440 10.240 705.345 820.585 ;
        RECT 1.215 2.215 705.345 10.240 ;
  END
END user_proj
END LIBRARY

