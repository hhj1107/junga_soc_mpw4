VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_proj
  CLASS BLOCK ;
  FOREIGN user_proj ;
  ORIGIN 0.000 0.000 ;
  SIZE 823.900 BY 834.620 ;
  PIN i_dout0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.610 830.620 534.890 834.620 ;
    END
  END i_dout0[0]
  PIN i_dout0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.070 830.620 627.350 834.620 ;
    END
  END i_dout0[10]
  PIN i_dout0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 384.920 4.000 385.520 ;
    END
  END i_dout0[11]
  PIN i_dout0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 645.470 830.620 645.750 834.620 ;
    END
  END i_dout0[12]
  PIN i_dout0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 459.720 823.900 460.320 ;
    END
  END i_dout0[13]
  PIN i_dout0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 797.270 0.000 797.550 4.000 ;
    END
  END i_dout0[14]
  PIN i_dout0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 520.920 823.900 521.520 ;
    END
  END i_dout0[15]
  PIN i_dout0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 801.870 0.000 802.150 4.000 ;
    END
  END i_dout0[16]
  PIN i_dout0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 545.400 823.900 546.000 ;
    END
  END i_dout0[17]
  PIN i_dout0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 696.530 830.620 696.810 834.620 ;
    END
  END i_dout0[18]
  PIN i_dout0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 595.040 823.900 595.640 ;
    END
  END i_dout0[19]
  PIN i_dout0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 42.880 823.900 43.480 ;
    END
  END i_dout0[1]
  PIN i_dout0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 710.330 830.620 710.610 834.620 ;
    END
  END i_dout0[20]
  PIN i_dout0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 631.760 823.900 632.360 ;
    END
  END i_dout0[21]
  PIN i_dout0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 719.530 830.620 719.810 834.620 ;
    END
  END i_dout0[22]
  PIN i_dout0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 620.880 4.000 621.480 ;
    END
  END i_dout0[23]
  PIN i_dout0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 756.790 830.620 757.070 834.620 ;
    END
  END i_dout0[24]
  PIN i_dout0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 765.990 830.620 766.270 834.620 ;
    END
  END i_dout0[25]
  PIN i_dout0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 754.160 823.900 754.760 ;
    END
  END i_dout0[26]
  PIN i_dout0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 731.040 4.000 731.640 ;
    END
  END i_dout0[27]
  PIN i_dout0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 766.400 823.900 767.000 ;
    END
  END i_dout0[28]
  PIN i_dout0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 788.990 830.620 789.270 834.620 ;
    END
  END i_dout0[29]
  PIN i_dout0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.680 4.000 118.280 ;
    END
  END i_dout0[2]
  PIN i_dout0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 798.190 830.620 798.470 834.620 ;
    END
  END i_dout0[30]
  PIN i_dout0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 821.190 830.620 821.470 834.620 ;
    END
  END i_dout0[31]
  PIN i_dout0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 759.550 0.000 759.830 4.000 ;
    END
  END i_dout0[3]
  PIN i_dout0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 226.480 823.900 227.080 ;
    END
  END i_dout0[4]
  PIN i_dout0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 263.200 823.900 263.800 ;
    END
  END i_dout0[5]
  PIN i_dout0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 243.480 4.000 244.080 ;
    END
  END i_dout0[6]
  PIN i_dout0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 776.110 0.000 776.390 4.000 ;
    END
  END i_dout0[7]
  PIN i_dout0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 306.040 4.000 306.640 ;
    END
  END i_dout0[8]
  PIN i_dout0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 786.690 0.000 786.970 4.000 ;
    END
  END i_dout0[9]
  PIN i_dout0_1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 741.610 0.000 741.890 4.000 ;
    END
  END i_dout0_1[0]
  PIN i_dout0_1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 398.520 823.900 399.120 ;
    END
  END i_dout0_1[10]
  PIN i_dout0_1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 369.280 4.000 369.880 ;
    END
  END i_dout0_1[11]
  PIN i_dout0_1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 794.050 0.000 794.330 4.000 ;
    END
  END i_dout0_1[12]
  PIN i_dout0_1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 447.480 823.900 448.080 ;
    END
  END i_dout0_1[13]
  PIN i_dout0_1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.070 830.620 650.350 834.620 ;
    END
  END i_dout0_1[14]
  PIN i_dout0_1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 663.870 830.620 664.150 834.620 ;
    END
  END i_dout0_1[15]
  PIN i_dout0_1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.070 830.620 673.350 834.620 ;
    END
  END i_dout0_1[16]
  PIN i_dout0_1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 526.360 4.000 526.960 ;
    END
  END i_dout0_1[17]
  PIN i_dout0_1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 687.330 830.620 687.610 834.620 ;
    END
  END i_dout0_1[18]
  PIN i_dout0_1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 570.560 823.900 571.160 ;
    END
  END i_dout0_1[19]
  PIN i_dout0_1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.010 830.620 553.290 834.620 ;
    END
  END i_dout0_1[1]
  PIN i_dout0_1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 573.960 4.000 574.560 ;
    END
  END i_dout0_1[20]
  PIN i_dout0_1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 809.230 0.000 809.510 4.000 ;
    END
  END i_dout0_1[21]
  PIN i_dout0_1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 810.610 0.000 810.890 4.000 ;
    END
  END i_dout0_1[22]
  PIN i_dout0_1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.930 830.620 738.210 834.620 ;
    END
  END i_dout0_1[23]
  PIN i_dout0_1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 752.190 830.620 752.470 834.620 ;
    END
  END i_dout0_1[24]
  PIN i_dout0_1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 729.680 823.900 730.280 ;
    END
  END i_dout0_1[25]
  PIN i_dout0_1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 684.120 4.000 684.720 ;
    END
  END i_dout0_1[26]
  PIN i_dout0_1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 816.590 0.000 816.870 4.000 ;
    END
  END i_dout0_1[27]
  PIN i_dout0_1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 763.000 4.000 763.600 ;
    END
  END i_dout0_1[28]
  PIN i_dout0_1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 778.640 4.000 779.240 ;
    END
  END i_dout0_1[29]
  PIN i_dout0_1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 566.810 830.620 567.090 834.620 ;
    END
  END i_dout0_1[2]
  PIN i_dout0_1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 794.280 4.000 794.880 ;
    END
  END i_dout0_1[30]
  PIN i_dout0_1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 811.990 830.620 812.270 834.620 ;
    END
  END i_dout0_1[31]
  PIN i_dout0_1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 758.170 0.000 758.450 4.000 ;
    END
  END i_dout0_1[3]
  PIN i_dout0_1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 214.240 823.900 214.840 ;
    END
  END i_dout0_1[4]
  PIN i_dout0_1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 765.990 0.000 766.270 4.000 ;
    END
  END i_dout0_1[5]
  PIN i_dout0_1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 768.750 0.000 769.030 4.000 ;
    END
  END i_dout0_1[6]
  PIN i_dout0_1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 774.730 0.000 775.010 4.000 ;
    END
  END i_dout0_1[7]
  PIN i_dout0_1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 617.870 830.620 618.150 834.620 ;
    END
  END i_dout0_1[8]
  PIN i_dout0_1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 322.360 4.000 322.960 ;
    END
  END i_dout0_1[9]
  PIN i_dout1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 7.520 4.000 8.120 ;
    END
  END i_dout1[0]
  PIN i_dout1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 631.670 830.620 631.950 834.620 ;
    END
  END i_dout1[10]
  PIN i_dout1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 791.290 0.000 791.570 4.000 ;
    END
  END i_dout1[11]
  PIN i_dout1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 423.000 823.900 423.600 ;
    END
  END i_dout1[12]
  PIN i_dout1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 471.960 823.900 472.560 ;
    END
  END i_dout1[13]
  PIN i_dout1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 654.670 830.620 654.950 834.620 ;
    END
  END i_dout1[14]
  PIN i_dout1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 463.800 4.000 464.400 ;
    END
  END i_dout1[15]
  PIN i_dout1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 495.080 4.000 495.680 ;
    END
  END i_dout1[16]
  PIN i_dout1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 557.640 823.900 558.240 ;
    END
  END i_dout1[17]
  PIN i_dout1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 542.680 4.000 543.280 ;
    END
  END i_dout1[18]
  PIN i_dout1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 607.280 823.900 607.880 ;
    END
  END i_dout1[19]
  PIN i_dout1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 67.360 823.900 67.960 ;
    END
  END i_dout1[1]
  PIN i_dout1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 605.240 4.000 605.840 ;
    END
  END i_dout1[20]
  PIN i_dout1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 644.000 823.900 644.600 ;
    END
  END i_dout1[21]
  PIN i_dout1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 724.130 830.620 724.410 834.620 ;
    END
  END i_dout1[22]
  PIN i_dout1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 680.720 823.900 681.320 ;
    END
  END i_dout1[23]
  PIN i_dout1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 761.390 830.620 761.670 834.620 ;
    END
  END i_dout1[24]
  PIN i_dout1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 668.480 4.000 669.080 ;
    END
  END i_dout1[25]
  PIN i_dout1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 699.760 4.000 700.360 ;
    END
  END i_dout1[26]
  PIN i_dout1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 775.190 830.620 775.470 834.620 ;
    END
  END i_dout1[27]
  PIN i_dout1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 778.640 823.900 779.240 ;
    END
  END i_dout1[28]
  PIN i_dout1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 821.190 0.000 821.470 4.000 ;
    END
  END i_dout1[29]
  PIN i_dout1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 104.080 823.900 104.680 ;
    END
  END i_dout1[2]
  PIN i_dout1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 802.790 830.620 803.070 834.620 ;
    END
  END i_dout1[30]
  PIN i_dout1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 809.920 4.000 810.520 ;
    END
  END i_dout1[31]
  PIN i_dout1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 571.410 830.620 571.690 834.620 ;
    END
  END i_dout1[3]
  PIN i_dout1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 238.720 823.900 239.320 ;
    END
  END i_dout1[4]
  PIN i_dout1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 275.440 823.900 276.040 ;
    END
  END i_dout1[5]
  PIN i_dout1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.010 830.620 599.290 834.620 ;
    END
  END i_dout1[6]
  PIN i_dout1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 259.120 4.000 259.720 ;
    END
  END i_dout1[7]
  PIN i_dout1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 780.710 0.000 780.990 4.000 ;
    END
  END i_dout1[8]
  PIN i_dout1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 353.640 4.000 354.240 ;
    END
  END i_dout1[9]
  PIN i_dout1_1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 743.450 0.000 743.730 4.000 ;
    END
  END i_dout1_1[0]
  PIN i_dout1_1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 410.760 823.900 411.360 ;
    END
  END i_dout1_1[10]
  PIN i_dout1_1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 640.870 830.620 641.150 834.620 ;
    END
  END i_dout1_1[11]
  PIN i_dout1_1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 416.200 4.000 416.800 ;
    END
  END i_dout1_1[12]
  PIN i_dout1_1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 432.520 4.000 433.120 ;
    END
  END i_dout1_1[13]
  PIN i_dout1_1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 496.440 823.900 497.040 ;
    END
  END i_dout1_1[14]
  PIN i_dout1_1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 798.650 0.000 798.930 4.000 ;
    END
  END i_dout1_1[15]
  PIN i_dout1_1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 800.030 0.000 800.310 4.000 ;
    END
  END i_dout1_1[16]
  PIN i_dout1_1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 533.160 823.900 533.760 ;
    END
  END i_dout1_1[17]
  PIN i_dout1_1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 691.930 830.620 692.210 834.620 ;
    END
  END i_dout1_1[18]
  PIN i_dout1_1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 582.800 823.900 583.400 ;
    END
  END i_dout1_1[19]
  PIN i_dout1_1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 55.120 823.900 55.720 ;
    END
  END i_dout1_1[1]
  PIN i_dout1_1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 589.600 4.000 590.200 ;
    END
  END i_dout1_1[20]
  PIN i_dout1_1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 619.520 823.900 620.120 ;
    END
  END i_dout1_1[21]
  PIN i_dout1_1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 668.480 823.900 669.080 ;
    END
  END i_dout1_1[22]
  PIN i_dout1_1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 742.530 830.620 742.810 834.620 ;
    END
  END i_dout1_1[23]
  PIN i_dout1_1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 692.960 823.900 693.560 ;
    END
  END i_dout1_1[24]
  PIN i_dout1_1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 652.840 4.000 653.440 ;
    END
  END i_dout1_1[25]
  PIN i_dout1_1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 813.830 0.000 814.110 4.000 ;
    END
  END i_dout1_1[26]
  PIN i_dout1_1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 770.590 830.620 770.870 834.620 ;
    END
  END i_dout1_1[27]
  PIN i_dout1_1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 819.810 0.000 820.090 4.000 ;
    END
  END i_dout1_1[28]
  PIN i_dout1_1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 784.390 830.620 784.670 834.620 ;
    END
  END i_dout1_1[29]
  PIN i_dout1_1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 101.360 4.000 101.960 ;
    END
  END i_dout1_1[2]
  PIN i_dout1_1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 793.590 830.620 793.870 834.620 ;
    END
  END i_dout1_1[30]
  PIN i_dout1_1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 816.590 830.620 816.870 834.620 ;
    END
  END i_dout1_1[31]
  PIN i_dout1_1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 140.800 823.900 141.400 ;
    END
  END i_dout1_1[3]
  PIN i_dout1_1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 164.600 4.000 165.200 ;
    END
  END i_dout1_1[4]
  PIN i_dout1_1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 195.880 4.000 196.480 ;
    END
  END i_dout1_1[5]
  PIN i_dout1_1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 300.600 823.900 301.200 ;
    END
  END i_dout1_1[6]
  PIN i_dout1_1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 613.270 830.620 613.550 834.620 ;
    END
  END i_dout1_1[7]
  PIN i_dout1_1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 290.400 4.000 291.000 ;
    END
  END i_dout1_1[8]
  PIN i_dout1_1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 338.000 4.000 338.600 ;
    END
  END i_dout1_1[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.390 830.620 2.670 834.620 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.850 830.620 141.130 834.620 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.110 830.620 155.390 834.620 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.910 830.620 169.190 834.620 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.710 830.620 182.990 834.620 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 830.620 196.790 834.620 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.310 830.620 210.590 834.620 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.110 830.620 224.390 834.620 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.370 830.620 238.650 834.620 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.170 830.620 252.450 834.620 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.970 830.620 266.250 834.620 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 830.620 16.470 834.620 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.770 830.620 280.050 834.620 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.570 830.620 293.850 834.620 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 307.830 830.620 308.110 834.620 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.630 830.620 321.910 834.620 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.430 830.620 335.710 834.620 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 349.230 830.620 349.510 834.620 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.030 830.620 363.310 834.620 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.290 830.620 377.570 834.620 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.090 830.620 391.370 834.620 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.890 830.620 405.170 834.620 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.990 830.620 30.270 834.620 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.690 830.620 418.970 834.620 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.490 830.620 432.770 834.620 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 446.290 830.620 446.570 834.620 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.550 830.620 460.830 834.620 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 474.350 830.620 474.630 834.620 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 488.150 830.620 488.430 834.620 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.950 830.620 502.230 834.620 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 515.750 830.620 516.030 834.620 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.790 830.620 44.070 834.620 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.590 830.620 57.870 834.620 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.390 830.620 71.670 834.620 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.650 830.620 85.930 834.620 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.450 830.620 99.730 834.620 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.250 830.620 113.530 834.620 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.050 830.620 127.330 834.620 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 830.620 7.270 834.620 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.450 830.620 145.730 834.620 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.710 830.620 159.990 834.620 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.510 830.620 173.790 834.620 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.310 830.620 187.590 834.620 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.110 830.620 201.390 834.620 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.910 830.620 215.190 834.620 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.170 830.620 229.450 834.620 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.970 830.620 243.250 834.620 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.770 830.620 257.050 834.620 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.570 830.620 270.850 834.620 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 830.620 21.070 834.620 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.370 830.620 284.650 834.620 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.170 830.620 298.450 834.620 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.430 830.620 312.710 834.620 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.230 830.620 326.510 834.620 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.030 830.620 340.310 834.620 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 353.830 830.620 354.110 834.620 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.630 830.620 367.910 834.620 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 381.890 830.620 382.170 834.620 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.690 830.620 395.970 834.620 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.490 830.620 409.770 834.620 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.590 830.620 34.870 834.620 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 423.290 830.620 423.570 834.620 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 437.090 830.620 437.370 834.620 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.890 830.620 451.170 834.620 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 465.150 830.620 465.430 834.620 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.950 830.620 479.230 834.620 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.750 830.620 493.030 834.620 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 506.550 830.620 506.830 834.620 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 520.350 830.620 520.630 834.620 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 830.620 48.670 834.620 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.190 830.620 62.470 834.620 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.990 830.620 76.270 834.620 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 830.620 90.530 834.620 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.050 830.620 104.330 834.620 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.850 830.620 118.130 834.620 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.650 830.620 131.930 834.620 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 830.620 11.870 834.620 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.050 830.620 150.330 834.620 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 830.620 164.590 834.620 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.110 830.620 178.390 834.620 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.910 830.620 192.190 834.620 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.710 830.620 205.990 834.620 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.510 830.620 219.790 834.620 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.770 830.620 234.050 834.620 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.570 830.620 247.850 834.620 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.370 830.620 261.650 834.620 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.170 830.620 275.450 834.620 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.390 830.620 25.670 834.620 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.970 830.620 289.250 834.620 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.230 830.620 303.510 834.620 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.030 830.620 317.310 834.620 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.830 830.620 331.110 834.620 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.630 830.620 344.910 834.620 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.430 830.620 358.710 834.620 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 372.230 830.620 372.510 834.620 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.490 830.620 386.770 834.620 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 400.290 830.620 400.570 834.620 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 414.090 830.620 414.370 834.620 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.190 830.620 39.470 834.620 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 427.890 830.620 428.170 834.620 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.690 830.620 441.970 834.620 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.950 830.620 456.230 834.620 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.750 830.620 470.030 834.620 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.550 830.620 483.830 834.620 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 497.350 830.620 497.630 834.620 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 511.150 830.620 511.430 834.620 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.950 830.620 525.230 834.620 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.990 830.620 53.270 834.620 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.790 830.620 67.070 834.620 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.050 830.620 81.330 834.620 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.850 830.620 95.130 834.620 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.650 830.620 108.930 834.620 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 830.620 122.730 834.620 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.250 830.620 136.530 834.620 ;
    END
  END io_out[9]
  PIN irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 734.250 0.000 734.530 4.000 ;
    END
  END irq[0]
  PIN irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 735.630 0.000 735.910 4.000 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.470 0.000 737.750 4.000 ;
    END
  END irq[2]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.250 0.000 159.530 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.670 0.000 608.950 4.000 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 612.810 0.000 613.090 4.000 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 617.410 0.000 617.690 4.000 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 622.010 0.000 622.290 4.000 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 626.610 0.000 626.890 4.000 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 630.750 0.000 631.030 4.000 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 635.350 0.000 635.630 4.000 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 639.950 0.000 640.230 4.000 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 644.550 0.000 644.830 4.000 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 649.150 0.000 649.430 4.000 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.870 0.000 204.150 4.000 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 653.290 0.000 653.570 4.000 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 657.890 0.000 658.170 4.000 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 662.490 0.000 662.770 4.000 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 667.090 0.000 667.370 4.000 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 671.230 0.000 671.510 4.000 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 675.830 0.000 676.110 4.000 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 680.430 0.000 680.710 4.000 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.030 0.000 685.310 4.000 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.170 0.000 689.450 4.000 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 693.770 0.000 694.050 4.000 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.470 0.000 208.750 4.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 698.370 0.000 698.650 4.000 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.970 0.000 703.250 4.000 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 707.570 0.000 707.850 4.000 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 711.710 0.000 711.990 4.000 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 716.310 0.000 716.590 4.000 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 720.910 0.000 721.190 4.000 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 725.510 0.000 725.790 4.000 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 729.650 0.000 729.930 4.000 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.070 0.000 213.350 4.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.670 0.000 217.950 4.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.810 0.000 222.090 4.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.410 0.000 226.690 4.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.010 0.000 231.290 4.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.610 0.000 235.890 4.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.210 0.000 240.490 4.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.350 0.000 244.630 4.000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.390 0.000 163.670 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.950 0.000 249.230 4.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.550 0.000 253.830 4.000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.150 0.000 258.430 4.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.290 0.000 262.570 4.000 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.890 0.000 267.170 4.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.490 0.000 271.770 4.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.090 0.000 276.370 4.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.230 0.000 280.510 4.000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.830 0.000 285.110 4.000 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.430 0.000 289.710 4.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.990 0.000 168.270 4.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.030 0.000 294.310 4.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.630 0.000 298.910 4.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.770 0.000 303.050 4.000 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 307.370 0.000 307.650 4.000 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.970 0.000 312.250 4.000 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.570 0.000 316.850 4.000 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 320.710 0.000 320.990 4.000 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.310 0.000 325.590 4.000 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.910 0.000 330.190 4.000 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.510 0.000 334.790 4.000 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.590 0.000 172.870 4.000 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.650 0.000 338.930 4.000 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.250 0.000 343.530 4.000 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.850 0.000 348.130 4.000 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.450 0.000 352.730 4.000 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.050 0.000 357.330 4.000 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.190 0.000 361.470 4.000 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.790 0.000 366.070 4.000 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.390 0.000 370.670 4.000 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.990 0.000 375.270 4.000 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.130 0.000 379.410 4.000 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 0.000 177.470 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.730 0.000 384.010 4.000 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 388.330 0.000 388.610 4.000 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.930 0.000 393.210 4.000 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.070 0.000 397.350 4.000 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 401.670 0.000 401.950 4.000 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 406.270 0.000 406.550 4.000 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.870 0.000 411.150 4.000 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.470 0.000 415.750 4.000 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 419.610 0.000 419.890 4.000 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 424.210 0.000 424.490 4.000 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.790 0.000 182.070 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.810 0.000 429.090 4.000 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 433.410 0.000 433.690 4.000 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 437.550 0.000 437.830 4.000 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 442.150 0.000 442.430 4.000 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 446.750 0.000 447.030 4.000 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 451.350 0.000 451.630 4.000 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.490 0.000 455.770 4.000 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.090 0.000 460.370 4.000 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 464.690 0.000 464.970 4.000 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.290 0.000 469.570 4.000 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.930 0.000 186.210 4.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.890 0.000 474.170 4.000 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.030 0.000 478.310 4.000 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 482.630 0.000 482.910 4.000 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 487.230 0.000 487.510 4.000 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 491.830 0.000 492.110 4.000 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.970 0.000 496.250 4.000 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 500.570 0.000 500.850 4.000 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.170 0.000 505.450 4.000 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 509.770 0.000 510.050 4.000 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 513.910 0.000 514.190 4.000 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.530 0.000 190.810 4.000 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.510 0.000 518.790 4.000 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 523.110 0.000 523.390 4.000 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 527.710 0.000 527.990 4.000 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 532.310 0.000 532.590 4.000 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 536.450 0.000 536.730 4.000 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.050 0.000 541.330 4.000 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 545.650 0.000 545.930 4.000 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 550.250 0.000 550.530 4.000 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 554.390 0.000 554.670 4.000 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 558.990 0.000 559.270 4.000 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.130 0.000 195.410 4.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 563.590 0.000 563.870 4.000 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 568.190 0.000 568.470 4.000 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 572.330 0.000 572.610 4.000 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.930 0.000 577.210 4.000 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.530 0.000 581.810 4.000 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.130 0.000 586.410 4.000 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 590.730 0.000 591.010 4.000 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 594.870 0.000 595.150 4.000 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.470 0.000 599.750 4.000 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 604.070 0.000 604.350 4.000 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.730 0.000 200.010 4.000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.630 0.000 160.910 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 610.050 0.000 610.330 4.000 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 614.650 0.000 614.930 4.000 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 618.790 0.000 619.070 4.000 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 623.390 0.000 623.670 4.000 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.990 0.000 628.270 4.000 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 632.590 0.000 632.870 4.000 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 636.730 0.000 637.010 4.000 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 641.330 0.000 641.610 4.000 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 645.930 0.000 646.210 4.000 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.530 0.000 650.810 4.000 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.710 0.000 205.990 4.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 655.130 0.000 655.410 4.000 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 659.270 0.000 659.550 4.000 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 663.870 0.000 664.150 4.000 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 668.470 0.000 668.750 4.000 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.070 0.000 673.350 4.000 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 677.210 0.000 677.490 4.000 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 681.810 0.000 682.090 4.000 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 686.410 0.000 686.690 4.000 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 691.010 0.000 691.290 4.000 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.150 0.000 695.430 4.000 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.850 0.000 210.130 4.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 699.750 0.000 700.030 4.000 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 704.350 0.000 704.630 4.000 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.950 0.000 709.230 4.000 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 713.550 0.000 713.830 4.000 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 717.690 0.000 717.970 4.000 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 722.290 0.000 722.570 4.000 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 726.890 0.000 727.170 4.000 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 731.490 0.000 731.770 4.000 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.450 0.000 214.730 4.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 0.000 219.330 4.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.650 0.000 223.930 4.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.790 0.000 228.070 4.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.390 0.000 232.670 4.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.990 0.000 237.270 4.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 0.000 241.870 4.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.190 0.000 246.470 4.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.230 0.000 165.510 4.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.330 0.000 250.610 4.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.930 0.000 255.210 4.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.530 0.000 259.810 4.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.130 0.000 264.410 4.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.270 0.000 268.550 4.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.870 0.000 273.150 4.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.470 0.000 277.750 4.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.070 0.000 282.350 4.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.210 0.000 286.490 4.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.810 0.000 291.090 4.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.370 0.000 169.650 4.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 295.410 0.000 295.690 4.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.010 0.000 300.290 4.000 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.610 0.000 304.890 4.000 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.750 0.000 309.030 4.000 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 313.350 0.000 313.630 4.000 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.950 0.000 318.230 4.000 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.550 0.000 322.830 4.000 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.690 0.000 326.970 4.000 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.290 0.000 331.570 4.000 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.890 0.000 336.170 4.000 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 0.000 174.250 4.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.490 0.000 340.770 4.000 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.630 0.000 344.910 4.000 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 349.230 0.000 349.510 4.000 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 353.830 0.000 354.110 4.000 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.430 0.000 358.710 4.000 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.030 0.000 363.310 4.000 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.170 0.000 367.450 4.000 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 371.770 0.000 372.050 4.000 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.370 0.000 376.650 4.000 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.970 0.000 381.250 4.000 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.570 0.000 178.850 4.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 385.110 0.000 385.390 4.000 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.710 0.000 389.990 4.000 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 394.310 0.000 394.590 4.000 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.910 0.000 399.190 4.000 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.050 0.000 403.330 4.000 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 407.650 0.000 407.930 4.000 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.250 0.000 412.530 4.000 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.850 0.000 417.130 4.000 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.450 0.000 421.730 4.000 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.590 0.000 425.870 4.000 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.170 0.000 183.450 4.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 430.190 0.000 430.470 4.000 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.790 0.000 435.070 4.000 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.390 0.000 439.670 4.000 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.530 0.000 443.810 4.000 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 448.130 0.000 448.410 4.000 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 452.730 0.000 453.010 4.000 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.330 0.000 457.610 4.000 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.470 0.000 461.750 4.000 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.070 0.000 466.350 4.000 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.670 0.000 470.950 4.000 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.770 0.000 188.050 4.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 475.270 0.000 475.550 4.000 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.870 0.000 480.150 4.000 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.010 0.000 484.290 4.000 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 488.610 0.000 488.890 4.000 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 493.210 0.000 493.490 4.000 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 497.810 0.000 498.090 4.000 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.950 0.000 502.230 4.000 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 506.550 0.000 506.830 4.000 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 511.150 0.000 511.430 4.000 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 515.750 0.000 516.030 4.000 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.910 0.000 192.190 4.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 519.890 0.000 520.170 4.000 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.490 0.000 524.770 4.000 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 529.090 0.000 529.370 4.000 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 533.690 0.000 533.970 4.000 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 538.290 0.000 538.570 4.000 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 542.430 0.000 542.710 4.000 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.030 0.000 547.310 4.000 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 551.630 0.000 551.910 4.000 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 556.230 0.000 556.510 4.000 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.370 0.000 560.650 4.000 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 0.000 196.790 4.000 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.970 0.000 565.250 4.000 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 569.570 0.000 569.850 4.000 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 574.170 0.000 574.450 4.000 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 578.310 0.000 578.590 4.000 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 582.910 0.000 583.190 4.000 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.510 0.000 587.790 4.000 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 592.110 0.000 592.390 4.000 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 596.710 0.000 596.990 4.000 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 600.850 0.000 601.130 4.000 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.450 0.000 605.730 4.000 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.110 0.000 201.390 4.000 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.010 0.000 162.290 4.000 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.430 0.000 611.710 4.000 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 616.030 0.000 616.310 4.000 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 620.630 0.000 620.910 4.000 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 624.770 0.000 625.050 4.000 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 629.370 0.000 629.650 4.000 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 633.970 0.000 634.250 4.000 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 638.570 0.000 638.850 4.000 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 642.710 0.000 642.990 4.000 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 647.310 0.000 647.590 4.000 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 651.910 0.000 652.190 4.000 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.090 0.000 207.370 4.000 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.510 0.000 656.790 4.000 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 661.110 0.000 661.390 4.000 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 665.250 0.000 665.530 4.000 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 669.850 0.000 670.130 4.000 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 674.450 0.000 674.730 4.000 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 679.050 0.000 679.330 4.000 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 683.190 0.000 683.470 4.000 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 687.790 0.000 688.070 4.000 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 692.390 0.000 692.670 4.000 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 696.990 0.000 697.270 4.000 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.690 0.000 211.970 4.000 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 701.130 0.000 701.410 4.000 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 705.730 0.000 706.010 4.000 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 710.330 0.000 710.610 4.000 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 714.930 0.000 715.210 4.000 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 719.530 0.000 719.810 4.000 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 723.670 0.000 723.950 4.000 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 728.270 0.000 728.550 4.000 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 732.870 0.000 733.150 4.000 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.830 0.000 216.110 4.000 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.430 0.000 220.710 4.000 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.030 0.000 225.310 4.000 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.630 0.000 229.910 4.000 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.770 0.000 234.050 4.000 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.370 0.000 238.650 4.000 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.970 0.000 243.250 4.000 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.570 0.000 247.850 4.000 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.610 0.000 166.890 4.000 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.170 0.000 252.450 4.000 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.310 0.000 256.590 4.000 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.910 0.000 261.190 4.000 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.510 0.000 265.790 4.000 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.110 0.000 270.390 4.000 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.250 0.000 274.530 4.000 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.850 0.000 279.130 4.000 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.450 0.000 283.730 4.000 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.050 0.000 288.330 4.000 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.190 0.000 292.470 4.000 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.210 0.000 171.490 4.000 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.790 0.000 297.070 4.000 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.390 0.000 301.670 4.000 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.990 0.000 306.270 4.000 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 310.590 0.000 310.870 4.000 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.730 0.000 315.010 4.000 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.330 0.000 319.610 4.000 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.930 0.000 324.210 4.000 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.530 0.000 328.810 4.000 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.670 0.000 332.950 4.000 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.270 0.000 337.550 4.000 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.350 0.000 175.630 4.000 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.870 0.000 342.150 4.000 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.470 0.000 346.750 4.000 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 350.610 0.000 350.890 4.000 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 355.210 0.000 355.490 4.000 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 359.810 0.000 360.090 4.000 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.410 0.000 364.690 4.000 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.010 0.000 369.290 4.000 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.150 0.000 373.430 4.000 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.750 0.000 378.030 4.000 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 382.350 0.000 382.630 4.000 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.950 0.000 180.230 4.000 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.950 0.000 387.230 4.000 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.090 0.000 391.370 4.000 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.690 0.000 395.970 4.000 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 400.290 0.000 400.570 4.000 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.890 0.000 405.170 4.000 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.030 0.000 409.310 4.000 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 413.630 0.000 413.910 4.000 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.230 0.000 418.510 4.000 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 422.830 0.000 423.110 4.000 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 427.430 0.000 427.710 4.000 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.550 0.000 184.830 4.000 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.570 0.000 431.850 4.000 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 436.170 0.000 436.450 4.000 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 440.770 0.000 441.050 4.000 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.370 0.000 445.650 4.000 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.510 0.000 449.790 4.000 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.110 0.000 454.390 4.000 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 458.710 0.000 458.990 4.000 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.310 0.000 463.590 4.000 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 467.450 0.000 467.730 4.000 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.050 0.000 472.330 4.000 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.150 0.000 189.430 4.000 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 476.650 0.000 476.930 4.000 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 481.250 0.000 481.530 4.000 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 485.850 0.000 486.130 4.000 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.990 0.000 490.270 4.000 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 494.590 0.000 494.870 4.000 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.190 0.000 499.470 4.000 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 503.790 0.000 504.070 4.000 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.930 0.000 508.210 4.000 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.530 0.000 512.810 4.000 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 517.130 0.000 517.410 4.000 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.750 0.000 194.030 4.000 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 521.730 0.000 522.010 4.000 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 525.870 0.000 526.150 4.000 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 530.470 0.000 530.750 4.000 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 535.070 0.000 535.350 4.000 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 539.670 0.000 539.950 4.000 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.270 0.000 544.550 4.000 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 548.410 0.000 548.690 4.000 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.010 0.000 553.290 4.000 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.610 0.000 557.890 4.000 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 562.210 0.000 562.490 4.000 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.890 0.000 198.170 4.000 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 566.350 0.000 566.630 4.000 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.950 0.000 571.230 4.000 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 575.550 0.000 575.830 4.000 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 580.150 0.000 580.430 4.000 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 584.290 0.000 584.570 4.000 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 588.890 0.000 589.170 4.000 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.490 0.000 593.770 4.000 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 598.090 0.000 598.370 4.000 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 602.690 0.000 602.970 4.000 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 606.830 0.000 607.110 4.000 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.490 0.000 202.770 4.000 ;
    END
  END la_oenb[9]
  PIN o_addr1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 539.210 830.620 539.490 834.620 ;
    END
  END o_addr1[0]
  PIN o_addr1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.610 830.620 557.890 834.620 ;
    END
  END o_addr1[1]
  PIN o_addr1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 752.190 0.000 752.470 4.000 ;
    END
  END o_addr1[2]
  PIN o_addr1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.960 4.000 149.560 ;
    END
  END o_addr1[3]
  PIN o_addr1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.240 4.000 180.840 ;
    END
  END o_addr1[4]
  PIN o_addr1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 767.370 0.000 767.650 4.000 ;
    END
  END o_addr1[5]
  PIN o_addr1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 770.130 0.000 770.410 4.000 ;
    END
  END o_addr1[6]
  PIN o_addr1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 274.760 4.000 275.360 ;
    END
  END o_addr1[7]
  PIN o_addr1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 783.930 0.000 784.210 4.000 ;
    END
  END o_addr1[8]
  PIN o_addr1_1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.160 4.000 23.760 ;
    END
  END o_addr1_1[0]
  PIN o_addr1_1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 79.600 823.900 80.200 ;
    END
  END o_addr1_1[1]
  PIN o_addr1_1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 750.810 0.000 751.090 4.000 ;
    END
  END o_addr1_1[2]
  PIN o_addr1_1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 153.040 823.900 153.640 ;
    END
  END o_addr1_1[3]
  PIN o_addr1_1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 762.770 0.000 763.050 4.000 ;
    END
  END o_addr1_1[4]
  PIN o_addr1_1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 211.520 4.000 212.120 ;
    END
  END o_addr1_1[5]
  PIN o_addr1_1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 604.070 830.620 604.350 834.620 ;
    END
  END o_addr1_1[6]
  PIN o_addr1_1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 777.950 0.000 778.230 4.000 ;
    END
  END o_addr1_1[7]
  PIN o_addr1_1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 782.090 0.000 782.370 4.000 ;
    END
  END o_addr1_1[8]
  PIN o_csb0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 6.160 823.900 6.760 ;
    END
  END o_csb0
  PIN o_csb0_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 738.850 0.000 739.130 4.000 ;
    END
  END o_csb0_1
  PIN o_csb1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 740.230 0.000 740.510 4.000 ;
    END
  END o_csb1
  PIN o_csb1_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 18.400 823.900 19.000 ;
    END
  END o_csb1_1
  PIN o_din0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.800 4.000 39.400 ;
    END
  END o_din0[0]
  PIN o_din0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 789.910 0.000 790.190 4.000 ;
    END
  END o_din0[10]
  PIN o_din0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 400.560 4.000 401.160 ;
    END
  END o_din0[11]
  PIN o_din0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 435.240 823.900 435.840 ;
    END
  END o_din0[12]
  PIN o_din0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 448.160 4.000 448.760 ;
    END
  END o_din0[13]
  PIN o_din0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 508.680 823.900 509.280 ;
    END
  END o_din0[14]
  PIN o_din0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 668.470 830.620 668.750 834.620 ;
    END
  END o_din0[15]
  PIN o_din0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 510.720 4.000 511.320 ;
    END
  END o_din0[16]
  PIN o_din0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 682.730 830.620 683.010 834.620 ;
    END
  END o_din0[17]
  PIN o_din0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 804.630 0.000 804.910 4.000 ;
    END
  END o_din0[18]
  PIN o_din0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 705.730 830.620 706.010 834.620 ;
    END
  END o_din0[19]
  PIN o_din0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 91.840 823.900 92.440 ;
    END
  END o_din0[1]
  PIN o_din0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 807.850 0.000 808.130 4.000 ;
    END
  END o_din0[20]
  PIN o_din0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 714.930 830.620 715.210 834.620 ;
    END
  END o_din0[21]
  PIN o_din0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 733.330 830.620 733.610 834.620 ;
    END
  END o_din0[22]
  PIN o_din0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 637.200 4.000 637.800 ;
    END
  END o_din0[23]
  PIN o_din0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 717.440 823.900 718.040 ;
    END
  END o_din0[24]
  PIN o_din0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 811.990 0.000 812.270 4.000 ;
    END
  END o_din0[25]
  PIN o_din0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 815.210 0.000 815.490 4.000 ;
    END
  END o_din0[26]
  PIN o_din0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 747.360 4.000 747.960 ;
    END
  END o_din0[27]
  PIN o_din0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 790.880 823.900 791.480 ;
    END
  END o_din0[28]
  PIN o_din0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 803.120 823.900 803.720 ;
    END
  END o_din0[29]
  PIN o_din0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 753.570 0.000 753.850 4.000 ;
    END
  END o_din0[2]
  PIN o_din0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 815.360 823.900 815.960 ;
    END
  END o_din0[30]
  PIN o_din0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 827.600 823.900 828.200 ;
    END
  END o_din0[31]
  PIN o_din0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 165.280 823.900 165.880 ;
    END
  END o_din0[3]
  PIN o_din0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 580.610 830.620 580.890 834.620 ;
    END
  END o_din0[4]
  PIN o_din0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 594.410 830.620 594.690 834.620 ;
    END
  END o_din0[5]
  PIN o_din0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 771.970 0.000 772.250 4.000 ;
    END
  END o_din0[6]
  PIN o_din0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 779.330 0.000 779.610 4.000 ;
    END
  END o_din0[7]
  PIN o_din0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 374.040 823.900 374.640 ;
    END
  END o_din0[8]
  PIN o_din0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 788.070 0.000 788.350 4.000 ;
    END
  END o_din0[9]
  PIN o_din0_1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END o_din0_1[0]
  PIN o_din0_1[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 636.270 830.620 636.550 834.620 ;
    END
  END o_din0_1[10]
  PIN o_din0_1[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 792.670 0.000 792.950 4.000 ;
    END
  END o_din0_1[11]
  PIN o_din0_1[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 795.890 0.000 796.170 4.000 ;
    END
  END o_din0_1[12]
  PIN o_din0_1[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 484.200 823.900 484.800 ;
    END
  END o_din0_1[13]
  PIN o_din0_1[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 659.270 830.620 659.550 834.620 ;
    END
  END o_din0_1[14]
  PIN o_din0_1[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 479.440 4.000 480.040 ;
    END
  END o_din0_1[15]
  PIN o_din0_1[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 803.250 0.000 803.530 4.000 ;
    END
  END o_din0_1[16]
  PIN o_din0_1[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 678.130 830.620 678.410 834.620 ;
    END
  END o_din0_1[17]
  PIN o_din0_1[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 701.130 830.620 701.410 834.620 ;
    END
  END o_din0_1[18]
  PIN o_din0_1[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 558.320 4.000 558.920 ;
    END
  END o_din0_1[19]
  PIN o_din0_1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 747.590 0.000 747.870 4.000 ;
    END
  END o_din0_1[1]
  PIN o_din0_1[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 806.010 0.000 806.290 4.000 ;
    END
  END o_din0_1[20]
  PIN o_din0_1[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 656.240 823.900 656.840 ;
    END
  END o_din0_1[21]
  PIN o_din0_1[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 728.730 830.620 729.010 834.620 ;
    END
  END o_din0_1[22]
  PIN o_din0_1[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 747.130 830.620 747.410 834.620 ;
    END
  END o_din0_1[23]
  PIN o_din0_1[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 705.200 823.900 705.800 ;
    END
  END o_din0_1[24]
  PIN o_din0_1[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 741.920 823.900 742.520 ;
    END
  END o_din0_1[25]
  PIN o_din0_1[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 715.400 4.000 716.000 ;
    END
  END o_din0_1[26]
  PIN o_din0_1[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 817.970 0.000 818.250 4.000 ;
    END
  END o_din0_1[27]
  PIN o_din0_1[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 779.790 830.620 780.070 834.620 ;
    END
  END o_din0_1[28]
  PIN o_din0_1[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 822.570 0.000 822.850 4.000 ;
    END
  END o_din0_1[29]
  PIN o_din0_1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 116.320 823.900 116.920 ;
    END
  END o_din0_1[2]
  PIN o_din0_1[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 807.390 830.620 807.670 834.620 ;
    END
  END o_din0_1[30]
  PIN o_din0_1[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 825.560 4.000 826.160 ;
    END
  END o_din0_1[31]
  PIN o_din0_1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 761.390 0.000 761.670 4.000 ;
    END
  END o_din0_1[3]
  PIN o_din0_1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 250.960 823.900 251.560 ;
    END
  END o_din0_1[4]
  PIN o_din0_1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 589.810 830.620 590.090 834.620 ;
    END
  END o_din0_1[5]
  PIN o_din0_1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.670 830.620 608.950 834.620 ;
    END
  END o_din0_1[6]
  PIN o_din0_1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 325.080 823.900 325.680 ;
    END
  END o_din0_1[7]
  PIN o_din0_1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 361.800 823.900 362.400 ;
    END
  END o_din0_1[8]
  PIN o_din0_1[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 622.470 830.620 622.750 834.620 ;
    END
  END o_din0_1[9]
  PIN o_waddr0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 543.810 830.620 544.090 834.620 ;
    END
  END o_waddr0[0]
  PIN o_waddr0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.080 4.000 70.680 ;
    END
  END o_waddr0[1]
  PIN o_waddr0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 755.410 0.000 755.690 4.000 ;
    END
  END o_waddr0[2]
  PIN o_waddr0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 189.760 823.900 190.360 ;
    END
  END o_waddr0[3]
  PIN o_waddr0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 764.150 0.000 764.430 4.000 ;
    END
  END o_waddr0[4]
  PIN o_waddr0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.840 4.000 228.440 ;
    END
  END o_waddr0[5]
  PIN o_waddr0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 312.840 823.900 313.440 ;
    END
  END o_waddr0[6]
  PIN o_waddr0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 349.560 823.900 350.160 ;
    END
  END o_waddr0[7]
  PIN o_waddr0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 785.310 0.000 785.590 4.000 ;
    END
  END o_waddr0[8]
  PIN o_waddr0_1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 744.830 0.000 745.110 4.000 ;
    END
  END o_waddr0_1[0]
  PIN o_waddr0_1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 562.210 830.620 562.490 834.620 ;
    END
  END o_waddr0_1[1]
  PIN o_waddr0_1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 128.560 823.900 129.160 ;
    END
  END o_waddr0_1[2]
  PIN o_waddr0_1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 177.520 823.900 178.120 ;
    END
  END o_waddr0_1[3]
  PIN o_waddr0_1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 585.210 830.620 585.490 834.620 ;
    END
  END o_waddr0_1[4]
  PIN o_waddr0_1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 288.360 823.900 288.960 ;
    END
  END o_waddr0_1[5]
  PIN o_waddr0_1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 773.350 0.000 773.630 4.000 ;
    END
  END o_waddr0_1[6]
  PIN o_waddr0_1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 337.320 823.900 337.920 ;
    END
  END o_waddr0_1[7]
  PIN o_waddr0_1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 386.280 823.900 386.880 ;
    END
  END o_waddr0_1[8]
  PIN o_web0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 530.010 830.620 530.290 834.620 ;
    END
  END o_web0
  PIN o_web0_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 30.640 823.900 31.240 ;
    END
  END o_web0_1
  PIN o_wmask0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 548.410 830.620 548.690 834.620 ;
    END
  END o_wmask0[0]
  PIN o_wmask0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 749.430 0.000 749.710 4.000 ;
    END
  END o_wmask0[1]
  PIN o_wmask0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 133.320 4.000 133.920 ;
    END
  END o_wmask0[2]
  PIN o_wmask0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.010 830.620 576.290 834.620 ;
    END
  END o_wmask0[3]
  PIN o_wmask0_1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 746.210 0.000 746.490 4.000 ;
    END
  END o_wmask0_1[0]
  PIN o_wmask0_1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.720 4.000 86.320 ;
    END
  END o_wmask0_1[1]
  PIN o_wmask0_1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 756.790 0.000 757.070 4.000 ;
    END
  END o_wmask0_1[2]
  PIN o_wmask0_1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 202.000 823.900 202.600 ;
    END
  END o_wmask0_1[3]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 821.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 821.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 821.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 821.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 821.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 821.680 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 821.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 821.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 821.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 821.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 821.680 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.550 0.000 0.830 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.930 0.000 2.210 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 0.000 3.590 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.290 0.000 9.570 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.350 0.000 60.630 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.950 0.000 65.230 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 0.000 69.370 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.690 0.000 73.970 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.290 0.000 78.570 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.890 0.000 83.170 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.630 0.000 91.910 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.230 0.000 96.510 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.830 0.000 101.110 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.270 0.000 15.550 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.970 0.000 105.250 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.170 0.000 114.450 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.770 0.000 119.050 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.370 0.000 123.650 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.510 0.000 127.790 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 0.000 132.390 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.710 0.000 136.990 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.310 0.000 141.590 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.450 0.000 145.730 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.250 0.000 21.530 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.050 0.000 150.330 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 0.000 154.930 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.230 0.000 27.510 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.210 0.000 33.490 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.810 0.000 38.090 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.410 0.000 42.690 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.550 0.000 46.830 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.150 0.000 51.430 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.750 0.000 56.030 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.690 0.000 4.970 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.670 0.000 10.950 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.730 0.000 62.010 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.330 0.000 66.610 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.070 0.000 75.350 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.670 0.000 79.950 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.270 0.000 84.550 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.870 0.000 89.150 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.010 0.000 93.290 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.610 0.000 97.890 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.210 0.000 102.490 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.650 0.000 16.930 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.810 0.000 107.090 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.950 0.000 111.230 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.550 0.000 115.830 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.150 0.000 120.430 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.750 0.000 125.030 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.350 0.000 129.630 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.490 0.000 133.770 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.090 0.000 138.370 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.690 0.000 142.970 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.290 0.000 147.570 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.430 0.000 151.710 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.030 0.000 156.310 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.610 0.000 28.890 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.590 0.000 34.870 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.190 0.000 39.470 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.790 0.000 44.070 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.530 0.000 52.810 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.130 0.000 57.410 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.510 0.000 12.790 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.110 0.000 63.390 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.310 0.000 72.590 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.910 0.000 77.190 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.050 0.000 81.330 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.650 0.000 85.930 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.850 0.000 95.130 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.990 0.000 99.270 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.590 0.000 103.870 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.490 0.000 18.770 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.190 0.000 108.470 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 0.000 113.070 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.930 0.000 117.210 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.530 0.000 121.810 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.130 0.000 126.410 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.730 0.000 131.010 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 0.000 135.610 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.470 0.000 139.750 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.070 0.000 144.350 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.670 0.000 148.950 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.470 0.000 24.750 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.270 0.000 153.550 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.410 0.000 157.690 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.450 0.000 30.730 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.430 0.000 36.710 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.570 0.000 40.850 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.770 0.000 50.050 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.370 0.000 54.650 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.510 0.000 58.790 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.890 0.000 14.170 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.870 0.000 20.150 4.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.830 0.000 32.110 4.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 0.000 6.810 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.910 0.000 8.190 4.000 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 8.245 823.715 827.815 ;
      LAYER met1 ;
        RECT 1.910 0.040 823.790 827.860 ;
      LAYER met2 ;
        RECT 0.550 830.340 2.110 830.620 ;
        RECT 2.950 830.340 6.710 830.620 ;
        RECT 7.550 830.340 11.310 830.620 ;
        RECT 12.150 830.340 15.910 830.620 ;
        RECT 16.750 830.340 20.510 830.620 ;
        RECT 21.350 830.340 25.110 830.620 ;
        RECT 25.950 830.340 29.710 830.620 ;
        RECT 30.550 830.340 34.310 830.620 ;
        RECT 35.150 830.340 38.910 830.620 ;
        RECT 39.750 830.340 43.510 830.620 ;
        RECT 44.350 830.340 48.110 830.620 ;
        RECT 48.950 830.340 52.710 830.620 ;
        RECT 53.550 830.340 57.310 830.620 ;
        RECT 58.150 830.340 61.910 830.620 ;
        RECT 62.750 830.340 66.510 830.620 ;
        RECT 67.350 830.340 71.110 830.620 ;
        RECT 71.950 830.340 75.710 830.620 ;
        RECT 76.550 830.340 80.770 830.620 ;
        RECT 81.610 830.340 85.370 830.620 ;
        RECT 86.210 830.340 89.970 830.620 ;
        RECT 90.810 830.340 94.570 830.620 ;
        RECT 95.410 830.340 99.170 830.620 ;
        RECT 100.010 830.340 103.770 830.620 ;
        RECT 104.610 830.340 108.370 830.620 ;
        RECT 109.210 830.340 112.970 830.620 ;
        RECT 113.810 830.340 117.570 830.620 ;
        RECT 118.410 830.340 122.170 830.620 ;
        RECT 123.010 830.340 126.770 830.620 ;
        RECT 127.610 830.340 131.370 830.620 ;
        RECT 132.210 830.340 135.970 830.620 ;
        RECT 136.810 830.340 140.570 830.620 ;
        RECT 141.410 830.340 145.170 830.620 ;
        RECT 146.010 830.340 149.770 830.620 ;
        RECT 150.610 830.340 154.830 830.620 ;
        RECT 155.670 830.340 159.430 830.620 ;
        RECT 160.270 830.340 164.030 830.620 ;
        RECT 164.870 830.340 168.630 830.620 ;
        RECT 169.470 830.340 173.230 830.620 ;
        RECT 174.070 830.340 177.830 830.620 ;
        RECT 178.670 830.340 182.430 830.620 ;
        RECT 183.270 830.340 187.030 830.620 ;
        RECT 187.870 830.340 191.630 830.620 ;
        RECT 192.470 830.340 196.230 830.620 ;
        RECT 197.070 830.340 200.830 830.620 ;
        RECT 201.670 830.340 205.430 830.620 ;
        RECT 206.270 830.340 210.030 830.620 ;
        RECT 210.870 830.340 214.630 830.620 ;
        RECT 215.470 830.340 219.230 830.620 ;
        RECT 220.070 830.340 223.830 830.620 ;
        RECT 224.670 830.340 228.890 830.620 ;
        RECT 229.730 830.340 233.490 830.620 ;
        RECT 234.330 830.340 238.090 830.620 ;
        RECT 238.930 830.340 242.690 830.620 ;
        RECT 243.530 830.340 247.290 830.620 ;
        RECT 248.130 830.340 251.890 830.620 ;
        RECT 252.730 830.340 256.490 830.620 ;
        RECT 257.330 830.340 261.090 830.620 ;
        RECT 261.930 830.340 265.690 830.620 ;
        RECT 266.530 830.340 270.290 830.620 ;
        RECT 271.130 830.340 274.890 830.620 ;
        RECT 275.730 830.340 279.490 830.620 ;
        RECT 280.330 830.340 284.090 830.620 ;
        RECT 284.930 830.340 288.690 830.620 ;
        RECT 289.530 830.340 293.290 830.620 ;
        RECT 294.130 830.340 297.890 830.620 ;
        RECT 298.730 830.340 302.950 830.620 ;
        RECT 303.790 830.340 307.550 830.620 ;
        RECT 308.390 830.340 312.150 830.620 ;
        RECT 312.990 830.340 316.750 830.620 ;
        RECT 317.590 830.340 321.350 830.620 ;
        RECT 322.190 830.340 325.950 830.620 ;
        RECT 326.790 830.340 330.550 830.620 ;
        RECT 331.390 830.340 335.150 830.620 ;
        RECT 335.990 830.340 339.750 830.620 ;
        RECT 340.590 830.340 344.350 830.620 ;
        RECT 345.190 830.340 348.950 830.620 ;
        RECT 349.790 830.340 353.550 830.620 ;
        RECT 354.390 830.340 358.150 830.620 ;
        RECT 358.990 830.340 362.750 830.620 ;
        RECT 363.590 830.340 367.350 830.620 ;
        RECT 368.190 830.340 371.950 830.620 ;
        RECT 372.790 830.340 377.010 830.620 ;
        RECT 377.850 830.340 381.610 830.620 ;
        RECT 382.450 830.340 386.210 830.620 ;
        RECT 387.050 830.340 390.810 830.620 ;
        RECT 391.650 830.340 395.410 830.620 ;
        RECT 396.250 830.340 400.010 830.620 ;
        RECT 400.850 830.340 404.610 830.620 ;
        RECT 405.450 830.340 409.210 830.620 ;
        RECT 410.050 830.340 413.810 830.620 ;
        RECT 414.650 830.340 418.410 830.620 ;
        RECT 419.250 830.340 423.010 830.620 ;
        RECT 423.850 830.340 427.610 830.620 ;
        RECT 428.450 830.340 432.210 830.620 ;
        RECT 433.050 830.340 436.810 830.620 ;
        RECT 437.650 830.340 441.410 830.620 ;
        RECT 442.250 830.340 446.010 830.620 ;
        RECT 446.850 830.340 450.610 830.620 ;
        RECT 451.450 830.340 455.670 830.620 ;
        RECT 456.510 830.340 460.270 830.620 ;
        RECT 461.110 830.340 464.870 830.620 ;
        RECT 465.710 830.340 469.470 830.620 ;
        RECT 470.310 830.340 474.070 830.620 ;
        RECT 474.910 830.340 478.670 830.620 ;
        RECT 479.510 830.340 483.270 830.620 ;
        RECT 484.110 830.340 487.870 830.620 ;
        RECT 488.710 830.340 492.470 830.620 ;
        RECT 493.310 830.340 497.070 830.620 ;
        RECT 497.910 830.340 501.670 830.620 ;
        RECT 502.510 830.340 506.270 830.620 ;
        RECT 507.110 830.340 510.870 830.620 ;
        RECT 511.710 830.340 515.470 830.620 ;
        RECT 516.310 830.340 520.070 830.620 ;
        RECT 520.910 830.340 524.670 830.620 ;
        RECT 525.510 830.340 529.730 830.620 ;
        RECT 530.570 830.340 534.330 830.620 ;
        RECT 535.170 830.340 538.930 830.620 ;
        RECT 539.770 830.340 543.530 830.620 ;
        RECT 544.370 830.340 548.130 830.620 ;
        RECT 548.970 830.340 552.730 830.620 ;
        RECT 553.570 830.340 557.330 830.620 ;
        RECT 558.170 830.340 561.930 830.620 ;
        RECT 562.770 830.340 566.530 830.620 ;
        RECT 567.370 830.340 571.130 830.620 ;
        RECT 571.970 830.340 575.730 830.620 ;
        RECT 576.570 830.340 580.330 830.620 ;
        RECT 581.170 830.340 584.930 830.620 ;
        RECT 585.770 830.340 589.530 830.620 ;
        RECT 590.370 830.340 594.130 830.620 ;
        RECT 594.970 830.340 598.730 830.620 ;
        RECT 599.570 830.340 603.790 830.620 ;
        RECT 604.630 830.340 608.390 830.620 ;
        RECT 609.230 830.340 612.990 830.620 ;
        RECT 613.830 830.340 617.590 830.620 ;
        RECT 618.430 830.340 622.190 830.620 ;
        RECT 623.030 830.340 626.790 830.620 ;
        RECT 627.630 830.340 631.390 830.620 ;
        RECT 632.230 830.340 635.990 830.620 ;
        RECT 636.830 830.340 640.590 830.620 ;
        RECT 641.430 830.340 645.190 830.620 ;
        RECT 646.030 830.340 649.790 830.620 ;
        RECT 650.630 830.340 654.390 830.620 ;
        RECT 655.230 830.340 658.990 830.620 ;
        RECT 659.830 830.340 663.590 830.620 ;
        RECT 664.430 830.340 668.190 830.620 ;
        RECT 669.030 830.340 672.790 830.620 ;
        RECT 673.630 830.340 677.850 830.620 ;
        RECT 678.690 830.340 682.450 830.620 ;
        RECT 683.290 830.340 687.050 830.620 ;
        RECT 687.890 830.340 691.650 830.620 ;
        RECT 692.490 830.340 696.250 830.620 ;
        RECT 697.090 830.340 700.850 830.620 ;
        RECT 701.690 830.340 705.450 830.620 ;
        RECT 706.290 830.340 710.050 830.620 ;
        RECT 710.890 830.340 714.650 830.620 ;
        RECT 715.490 830.340 719.250 830.620 ;
        RECT 720.090 830.340 723.850 830.620 ;
        RECT 724.690 830.340 728.450 830.620 ;
        RECT 729.290 830.340 733.050 830.620 ;
        RECT 733.890 830.340 737.650 830.620 ;
        RECT 738.490 830.340 742.250 830.620 ;
        RECT 743.090 830.340 746.850 830.620 ;
        RECT 747.690 830.340 751.910 830.620 ;
        RECT 752.750 830.340 756.510 830.620 ;
        RECT 757.350 830.340 761.110 830.620 ;
        RECT 761.950 830.340 765.710 830.620 ;
        RECT 766.550 830.340 770.310 830.620 ;
        RECT 771.150 830.340 774.910 830.620 ;
        RECT 775.750 830.340 779.510 830.620 ;
        RECT 780.350 830.340 784.110 830.620 ;
        RECT 784.950 830.340 788.710 830.620 ;
        RECT 789.550 830.340 793.310 830.620 ;
        RECT 794.150 830.340 797.910 830.620 ;
        RECT 798.750 830.340 802.510 830.620 ;
        RECT 803.350 830.340 807.110 830.620 ;
        RECT 807.950 830.340 811.710 830.620 ;
        RECT 812.550 830.340 816.310 830.620 ;
        RECT 817.150 830.340 820.910 830.620 ;
        RECT 821.750 830.340 823.770 830.620 ;
        RECT 0.550 4.280 823.770 830.340 ;
        RECT 1.110 0.010 1.650 4.280 ;
        RECT 2.490 0.010 3.030 4.280 ;
        RECT 3.870 0.010 4.410 4.280 ;
        RECT 5.250 0.010 6.250 4.280 ;
        RECT 7.090 0.010 7.630 4.280 ;
        RECT 8.470 0.010 9.010 4.280 ;
        RECT 9.850 0.010 10.390 4.280 ;
        RECT 11.230 0.010 12.230 4.280 ;
        RECT 13.070 0.010 13.610 4.280 ;
        RECT 14.450 0.010 14.990 4.280 ;
        RECT 15.830 0.010 16.370 4.280 ;
        RECT 17.210 0.010 18.210 4.280 ;
        RECT 19.050 0.010 19.590 4.280 ;
        RECT 20.430 0.010 20.970 4.280 ;
        RECT 21.810 0.010 22.350 4.280 ;
        RECT 23.190 0.010 24.190 4.280 ;
        RECT 25.030 0.010 25.570 4.280 ;
        RECT 26.410 0.010 26.950 4.280 ;
        RECT 27.790 0.010 28.330 4.280 ;
        RECT 29.170 0.010 30.170 4.280 ;
        RECT 31.010 0.010 31.550 4.280 ;
        RECT 32.390 0.010 32.930 4.280 ;
        RECT 33.770 0.010 34.310 4.280 ;
        RECT 35.150 0.010 36.150 4.280 ;
        RECT 36.990 0.010 37.530 4.280 ;
        RECT 38.370 0.010 38.910 4.280 ;
        RECT 39.750 0.010 40.290 4.280 ;
        RECT 41.130 0.010 42.130 4.280 ;
        RECT 42.970 0.010 43.510 4.280 ;
        RECT 44.350 0.010 44.890 4.280 ;
        RECT 45.730 0.010 46.270 4.280 ;
        RECT 47.110 0.010 48.110 4.280 ;
        RECT 48.950 0.010 49.490 4.280 ;
        RECT 50.330 0.010 50.870 4.280 ;
        RECT 51.710 0.010 52.250 4.280 ;
        RECT 53.090 0.010 54.090 4.280 ;
        RECT 54.930 0.010 55.470 4.280 ;
        RECT 56.310 0.010 56.850 4.280 ;
        RECT 57.690 0.010 58.230 4.280 ;
        RECT 59.070 0.010 60.070 4.280 ;
        RECT 60.910 0.010 61.450 4.280 ;
        RECT 62.290 0.010 62.830 4.280 ;
        RECT 63.670 0.010 64.670 4.280 ;
        RECT 65.510 0.010 66.050 4.280 ;
        RECT 66.890 0.010 67.430 4.280 ;
        RECT 68.270 0.010 68.810 4.280 ;
        RECT 69.650 0.010 70.650 4.280 ;
        RECT 71.490 0.010 72.030 4.280 ;
        RECT 72.870 0.010 73.410 4.280 ;
        RECT 74.250 0.010 74.790 4.280 ;
        RECT 75.630 0.010 76.630 4.280 ;
        RECT 77.470 0.010 78.010 4.280 ;
        RECT 78.850 0.010 79.390 4.280 ;
        RECT 80.230 0.010 80.770 4.280 ;
        RECT 81.610 0.010 82.610 4.280 ;
        RECT 83.450 0.010 83.990 4.280 ;
        RECT 84.830 0.010 85.370 4.280 ;
        RECT 86.210 0.010 86.750 4.280 ;
        RECT 87.590 0.010 88.590 4.280 ;
        RECT 89.430 0.010 89.970 4.280 ;
        RECT 90.810 0.010 91.350 4.280 ;
        RECT 92.190 0.010 92.730 4.280 ;
        RECT 93.570 0.010 94.570 4.280 ;
        RECT 95.410 0.010 95.950 4.280 ;
        RECT 96.790 0.010 97.330 4.280 ;
        RECT 98.170 0.010 98.710 4.280 ;
        RECT 99.550 0.010 100.550 4.280 ;
        RECT 101.390 0.010 101.930 4.280 ;
        RECT 102.770 0.010 103.310 4.280 ;
        RECT 104.150 0.010 104.690 4.280 ;
        RECT 105.530 0.010 106.530 4.280 ;
        RECT 107.370 0.010 107.910 4.280 ;
        RECT 108.750 0.010 109.290 4.280 ;
        RECT 110.130 0.010 110.670 4.280 ;
        RECT 111.510 0.010 112.510 4.280 ;
        RECT 113.350 0.010 113.890 4.280 ;
        RECT 114.730 0.010 115.270 4.280 ;
        RECT 116.110 0.010 116.650 4.280 ;
        RECT 117.490 0.010 118.490 4.280 ;
        RECT 119.330 0.010 119.870 4.280 ;
        RECT 120.710 0.010 121.250 4.280 ;
        RECT 122.090 0.010 123.090 4.280 ;
        RECT 123.930 0.010 124.470 4.280 ;
        RECT 125.310 0.010 125.850 4.280 ;
        RECT 126.690 0.010 127.230 4.280 ;
        RECT 128.070 0.010 129.070 4.280 ;
        RECT 129.910 0.010 130.450 4.280 ;
        RECT 131.290 0.010 131.830 4.280 ;
        RECT 132.670 0.010 133.210 4.280 ;
        RECT 134.050 0.010 135.050 4.280 ;
        RECT 135.890 0.010 136.430 4.280 ;
        RECT 137.270 0.010 137.810 4.280 ;
        RECT 138.650 0.010 139.190 4.280 ;
        RECT 140.030 0.010 141.030 4.280 ;
        RECT 141.870 0.010 142.410 4.280 ;
        RECT 143.250 0.010 143.790 4.280 ;
        RECT 144.630 0.010 145.170 4.280 ;
        RECT 146.010 0.010 147.010 4.280 ;
        RECT 147.850 0.010 148.390 4.280 ;
        RECT 149.230 0.010 149.770 4.280 ;
        RECT 150.610 0.010 151.150 4.280 ;
        RECT 151.990 0.010 152.990 4.280 ;
        RECT 153.830 0.010 154.370 4.280 ;
        RECT 155.210 0.010 155.750 4.280 ;
        RECT 156.590 0.010 157.130 4.280 ;
        RECT 157.970 0.010 158.970 4.280 ;
        RECT 159.810 0.010 160.350 4.280 ;
        RECT 161.190 0.010 161.730 4.280 ;
        RECT 162.570 0.010 163.110 4.280 ;
        RECT 163.950 0.010 164.950 4.280 ;
        RECT 165.790 0.010 166.330 4.280 ;
        RECT 167.170 0.010 167.710 4.280 ;
        RECT 168.550 0.010 169.090 4.280 ;
        RECT 169.930 0.010 170.930 4.280 ;
        RECT 171.770 0.010 172.310 4.280 ;
        RECT 173.150 0.010 173.690 4.280 ;
        RECT 174.530 0.010 175.070 4.280 ;
        RECT 175.910 0.010 176.910 4.280 ;
        RECT 177.750 0.010 178.290 4.280 ;
        RECT 179.130 0.010 179.670 4.280 ;
        RECT 180.510 0.010 181.510 4.280 ;
        RECT 182.350 0.010 182.890 4.280 ;
        RECT 183.730 0.010 184.270 4.280 ;
        RECT 185.110 0.010 185.650 4.280 ;
        RECT 186.490 0.010 187.490 4.280 ;
        RECT 188.330 0.010 188.870 4.280 ;
        RECT 189.710 0.010 190.250 4.280 ;
        RECT 191.090 0.010 191.630 4.280 ;
        RECT 192.470 0.010 193.470 4.280 ;
        RECT 194.310 0.010 194.850 4.280 ;
        RECT 195.690 0.010 196.230 4.280 ;
        RECT 197.070 0.010 197.610 4.280 ;
        RECT 198.450 0.010 199.450 4.280 ;
        RECT 200.290 0.010 200.830 4.280 ;
        RECT 201.670 0.010 202.210 4.280 ;
        RECT 203.050 0.010 203.590 4.280 ;
        RECT 204.430 0.010 205.430 4.280 ;
        RECT 206.270 0.010 206.810 4.280 ;
        RECT 207.650 0.010 208.190 4.280 ;
        RECT 209.030 0.010 209.570 4.280 ;
        RECT 210.410 0.010 211.410 4.280 ;
        RECT 212.250 0.010 212.790 4.280 ;
        RECT 213.630 0.010 214.170 4.280 ;
        RECT 215.010 0.010 215.550 4.280 ;
        RECT 216.390 0.010 217.390 4.280 ;
        RECT 218.230 0.010 218.770 4.280 ;
        RECT 219.610 0.010 220.150 4.280 ;
        RECT 220.990 0.010 221.530 4.280 ;
        RECT 222.370 0.010 223.370 4.280 ;
        RECT 224.210 0.010 224.750 4.280 ;
        RECT 225.590 0.010 226.130 4.280 ;
        RECT 226.970 0.010 227.510 4.280 ;
        RECT 228.350 0.010 229.350 4.280 ;
        RECT 230.190 0.010 230.730 4.280 ;
        RECT 231.570 0.010 232.110 4.280 ;
        RECT 232.950 0.010 233.490 4.280 ;
        RECT 234.330 0.010 235.330 4.280 ;
        RECT 236.170 0.010 236.710 4.280 ;
        RECT 237.550 0.010 238.090 4.280 ;
        RECT 238.930 0.010 239.930 4.280 ;
        RECT 240.770 0.010 241.310 4.280 ;
        RECT 242.150 0.010 242.690 4.280 ;
        RECT 243.530 0.010 244.070 4.280 ;
        RECT 244.910 0.010 245.910 4.280 ;
        RECT 246.750 0.010 247.290 4.280 ;
        RECT 248.130 0.010 248.670 4.280 ;
        RECT 249.510 0.010 250.050 4.280 ;
        RECT 250.890 0.010 251.890 4.280 ;
        RECT 252.730 0.010 253.270 4.280 ;
        RECT 254.110 0.010 254.650 4.280 ;
        RECT 255.490 0.010 256.030 4.280 ;
        RECT 256.870 0.010 257.870 4.280 ;
        RECT 258.710 0.010 259.250 4.280 ;
        RECT 260.090 0.010 260.630 4.280 ;
        RECT 261.470 0.010 262.010 4.280 ;
        RECT 262.850 0.010 263.850 4.280 ;
        RECT 264.690 0.010 265.230 4.280 ;
        RECT 266.070 0.010 266.610 4.280 ;
        RECT 267.450 0.010 267.990 4.280 ;
        RECT 268.830 0.010 269.830 4.280 ;
        RECT 270.670 0.010 271.210 4.280 ;
        RECT 272.050 0.010 272.590 4.280 ;
        RECT 273.430 0.010 273.970 4.280 ;
        RECT 274.810 0.010 275.810 4.280 ;
        RECT 276.650 0.010 277.190 4.280 ;
        RECT 278.030 0.010 278.570 4.280 ;
        RECT 279.410 0.010 279.950 4.280 ;
        RECT 280.790 0.010 281.790 4.280 ;
        RECT 282.630 0.010 283.170 4.280 ;
        RECT 284.010 0.010 284.550 4.280 ;
        RECT 285.390 0.010 285.930 4.280 ;
        RECT 286.770 0.010 287.770 4.280 ;
        RECT 288.610 0.010 289.150 4.280 ;
        RECT 289.990 0.010 290.530 4.280 ;
        RECT 291.370 0.010 291.910 4.280 ;
        RECT 292.750 0.010 293.750 4.280 ;
        RECT 294.590 0.010 295.130 4.280 ;
        RECT 295.970 0.010 296.510 4.280 ;
        RECT 297.350 0.010 298.350 4.280 ;
        RECT 299.190 0.010 299.730 4.280 ;
        RECT 300.570 0.010 301.110 4.280 ;
        RECT 301.950 0.010 302.490 4.280 ;
        RECT 303.330 0.010 304.330 4.280 ;
        RECT 305.170 0.010 305.710 4.280 ;
        RECT 306.550 0.010 307.090 4.280 ;
        RECT 307.930 0.010 308.470 4.280 ;
        RECT 309.310 0.010 310.310 4.280 ;
        RECT 311.150 0.010 311.690 4.280 ;
        RECT 312.530 0.010 313.070 4.280 ;
        RECT 313.910 0.010 314.450 4.280 ;
        RECT 315.290 0.010 316.290 4.280 ;
        RECT 317.130 0.010 317.670 4.280 ;
        RECT 318.510 0.010 319.050 4.280 ;
        RECT 319.890 0.010 320.430 4.280 ;
        RECT 321.270 0.010 322.270 4.280 ;
        RECT 323.110 0.010 323.650 4.280 ;
        RECT 324.490 0.010 325.030 4.280 ;
        RECT 325.870 0.010 326.410 4.280 ;
        RECT 327.250 0.010 328.250 4.280 ;
        RECT 329.090 0.010 329.630 4.280 ;
        RECT 330.470 0.010 331.010 4.280 ;
        RECT 331.850 0.010 332.390 4.280 ;
        RECT 333.230 0.010 334.230 4.280 ;
        RECT 335.070 0.010 335.610 4.280 ;
        RECT 336.450 0.010 336.990 4.280 ;
        RECT 337.830 0.010 338.370 4.280 ;
        RECT 339.210 0.010 340.210 4.280 ;
        RECT 341.050 0.010 341.590 4.280 ;
        RECT 342.430 0.010 342.970 4.280 ;
        RECT 343.810 0.010 344.350 4.280 ;
        RECT 345.190 0.010 346.190 4.280 ;
        RECT 347.030 0.010 347.570 4.280 ;
        RECT 348.410 0.010 348.950 4.280 ;
        RECT 349.790 0.010 350.330 4.280 ;
        RECT 351.170 0.010 352.170 4.280 ;
        RECT 353.010 0.010 353.550 4.280 ;
        RECT 354.390 0.010 354.930 4.280 ;
        RECT 355.770 0.010 356.770 4.280 ;
        RECT 357.610 0.010 358.150 4.280 ;
        RECT 358.990 0.010 359.530 4.280 ;
        RECT 360.370 0.010 360.910 4.280 ;
        RECT 361.750 0.010 362.750 4.280 ;
        RECT 363.590 0.010 364.130 4.280 ;
        RECT 364.970 0.010 365.510 4.280 ;
        RECT 366.350 0.010 366.890 4.280 ;
        RECT 367.730 0.010 368.730 4.280 ;
        RECT 369.570 0.010 370.110 4.280 ;
        RECT 370.950 0.010 371.490 4.280 ;
        RECT 372.330 0.010 372.870 4.280 ;
        RECT 373.710 0.010 374.710 4.280 ;
        RECT 375.550 0.010 376.090 4.280 ;
        RECT 376.930 0.010 377.470 4.280 ;
        RECT 378.310 0.010 378.850 4.280 ;
        RECT 379.690 0.010 380.690 4.280 ;
        RECT 381.530 0.010 382.070 4.280 ;
        RECT 382.910 0.010 383.450 4.280 ;
        RECT 384.290 0.010 384.830 4.280 ;
        RECT 385.670 0.010 386.670 4.280 ;
        RECT 387.510 0.010 388.050 4.280 ;
        RECT 388.890 0.010 389.430 4.280 ;
        RECT 390.270 0.010 390.810 4.280 ;
        RECT 391.650 0.010 392.650 4.280 ;
        RECT 393.490 0.010 394.030 4.280 ;
        RECT 394.870 0.010 395.410 4.280 ;
        RECT 396.250 0.010 396.790 4.280 ;
        RECT 397.630 0.010 398.630 4.280 ;
        RECT 399.470 0.010 400.010 4.280 ;
        RECT 400.850 0.010 401.390 4.280 ;
        RECT 402.230 0.010 402.770 4.280 ;
        RECT 403.610 0.010 404.610 4.280 ;
        RECT 405.450 0.010 405.990 4.280 ;
        RECT 406.830 0.010 407.370 4.280 ;
        RECT 408.210 0.010 408.750 4.280 ;
        RECT 409.590 0.010 410.590 4.280 ;
        RECT 411.430 0.010 411.970 4.280 ;
        RECT 412.810 0.010 413.350 4.280 ;
        RECT 414.190 0.010 415.190 4.280 ;
        RECT 416.030 0.010 416.570 4.280 ;
        RECT 417.410 0.010 417.950 4.280 ;
        RECT 418.790 0.010 419.330 4.280 ;
        RECT 420.170 0.010 421.170 4.280 ;
        RECT 422.010 0.010 422.550 4.280 ;
        RECT 423.390 0.010 423.930 4.280 ;
        RECT 424.770 0.010 425.310 4.280 ;
        RECT 426.150 0.010 427.150 4.280 ;
        RECT 427.990 0.010 428.530 4.280 ;
        RECT 429.370 0.010 429.910 4.280 ;
        RECT 430.750 0.010 431.290 4.280 ;
        RECT 432.130 0.010 433.130 4.280 ;
        RECT 433.970 0.010 434.510 4.280 ;
        RECT 435.350 0.010 435.890 4.280 ;
        RECT 436.730 0.010 437.270 4.280 ;
        RECT 438.110 0.010 439.110 4.280 ;
        RECT 439.950 0.010 440.490 4.280 ;
        RECT 441.330 0.010 441.870 4.280 ;
        RECT 442.710 0.010 443.250 4.280 ;
        RECT 444.090 0.010 445.090 4.280 ;
        RECT 445.930 0.010 446.470 4.280 ;
        RECT 447.310 0.010 447.850 4.280 ;
        RECT 448.690 0.010 449.230 4.280 ;
        RECT 450.070 0.010 451.070 4.280 ;
        RECT 451.910 0.010 452.450 4.280 ;
        RECT 453.290 0.010 453.830 4.280 ;
        RECT 454.670 0.010 455.210 4.280 ;
        RECT 456.050 0.010 457.050 4.280 ;
        RECT 457.890 0.010 458.430 4.280 ;
        RECT 459.270 0.010 459.810 4.280 ;
        RECT 460.650 0.010 461.190 4.280 ;
        RECT 462.030 0.010 463.030 4.280 ;
        RECT 463.870 0.010 464.410 4.280 ;
        RECT 465.250 0.010 465.790 4.280 ;
        RECT 466.630 0.010 467.170 4.280 ;
        RECT 468.010 0.010 469.010 4.280 ;
        RECT 469.850 0.010 470.390 4.280 ;
        RECT 471.230 0.010 471.770 4.280 ;
        RECT 472.610 0.010 473.610 4.280 ;
        RECT 474.450 0.010 474.990 4.280 ;
        RECT 475.830 0.010 476.370 4.280 ;
        RECT 477.210 0.010 477.750 4.280 ;
        RECT 478.590 0.010 479.590 4.280 ;
        RECT 480.430 0.010 480.970 4.280 ;
        RECT 481.810 0.010 482.350 4.280 ;
        RECT 483.190 0.010 483.730 4.280 ;
        RECT 484.570 0.010 485.570 4.280 ;
        RECT 486.410 0.010 486.950 4.280 ;
        RECT 487.790 0.010 488.330 4.280 ;
        RECT 489.170 0.010 489.710 4.280 ;
        RECT 490.550 0.010 491.550 4.280 ;
        RECT 492.390 0.010 492.930 4.280 ;
        RECT 493.770 0.010 494.310 4.280 ;
        RECT 495.150 0.010 495.690 4.280 ;
        RECT 496.530 0.010 497.530 4.280 ;
        RECT 498.370 0.010 498.910 4.280 ;
        RECT 499.750 0.010 500.290 4.280 ;
        RECT 501.130 0.010 501.670 4.280 ;
        RECT 502.510 0.010 503.510 4.280 ;
        RECT 504.350 0.010 504.890 4.280 ;
        RECT 505.730 0.010 506.270 4.280 ;
        RECT 507.110 0.010 507.650 4.280 ;
        RECT 508.490 0.010 509.490 4.280 ;
        RECT 510.330 0.010 510.870 4.280 ;
        RECT 511.710 0.010 512.250 4.280 ;
        RECT 513.090 0.010 513.630 4.280 ;
        RECT 514.470 0.010 515.470 4.280 ;
        RECT 516.310 0.010 516.850 4.280 ;
        RECT 517.690 0.010 518.230 4.280 ;
        RECT 519.070 0.010 519.610 4.280 ;
        RECT 520.450 0.010 521.450 4.280 ;
        RECT 522.290 0.010 522.830 4.280 ;
        RECT 523.670 0.010 524.210 4.280 ;
        RECT 525.050 0.010 525.590 4.280 ;
        RECT 526.430 0.010 527.430 4.280 ;
        RECT 528.270 0.010 528.810 4.280 ;
        RECT 529.650 0.010 530.190 4.280 ;
        RECT 531.030 0.010 532.030 4.280 ;
        RECT 532.870 0.010 533.410 4.280 ;
        RECT 534.250 0.010 534.790 4.280 ;
        RECT 535.630 0.010 536.170 4.280 ;
        RECT 537.010 0.010 538.010 4.280 ;
        RECT 538.850 0.010 539.390 4.280 ;
        RECT 540.230 0.010 540.770 4.280 ;
        RECT 541.610 0.010 542.150 4.280 ;
        RECT 542.990 0.010 543.990 4.280 ;
        RECT 544.830 0.010 545.370 4.280 ;
        RECT 546.210 0.010 546.750 4.280 ;
        RECT 547.590 0.010 548.130 4.280 ;
        RECT 548.970 0.010 549.970 4.280 ;
        RECT 550.810 0.010 551.350 4.280 ;
        RECT 552.190 0.010 552.730 4.280 ;
        RECT 553.570 0.010 554.110 4.280 ;
        RECT 554.950 0.010 555.950 4.280 ;
        RECT 556.790 0.010 557.330 4.280 ;
        RECT 558.170 0.010 558.710 4.280 ;
        RECT 559.550 0.010 560.090 4.280 ;
        RECT 560.930 0.010 561.930 4.280 ;
        RECT 562.770 0.010 563.310 4.280 ;
        RECT 564.150 0.010 564.690 4.280 ;
        RECT 565.530 0.010 566.070 4.280 ;
        RECT 566.910 0.010 567.910 4.280 ;
        RECT 568.750 0.010 569.290 4.280 ;
        RECT 570.130 0.010 570.670 4.280 ;
        RECT 571.510 0.010 572.050 4.280 ;
        RECT 572.890 0.010 573.890 4.280 ;
        RECT 574.730 0.010 575.270 4.280 ;
        RECT 576.110 0.010 576.650 4.280 ;
        RECT 577.490 0.010 578.030 4.280 ;
        RECT 578.870 0.010 579.870 4.280 ;
        RECT 580.710 0.010 581.250 4.280 ;
        RECT 582.090 0.010 582.630 4.280 ;
        RECT 583.470 0.010 584.010 4.280 ;
        RECT 584.850 0.010 585.850 4.280 ;
        RECT 586.690 0.010 587.230 4.280 ;
        RECT 588.070 0.010 588.610 4.280 ;
        RECT 589.450 0.010 590.450 4.280 ;
        RECT 591.290 0.010 591.830 4.280 ;
        RECT 592.670 0.010 593.210 4.280 ;
        RECT 594.050 0.010 594.590 4.280 ;
        RECT 595.430 0.010 596.430 4.280 ;
        RECT 597.270 0.010 597.810 4.280 ;
        RECT 598.650 0.010 599.190 4.280 ;
        RECT 600.030 0.010 600.570 4.280 ;
        RECT 601.410 0.010 602.410 4.280 ;
        RECT 603.250 0.010 603.790 4.280 ;
        RECT 604.630 0.010 605.170 4.280 ;
        RECT 606.010 0.010 606.550 4.280 ;
        RECT 607.390 0.010 608.390 4.280 ;
        RECT 609.230 0.010 609.770 4.280 ;
        RECT 610.610 0.010 611.150 4.280 ;
        RECT 611.990 0.010 612.530 4.280 ;
        RECT 613.370 0.010 614.370 4.280 ;
        RECT 615.210 0.010 615.750 4.280 ;
        RECT 616.590 0.010 617.130 4.280 ;
        RECT 617.970 0.010 618.510 4.280 ;
        RECT 619.350 0.010 620.350 4.280 ;
        RECT 621.190 0.010 621.730 4.280 ;
        RECT 622.570 0.010 623.110 4.280 ;
        RECT 623.950 0.010 624.490 4.280 ;
        RECT 625.330 0.010 626.330 4.280 ;
        RECT 627.170 0.010 627.710 4.280 ;
        RECT 628.550 0.010 629.090 4.280 ;
        RECT 629.930 0.010 630.470 4.280 ;
        RECT 631.310 0.010 632.310 4.280 ;
        RECT 633.150 0.010 633.690 4.280 ;
        RECT 634.530 0.010 635.070 4.280 ;
        RECT 635.910 0.010 636.450 4.280 ;
        RECT 637.290 0.010 638.290 4.280 ;
        RECT 639.130 0.010 639.670 4.280 ;
        RECT 640.510 0.010 641.050 4.280 ;
        RECT 641.890 0.010 642.430 4.280 ;
        RECT 643.270 0.010 644.270 4.280 ;
        RECT 645.110 0.010 645.650 4.280 ;
        RECT 646.490 0.010 647.030 4.280 ;
        RECT 647.870 0.010 648.870 4.280 ;
        RECT 649.710 0.010 650.250 4.280 ;
        RECT 651.090 0.010 651.630 4.280 ;
        RECT 652.470 0.010 653.010 4.280 ;
        RECT 653.850 0.010 654.850 4.280 ;
        RECT 655.690 0.010 656.230 4.280 ;
        RECT 657.070 0.010 657.610 4.280 ;
        RECT 658.450 0.010 658.990 4.280 ;
        RECT 659.830 0.010 660.830 4.280 ;
        RECT 661.670 0.010 662.210 4.280 ;
        RECT 663.050 0.010 663.590 4.280 ;
        RECT 664.430 0.010 664.970 4.280 ;
        RECT 665.810 0.010 666.810 4.280 ;
        RECT 667.650 0.010 668.190 4.280 ;
        RECT 669.030 0.010 669.570 4.280 ;
        RECT 670.410 0.010 670.950 4.280 ;
        RECT 671.790 0.010 672.790 4.280 ;
        RECT 673.630 0.010 674.170 4.280 ;
        RECT 675.010 0.010 675.550 4.280 ;
        RECT 676.390 0.010 676.930 4.280 ;
        RECT 677.770 0.010 678.770 4.280 ;
        RECT 679.610 0.010 680.150 4.280 ;
        RECT 680.990 0.010 681.530 4.280 ;
        RECT 682.370 0.010 682.910 4.280 ;
        RECT 683.750 0.010 684.750 4.280 ;
        RECT 685.590 0.010 686.130 4.280 ;
        RECT 686.970 0.010 687.510 4.280 ;
        RECT 688.350 0.010 688.890 4.280 ;
        RECT 689.730 0.010 690.730 4.280 ;
        RECT 691.570 0.010 692.110 4.280 ;
        RECT 692.950 0.010 693.490 4.280 ;
        RECT 694.330 0.010 694.870 4.280 ;
        RECT 695.710 0.010 696.710 4.280 ;
        RECT 697.550 0.010 698.090 4.280 ;
        RECT 698.930 0.010 699.470 4.280 ;
        RECT 700.310 0.010 700.850 4.280 ;
        RECT 701.690 0.010 702.690 4.280 ;
        RECT 703.530 0.010 704.070 4.280 ;
        RECT 704.910 0.010 705.450 4.280 ;
        RECT 706.290 0.010 707.290 4.280 ;
        RECT 708.130 0.010 708.670 4.280 ;
        RECT 709.510 0.010 710.050 4.280 ;
        RECT 710.890 0.010 711.430 4.280 ;
        RECT 712.270 0.010 713.270 4.280 ;
        RECT 714.110 0.010 714.650 4.280 ;
        RECT 715.490 0.010 716.030 4.280 ;
        RECT 716.870 0.010 717.410 4.280 ;
        RECT 718.250 0.010 719.250 4.280 ;
        RECT 720.090 0.010 720.630 4.280 ;
        RECT 721.470 0.010 722.010 4.280 ;
        RECT 722.850 0.010 723.390 4.280 ;
        RECT 724.230 0.010 725.230 4.280 ;
        RECT 726.070 0.010 726.610 4.280 ;
        RECT 727.450 0.010 727.990 4.280 ;
        RECT 728.830 0.010 729.370 4.280 ;
        RECT 730.210 0.010 731.210 4.280 ;
        RECT 732.050 0.010 732.590 4.280 ;
        RECT 733.430 0.010 733.970 4.280 ;
        RECT 734.810 0.010 735.350 4.280 ;
        RECT 736.190 0.010 737.190 4.280 ;
        RECT 738.030 0.010 738.570 4.280 ;
        RECT 739.410 0.010 739.950 4.280 ;
        RECT 740.790 0.010 741.330 4.280 ;
        RECT 742.170 0.010 743.170 4.280 ;
        RECT 744.010 0.010 744.550 4.280 ;
        RECT 745.390 0.010 745.930 4.280 ;
        RECT 746.770 0.010 747.310 4.280 ;
        RECT 748.150 0.010 749.150 4.280 ;
        RECT 749.990 0.010 750.530 4.280 ;
        RECT 751.370 0.010 751.910 4.280 ;
        RECT 752.750 0.010 753.290 4.280 ;
        RECT 754.130 0.010 755.130 4.280 ;
        RECT 755.970 0.010 756.510 4.280 ;
        RECT 757.350 0.010 757.890 4.280 ;
        RECT 758.730 0.010 759.270 4.280 ;
        RECT 760.110 0.010 761.110 4.280 ;
        RECT 761.950 0.010 762.490 4.280 ;
        RECT 763.330 0.010 763.870 4.280 ;
        RECT 764.710 0.010 765.710 4.280 ;
        RECT 766.550 0.010 767.090 4.280 ;
        RECT 767.930 0.010 768.470 4.280 ;
        RECT 769.310 0.010 769.850 4.280 ;
        RECT 770.690 0.010 771.690 4.280 ;
        RECT 772.530 0.010 773.070 4.280 ;
        RECT 773.910 0.010 774.450 4.280 ;
        RECT 775.290 0.010 775.830 4.280 ;
        RECT 776.670 0.010 777.670 4.280 ;
        RECT 778.510 0.010 779.050 4.280 ;
        RECT 779.890 0.010 780.430 4.280 ;
        RECT 781.270 0.010 781.810 4.280 ;
        RECT 782.650 0.010 783.650 4.280 ;
        RECT 784.490 0.010 785.030 4.280 ;
        RECT 785.870 0.010 786.410 4.280 ;
        RECT 787.250 0.010 787.790 4.280 ;
        RECT 788.630 0.010 789.630 4.280 ;
        RECT 790.470 0.010 791.010 4.280 ;
        RECT 791.850 0.010 792.390 4.280 ;
        RECT 793.230 0.010 793.770 4.280 ;
        RECT 794.610 0.010 795.610 4.280 ;
        RECT 796.450 0.010 796.990 4.280 ;
        RECT 797.830 0.010 798.370 4.280 ;
        RECT 799.210 0.010 799.750 4.280 ;
        RECT 800.590 0.010 801.590 4.280 ;
        RECT 802.430 0.010 802.970 4.280 ;
        RECT 803.810 0.010 804.350 4.280 ;
        RECT 805.190 0.010 805.730 4.280 ;
        RECT 806.570 0.010 807.570 4.280 ;
        RECT 808.410 0.010 808.950 4.280 ;
        RECT 809.790 0.010 810.330 4.280 ;
        RECT 811.170 0.010 811.710 4.280 ;
        RECT 812.550 0.010 813.550 4.280 ;
        RECT 814.390 0.010 814.930 4.280 ;
        RECT 815.770 0.010 816.310 4.280 ;
        RECT 817.150 0.010 817.690 4.280 ;
        RECT 818.530 0.010 819.530 4.280 ;
        RECT 820.370 0.010 820.910 4.280 ;
        RECT 821.750 0.010 822.290 4.280 ;
        RECT 823.130 0.010 823.770 4.280 ;
      LAYER met3 ;
        RECT 0.525 827.200 819.500 828.065 ;
        RECT 0.525 826.560 823.795 827.200 ;
        RECT 4.400 825.160 823.795 826.560 ;
        RECT 0.525 816.360 823.795 825.160 ;
        RECT 0.525 814.960 819.500 816.360 ;
        RECT 0.525 810.920 823.795 814.960 ;
        RECT 4.400 809.520 823.795 810.920 ;
        RECT 0.525 804.120 823.795 809.520 ;
        RECT 0.525 802.720 819.500 804.120 ;
        RECT 0.525 795.280 823.795 802.720 ;
        RECT 4.400 793.880 823.795 795.280 ;
        RECT 0.525 791.880 823.795 793.880 ;
        RECT 0.525 790.480 819.500 791.880 ;
        RECT 0.525 779.640 823.795 790.480 ;
        RECT 4.400 778.240 819.500 779.640 ;
        RECT 0.525 767.400 823.795 778.240 ;
        RECT 0.525 766.000 819.500 767.400 ;
        RECT 0.525 764.000 823.795 766.000 ;
        RECT 4.400 762.600 823.795 764.000 ;
        RECT 0.525 755.160 823.795 762.600 ;
        RECT 0.525 753.760 819.500 755.160 ;
        RECT 0.525 748.360 823.795 753.760 ;
        RECT 4.400 746.960 823.795 748.360 ;
        RECT 0.525 742.920 823.795 746.960 ;
        RECT 0.525 741.520 819.500 742.920 ;
        RECT 0.525 732.040 823.795 741.520 ;
        RECT 4.400 730.680 823.795 732.040 ;
        RECT 4.400 730.640 819.500 730.680 ;
        RECT 0.525 729.280 819.500 730.640 ;
        RECT 0.525 718.440 823.795 729.280 ;
        RECT 0.525 717.040 819.500 718.440 ;
        RECT 0.525 716.400 823.795 717.040 ;
        RECT 4.400 715.000 823.795 716.400 ;
        RECT 0.525 706.200 823.795 715.000 ;
        RECT 0.525 704.800 819.500 706.200 ;
        RECT 0.525 700.760 823.795 704.800 ;
        RECT 4.400 699.360 823.795 700.760 ;
        RECT 0.525 693.960 823.795 699.360 ;
        RECT 0.525 692.560 819.500 693.960 ;
        RECT 0.525 685.120 823.795 692.560 ;
        RECT 4.400 683.720 823.795 685.120 ;
        RECT 0.525 681.720 823.795 683.720 ;
        RECT 0.525 680.320 819.500 681.720 ;
        RECT 0.525 669.480 823.795 680.320 ;
        RECT 4.400 668.080 819.500 669.480 ;
        RECT 0.525 657.240 823.795 668.080 ;
        RECT 0.525 655.840 819.500 657.240 ;
        RECT 0.525 653.840 823.795 655.840 ;
        RECT 4.400 652.440 823.795 653.840 ;
        RECT 0.525 645.000 823.795 652.440 ;
        RECT 0.525 643.600 819.500 645.000 ;
        RECT 0.525 638.200 823.795 643.600 ;
        RECT 4.400 636.800 823.795 638.200 ;
        RECT 0.525 632.760 823.795 636.800 ;
        RECT 0.525 631.360 819.500 632.760 ;
        RECT 0.525 621.880 823.795 631.360 ;
        RECT 4.400 620.520 823.795 621.880 ;
        RECT 4.400 620.480 819.500 620.520 ;
        RECT 0.525 619.120 819.500 620.480 ;
        RECT 0.525 608.280 823.795 619.120 ;
        RECT 0.525 606.880 819.500 608.280 ;
        RECT 0.525 606.240 823.795 606.880 ;
        RECT 4.400 604.840 823.795 606.240 ;
        RECT 0.525 596.040 823.795 604.840 ;
        RECT 0.525 594.640 819.500 596.040 ;
        RECT 0.525 590.600 823.795 594.640 ;
        RECT 4.400 589.200 823.795 590.600 ;
        RECT 0.525 583.800 823.795 589.200 ;
        RECT 0.525 582.400 819.500 583.800 ;
        RECT 0.525 574.960 823.795 582.400 ;
        RECT 4.400 573.560 823.795 574.960 ;
        RECT 0.525 571.560 823.795 573.560 ;
        RECT 0.525 570.160 819.500 571.560 ;
        RECT 0.525 559.320 823.795 570.160 ;
        RECT 4.400 558.640 823.795 559.320 ;
        RECT 4.400 557.920 819.500 558.640 ;
        RECT 0.525 557.240 819.500 557.920 ;
        RECT 0.525 546.400 823.795 557.240 ;
        RECT 0.525 545.000 819.500 546.400 ;
        RECT 0.525 543.680 823.795 545.000 ;
        RECT 4.400 542.280 823.795 543.680 ;
        RECT 0.525 534.160 823.795 542.280 ;
        RECT 0.525 532.760 819.500 534.160 ;
        RECT 0.525 527.360 823.795 532.760 ;
        RECT 4.400 525.960 823.795 527.360 ;
        RECT 0.525 521.920 823.795 525.960 ;
        RECT 0.525 520.520 819.500 521.920 ;
        RECT 0.525 511.720 823.795 520.520 ;
        RECT 4.400 510.320 823.795 511.720 ;
        RECT 0.525 509.680 823.795 510.320 ;
        RECT 0.525 508.280 819.500 509.680 ;
        RECT 0.525 497.440 823.795 508.280 ;
        RECT 0.525 496.080 819.500 497.440 ;
        RECT 4.400 496.040 819.500 496.080 ;
        RECT 4.400 494.680 823.795 496.040 ;
        RECT 0.525 485.200 823.795 494.680 ;
        RECT 0.525 483.800 819.500 485.200 ;
        RECT 0.525 480.440 823.795 483.800 ;
        RECT 4.400 479.040 823.795 480.440 ;
        RECT 0.525 472.960 823.795 479.040 ;
        RECT 0.525 471.560 819.500 472.960 ;
        RECT 0.525 464.800 823.795 471.560 ;
        RECT 4.400 463.400 823.795 464.800 ;
        RECT 0.525 460.720 823.795 463.400 ;
        RECT 0.525 459.320 819.500 460.720 ;
        RECT 0.525 449.160 823.795 459.320 ;
        RECT 4.400 448.480 823.795 449.160 ;
        RECT 4.400 447.760 819.500 448.480 ;
        RECT 0.525 447.080 819.500 447.760 ;
        RECT 0.525 436.240 823.795 447.080 ;
        RECT 0.525 434.840 819.500 436.240 ;
        RECT 0.525 433.520 823.795 434.840 ;
        RECT 4.400 432.120 823.795 433.520 ;
        RECT 0.525 424.000 823.795 432.120 ;
        RECT 0.525 422.600 819.500 424.000 ;
        RECT 0.525 417.200 823.795 422.600 ;
        RECT 4.400 415.800 823.795 417.200 ;
        RECT 0.525 411.760 823.795 415.800 ;
        RECT 0.525 410.360 819.500 411.760 ;
        RECT 0.525 401.560 823.795 410.360 ;
        RECT 4.400 400.160 823.795 401.560 ;
        RECT 0.525 399.520 823.795 400.160 ;
        RECT 0.525 398.120 819.500 399.520 ;
        RECT 0.525 387.280 823.795 398.120 ;
        RECT 0.525 385.920 819.500 387.280 ;
        RECT 4.400 385.880 819.500 385.920 ;
        RECT 4.400 384.520 823.795 385.880 ;
        RECT 0.525 375.040 823.795 384.520 ;
        RECT 0.525 373.640 819.500 375.040 ;
        RECT 0.525 370.280 823.795 373.640 ;
        RECT 4.400 368.880 823.795 370.280 ;
        RECT 0.525 362.800 823.795 368.880 ;
        RECT 0.525 361.400 819.500 362.800 ;
        RECT 0.525 354.640 823.795 361.400 ;
        RECT 4.400 353.240 823.795 354.640 ;
        RECT 0.525 350.560 823.795 353.240 ;
        RECT 0.525 349.160 819.500 350.560 ;
        RECT 0.525 339.000 823.795 349.160 ;
        RECT 4.400 338.320 823.795 339.000 ;
        RECT 4.400 337.600 819.500 338.320 ;
        RECT 0.525 336.920 819.500 337.600 ;
        RECT 0.525 326.080 823.795 336.920 ;
        RECT 0.525 324.680 819.500 326.080 ;
        RECT 0.525 323.360 823.795 324.680 ;
        RECT 4.400 321.960 823.795 323.360 ;
        RECT 0.525 313.840 823.795 321.960 ;
        RECT 0.525 312.440 819.500 313.840 ;
        RECT 0.525 307.040 823.795 312.440 ;
        RECT 4.400 305.640 823.795 307.040 ;
        RECT 0.525 301.600 823.795 305.640 ;
        RECT 0.525 300.200 819.500 301.600 ;
        RECT 0.525 291.400 823.795 300.200 ;
        RECT 4.400 290.000 823.795 291.400 ;
        RECT 0.525 289.360 823.795 290.000 ;
        RECT 0.525 287.960 819.500 289.360 ;
        RECT 0.525 276.440 823.795 287.960 ;
        RECT 0.525 275.760 819.500 276.440 ;
        RECT 4.400 275.040 819.500 275.760 ;
        RECT 4.400 274.360 823.795 275.040 ;
        RECT 0.525 264.200 823.795 274.360 ;
        RECT 0.525 262.800 819.500 264.200 ;
        RECT 0.525 260.120 823.795 262.800 ;
        RECT 4.400 258.720 823.795 260.120 ;
        RECT 0.525 251.960 823.795 258.720 ;
        RECT 0.525 250.560 819.500 251.960 ;
        RECT 0.525 244.480 823.795 250.560 ;
        RECT 4.400 243.080 823.795 244.480 ;
        RECT 0.525 239.720 823.795 243.080 ;
        RECT 0.525 238.320 819.500 239.720 ;
        RECT 0.525 228.840 823.795 238.320 ;
        RECT 4.400 227.480 823.795 228.840 ;
        RECT 4.400 227.440 819.500 227.480 ;
        RECT 0.525 226.080 819.500 227.440 ;
        RECT 0.525 215.240 823.795 226.080 ;
        RECT 0.525 213.840 819.500 215.240 ;
        RECT 0.525 212.520 823.795 213.840 ;
        RECT 4.400 211.120 823.795 212.520 ;
        RECT 0.525 203.000 823.795 211.120 ;
        RECT 0.525 201.600 819.500 203.000 ;
        RECT 0.525 196.880 823.795 201.600 ;
        RECT 4.400 195.480 823.795 196.880 ;
        RECT 0.525 190.760 823.795 195.480 ;
        RECT 0.525 189.360 819.500 190.760 ;
        RECT 0.525 181.240 823.795 189.360 ;
        RECT 4.400 179.840 823.795 181.240 ;
        RECT 0.525 178.520 823.795 179.840 ;
        RECT 0.525 177.120 819.500 178.520 ;
        RECT 0.525 166.280 823.795 177.120 ;
        RECT 0.525 165.600 819.500 166.280 ;
        RECT 4.400 164.880 819.500 165.600 ;
        RECT 4.400 164.200 823.795 164.880 ;
        RECT 0.525 154.040 823.795 164.200 ;
        RECT 0.525 152.640 819.500 154.040 ;
        RECT 0.525 149.960 823.795 152.640 ;
        RECT 4.400 148.560 823.795 149.960 ;
        RECT 0.525 141.800 823.795 148.560 ;
        RECT 0.525 140.400 819.500 141.800 ;
        RECT 0.525 134.320 823.795 140.400 ;
        RECT 4.400 132.920 823.795 134.320 ;
        RECT 0.525 129.560 823.795 132.920 ;
        RECT 0.525 128.160 819.500 129.560 ;
        RECT 0.525 118.680 823.795 128.160 ;
        RECT 4.400 117.320 823.795 118.680 ;
        RECT 4.400 117.280 819.500 117.320 ;
        RECT 0.525 115.920 819.500 117.280 ;
        RECT 0.525 105.080 823.795 115.920 ;
        RECT 0.525 103.680 819.500 105.080 ;
        RECT 0.525 102.360 823.795 103.680 ;
        RECT 4.400 100.960 823.795 102.360 ;
        RECT 0.525 92.840 823.795 100.960 ;
        RECT 0.525 91.440 819.500 92.840 ;
        RECT 0.525 86.720 823.795 91.440 ;
        RECT 4.400 85.320 823.795 86.720 ;
        RECT 0.525 80.600 823.795 85.320 ;
        RECT 0.525 79.200 819.500 80.600 ;
        RECT 0.525 71.080 823.795 79.200 ;
        RECT 4.400 69.680 823.795 71.080 ;
        RECT 0.525 68.360 823.795 69.680 ;
        RECT 0.525 66.960 819.500 68.360 ;
        RECT 0.525 56.120 823.795 66.960 ;
        RECT 0.525 55.440 819.500 56.120 ;
        RECT 4.400 54.720 819.500 55.440 ;
        RECT 4.400 54.040 823.795 54.720 ;
        RECT 0.525 43.880 823.795 54.040 ;
        RECT 0.525 42.480 819.500 43.880 ;
        RECT 0.525 39.800 823.795 42.480 ;
        RECT 4.400 38.400 823.795 39.800 ;
        RECT 0.525 31.640 823.795 38.400 ;
        RECT 0.525 30.240 819.500 31.640 ;
        RECT 0.525 24.160 823.795 30.240 ;
        RECT 4.400 22.760 823.795 24.160 ;
        RECT 0.525 19.400 823.795 22.760 ;
        RECT 0.525 18.000 819.500 19.400 ;
        RECT 0.525 8.520 823.795 18.000 ;
        RECT 4.400 7.160 823.795 8.520 ;
        RECT 4.400 7.120 819.500 7.160 ;
        RECT 0.525 5.760 819.500 7.120 ;
        RECT 0.525 1.535 823.795 5.760 ;
      LAYER met4 ;
        RECT 5.815 10.240 20.640 781.825 ;
        RECT 23.040 10.240 97.440 781.825 ;
        RECT 99.840 10.240 174.240 781.825 ;
        RECT 176.640 10.240 251.040 781.825 ;
        RECT 253.440 10.240 327.840 781.825 ;
        RECT 330.240 10.240 404.640 781.825 ;
        RECT 407.040 10.240 481.440 781.825 ;
        RECT 483.840 10.240 558.240 781.825 ;
        RECT 560.640 10.240 635.040 781.825 ;
        RECT 637.440 10.240 711.840 781.825 ;
        RECT 714.240 10.240 788.640 781.825 ;
        RECT 791.040 10.240 817.585 781.825 ;
        RECT 5.815 2.895 817.585 10.240 ;
  END
END user_proj
END LIBRARY

