magic
tech sky130A
magscale 1 2
timestamp 1640373242
<< locali >>
rect 146309 504747 146343 504917
rect 155969 503727 156003 504577
rect 93719 503421 93869 503455
rect 196725 502367 196759 503421
rect 196725 483871 196759 487305
rect 219633 481423 219667 483361
rect 219725 480743 219759 486421
rect 219817 476117 219851 483225
rect 219817 476083 220771 476117
rect 219817 470543 219851 470645
rect 219817 451231 219851 451333
rect 219817 431919 219851 432021
rect 219725 422263 219759 422365
rect 220737 422297 220771 476083
rect 220001 422263 220771 422297
rect 219449 402883 219483 403053
rect 219541 402815 219575 412573
rect 219817 412539 219851 412709
rect 220001 412675 220035 422263
rect 187559 399993 187709 400027
rect 219483 398769 219575 398803
rect 219449 397919 219483 398565
rect 219541 398531 219575 398769
rect 219633 398735 219667 402917
rect 219541 397783 219575 398361
rect 108405 396695 108439 397069
rect 95893 396491 95927 396593
rect 221197 58395 221231 59177
rect 64521 57647 64555 57953
rect 66729 57307 66763 57681
rect 67005 57579 67039 57885
rect 70869 57783 70903 57953
rect 152381 57885 152691 57919
rect 152381 57851 152415 57885
rect 69121 57511 69155 57681
rect 66821 57307 66855 57477
rect 64889 56763 64923 57273
rect 64739 56729 64831 56763
rect 64245 56559 64279 56661
rect 64797 56627 64831 56729
rect 64981 56559 65015 56729
rect 66729 56559 66763 56865
rect 67925 56763 67959 57409
rect 68845 56899 68879 57205
rect 95433 57035 95467 57477
rect 102885 57443 102919 57749
rect 110521 57103 110555 57817
rect 111993 56899 112027 57341
rect 113097 56967 113131 57545
rect 68477 56559 68511 56797
rect 122665 56763 122699 57137
rect 122849 56627 122883 57681
rect 123309 56831 123343 57749
rect 135119 57613 135211 57647
rect 136407 57613 136741 57647
rect 138247 57613 138397 57647
rect 124781 56831 124815 57137
rect 124873 56899 124907 57137
rect 134901 57103 134935 57477
rect 124689 56763 124723 56797
rect 124965 56763 124999 56865
rect 124689 56729 124999 56763
rect 133889 56763 133923 57069
rect 135177 56831 135211 57613
rect 137201 57103 137235 57205
rect 137201 57069 137385 57103
rect 138121 56763 138155 57205
rect 140145 56763 140179 57341
rect 141341 56967 141375 57681
rect 143089 56899 143123 57545
rect 149345 57171 149379 57817
rect 152473 57647 152507 57817
rect 152657 57715 152691 57885
rect 152289 57613 152507 57647
rect 152289 57443 152323 57613
rect 152473 57307 152507 57545
rect 152415 57273 152507 57307
rect 152565 57239 152599 57681
rect 152657 57171 152691 57341
rect 152415 57137 152691 57171
rect 146401 56763 146435 57137
rect 138063 56729 138155 56763
rect 138213 56695 138247 56729
rect 138155 56661 138247 56695
rect 146309 56627 146343 56729
rect 156889 56559 156923 57681
rect 168297 57647 168331 57817
rect 171057 57783 171091 57817
rect 170815 57749 171091 57783
rect 157165 57035 157199 57613
rect 157073 56627 157107 57001
rect 157993 56627 158027 57545
rect 158821 56763 158855 57477
rect 159005 57171 159039 57409
rect 159097 57069 159373 57103
rect 159097 56967 159131 57069
rect 162133 57035 162167 57205
rect 162225 56899 162259 57613
rect 162133 56491 162167 56797
rect 166733 56559 166767 57409
rect 166917 56627 166951 56933
rect 170597 56695 170631 57205
rect 171149 56831 171183 57273
rect 177957 57137 178049 57171
rect 176577 56763 176611 57069
rect 177957 57035 177991 57137
rect 182465 56695 182499 57341
rect 183937 56899 183971 57069
rect 185535 57001 185685 57035
rect 200957 56831 200991 57477
rect 201785 56695 201819 57817
rect 223129 57103 223163 57613
rect 166917 56593 167101 56627
rect 205097 5015 205131 5117
rect 195253 4743 195287 4845
rect 205005 4675 205039 4981
rect 205189 4879 205223 5117
rect 59829 4063 59863 4097
rect 59829 4029 60013 4063
rect 64245 3995 64279 4097
rect 57989 2907 58023 3349
rect 58725 3247 58759 3417
rect 58909 3315 58943 3893
rect 60047 3893 60197 3927
rect 59001 3723 59035 3893
rect 59921 3451 59955 3825
rect 111717 3315 111751 4029
rect 476497 3315 476531 3621
<< viali >>
rect 146309 504917 146343 504951
rect 146309 504713 146343 504747
rect 155969 504577 156003 504611
rect 155969 503693 156003 503727
rect 93685 503421 93719 503455
rect 93869 503421 93903 503455
rect 196725 503421 196759 503455
rect 196725 502333 196759 502367
rect 196725 487305 196759 487339
rect 196725 483837 196759 483871
rect 219725 486421 219759 486455
rect 219633 483361 219667 483395
rect 219633 481389 219667 481423
rect 219725 480709 219759 480743
rect 219817 483225 219851 483259
rect 219817 470645 219851 470679
rect 219817 470509 219851 470543
rect 219817 451333 219851 451367
rect 219817 451197 219851 451231
rect 219817 432021 219851 432055
rect 219817 431885 219851 431919
rect 219725 422365 219759 422399
rect 219725 422229 219759 422263
rect 219817 412709 219851 412743
rect 219541 412573 219575 412607
rect 219449 403053 219483 403087
rect 219449 402849 219483 402883
rect 220001 412641 220035 412675
rect 219817 412505 219851 412539
rect 219541 402781 219575 402815
rect 219633 402917 219667 402951
rect 187525 399993 187559 400027
rect 187709 399993 187743 400027
rect 219449 398769 219483 398803
rect 219449 398565 219483 398599
rect 219633 398701 219667 398735
rect 219541 398497 219575 398531
rect 219449 397885 219483 397919
rect 219541 398361 219575 398395
rect 219541 397749 219575 397783
rect 108405 397069 108439 397103
rect 108405 396661 108439 396695
rect 95893 396593 95927 396627
rect 95893 396457 95927 396491
rect 221197 59177 221231 59211
rect 221197 58361 221231 58395
rect 64521 57953 64555 57987
rect 70869 57953 70903 57987
rect 67005 57885 67039 57919
rect 64521 57613 64555 57647
rect 66729 57681 66763 57715
rect 110521 57817 110555 57851
rect 70869 57749 70903 57783
rect 102885 57749 102919 57783
rect 67005 57545 67039 57579
rect 69121 57681 69155 57715
rect 64889 57273 64923 57307
rect 66729 57273 66763 57307
rect 66821 57477 66855 57511
rect 69121 57477 69155 57511
rect 95433 57477 95467 57511
rect 66821 57273 66855 57307
rect 67925 57409 67959 57443
rect 66729 56865 66763 56899
rect 64705 56729 64739 56763
rect 64889 56729 64923 56763
rect 64981 56729 65015 56763
rect 64245 56661 64279 56695
rect 64797 56593 64831 56627
rect 64245 56525 64279 56559
rect 64981 56525 65015 56559
rect 68845 57205 68879 57239
rect 102885 57409 102919 57443
rect 149345 57817 149379 57851
rect 152381 57817 152415 57851
rect 152473 57817 152507 57851
rect 123309 57749 123343 57783
rect 122849 57681 122883 57715
rect 113097 57545 113131 57579
rect 110521 57069 110555 57103
rect 111993 57341 112027 57375
rect 95433 57001 95467 57035
rect 68845 56865 68879 56899
rect 113097 56933 113131 56967
rect 122665 57137 122699 57171
rect 111993 56865 112027 56899
rect 67925 56729 67959 56763
rect 68477 56797 68511 56831
rect 66729 56525 66763 56559
rect 122665 56729 122699 56763
rect 141341 57681 141375 57715
rect 135085 57613 135119 57647
rect 136373 57613 136407 57647
rect 136741 57613 136775 57647
rect 138213 57613 138247 57647
rect 138397 57613 138431 57647
rect 134901 57477 134935 57511
rect 124781 57137 124815 57171
rect 124873 57137 124907 57171
rect 133889 57069 133923 57103
rect 134901 57069 134935 57103
rect 124873 56865 124907 56899
rect 124965 56865 124999 56899
rect 123309 56797 123343 56831
rect 124689 56797 124723 56831
rect 124781 56797 124815 56831
rect 140145 57341 140179 57375
rect 137201 57205 137235 57239
rect 138121 57205 138155 57239
rect 137385 57069 137419 57103
rect 135177 56797 135211 56831
rect 141341 56933 141375 56967
rect 143089 57545 143123 57579
rect 168297 57817 168331 57851
rect 152565 57681 152599 57715
rect 152657 57681 152691 57715
rect 156889 57681 156923 57715
rect 152289 57409 152323 57443
rect 152473 57545 152507 57579
rect 152381 57273 152415 57307
rect 152565 57205 152599 57239
rect 152657 57341 152691 57375
rect 143089 56865 143123 56899
rect 146401 57137 146435 57171
rect 149345 57137 149379 57171
rect 152381 57137 152415 57171
rect 133889 56729 133923 56763
rect 138029 56729 138063 56763
rect 138213 56729 138247 56763
rect 140145 56729 140179 56763
rect 146309 56729 146343 56763
rect 146401 56729 146435 56763
rect 138121 56661 138155 56695
rect 122849 56593 122883 56627
rect 146309 56593 146343 56627
rect 68477 56525 68511 56559
rect 171057 57817 171091 57851
rect 170781 57749 170815 57783
rect 201785 57817 201819 57851
rect 157165 57613 157199 57647
rect 162225 57613 162259 57647
rect 168297 57613 168331 57647
rect 157073 57001 157107 57035
rect 157165 57001 157199 57035
rect 157993 57545 158027 57579
rect 157073 56593 157107 56627
rect 158821 57477 158855 57511
rect 159005 57409 159039 57443
rect 159005 57137 159039 57171
rect 162133 57205 162167 57239
rect 159373 57069 159407 57103
rect 162133 57001 162167 57035
rect 159097 56933 159131 56967
rect 200957 57477 200991 57511
rect 162225 56865 162259 56899
rect 166733 57409 166767 57443
rect 158821 56729 158855 56763
rect 162133 56797 162167 56831
rect 157993 56593 158027 56627
rect 156889 56525 156923 56559
rect 182465 57341 182499 57375
rect 171149 57273 171183 57307
rect 170597 57205 170631 57239
rect 166917 56933 166951 56967
rect 178049 57137 178083 57171
rect 171149 56797 171183 56831
rect 176577 57069 176611 57103
rect 177957 57001 177991 57035
rect 176577 56729 176611 56763
rect 170597 56661 170631 56695
rect 183937 57069 183971 57103
rect 185501 57001 185535 57035
rect 185685 57001 185719 57035
rect 183937 56865 183971 56899
rect 200957 56797 200991 56831
rect 182465 56661 182499 56695
rect 223129 57613 223163 57647
rect 223129 57069 223163 57103
rect 201785 56661 201819 56695
rect 167101 56593 167135 56627
rect 166733 56525 166767 56559
rect 162133 56457 162167 56491
rect 205097 5117 205131 5151
rect 205005 4981 205039 5015
rect 205097 4981 205131 5015
rect 205189 5117 205223 5151
rect 195253 4845 195287 4879
rect 195253 4709 195287 4743
rect 205189 4845 205223 4879
rect 205005 4641 205039 4675
rect 59829 4097 59863 4131
rect 64245 4097 64279 4131
rect 60013 4029 60047 4063
rect 64245 3961 64279 3995
rect 111717 4029 111751 4063
rect 58909 3893 58943 3927
rect 58725 3417 58759 3451
rect 57989 3349 58023 3383
rect 59001 3893 59035 3927
rect 60013 3893 60047 3927
rect 60197 3893 60231 3927
rect 59001 3689 59035 3723
rect 59921 3825 59955 3859
rect 59921 3417 59955 3451
rect 58909 3281 58943 3315
rect 111717 3281 111751 3315
rect 476497 3621 476531 3655
rect 476497 3281 476531 3315
rect 58725 3213 58759 3247
rect 57989 2873 58023 2907
<< metal1 >>
rect 201494 702992 201500 703044
rect 201552 703032 201558 703044
rect 202782 703032 202788 703044
rect 201552 703004 202788 703032
rect 201552 702992 201558 703004
rect 202782 702992 202788 703004
rect 202840 702992 202846 703044
rect 204898 700680 204904 700732
rect 204956 700720 204962 700732
rect 235166 700720 235172 700732
rect 204956 700692 235172 700720
rect 204956 700680 204962 700692
rect 235166 700680 235172 700692
rect 235224 700680 235230 700732
rect 206370 700612 206376 700664
rect 206428 700652 206434 700664
rect 267642 700652 267648 700664
rect 206428 700624 267648 700652
rect 206428 700612 206434 700624
rect 267642 700612 267648 700624
rect 267700 700612 267706 700664
rect 213270 700544 213276 700596
rect 213328 700584 213334 700596
rect 283834 700584 283840 700596
rect 213328 700556 283840 700584
rect 213328 700544 213334 700556
rect 283834 700544 283840 700556
rect 283892 700544 283898 700596
rect 377398 700544 377404 700596
rect 377456 700584 377462 700596
rect 397454 700584 397460 700596
rect 377456 700556 397460 700584
rect 377456 700544 377462 700556
rect 397454 700544 397460 700556
rect 397512 700544 397518 700596
rect 446398 700544 446404 700596
rect 446456 700584 446462 700596
rect 494790 700584 494796 700596
rect 446456 700556 494796 700584
rect 446456 700544 446462 700556
rect 494790 700544 494796 700556
rect 494848 700544 494854 700596
rect 197998 700476 198004 700528
rect 198056 700516 198062 700528
rect 300118 700516 300124 700528
rect 198056 700488 300124 700516
rect 198056 700476 198062 700488
rect 300118 700476 300124 700488
rect 300176 700476 300182 700528
rect 376018 700476 376024 700528
rect 376076 700516 376082 700528
rect 462314 700516 462320 700528
rect 376076 700488 462320 700516
rect 376076 700476 376082 700488
rect 462314 700476 462320 700488
rect 462372 700476 462378 700528
rect 215938 700408 215944 700460
rect 215996 700448 216002 700460
rect 332502 700448 332508 700460
rect 215996 700420 332508 700448
rect 215996 700408 216002 700420
rect 332502 700408 332508 700420
rect 332560 700408 332566 700460
rect 388438 700408 388444 700460
rect 388496 700448 388502 700460
rect 478506 700448 478512 700460
rect 388496 700420 478512 700448
rect 388496 700408 388502 700420
rect 478506 700408 478512 700420
rect 478564 700408 478570 700460
rect 40494 700340 40500 700392
rect 40552 700380 40558 700392
rect 41322 700380 41328 700392
rect 40552 700352 41328 700380
rect 40552 700340 40558 700352
rect 41322 700340 41328 700352
rect 41380 700340 41386 700392
rect 170306 700340 170312 700392
rect 170364 700380 170370 700392
rect 196526 700380 196532 700392
rect 170364 700352 196532 700380
rect 170364 700340 170370 700352
rect 196526 700340 196532 700352
rect 196584 700340 196590 700392
rect 209038 700340 209044 700392
rect 209096 700380 209102 700392
rect 348786 700380 348792 700392
rect 209096 700352 348792 700380
rect 209096 700340 209102 700352
rect 348786 700340 348792 700352
rect 348844 700340 348850 700392
rect 374638 700340 374644 700392
rect 374696 700380 374702 700392
rect 527174 700380 527180 700392
rect 374696 700352 527180 700380
rect 374696 700340 374702 700352
rect 527174 700340 527180 700352
rect 527232 700340 527238 700392
rect 24302 700272 24308 700324
rect 24360 700312 24366 700324
rect 33778 700312 33784 700324
rect 24360 700284 33784 700312
rect 24360 700272 24366 700284
rect 33778 700272 33784 700284
rect 33836 700272 33842 700324
rect 59262 700272 59268 700324
rect 59320 700312 59326 700324
rect 72970 700312 72976 700324
rect 59320 700284 72976 700312
rect 59320 700272 59326 700284
rect 72970 700272 72976 700284
rect 73028 700272 73034 700324
rect 154114 700272 154120 700324
rect 154172 700312 154178 700324
rect 196618 700312 196624 700324
rect 154172 700284 196624 700312
rect 154172 700272 154178 700284
rect 196618 700272 196624 700284
rect 196676 700272 196682 700324
rect 214558 700272 214564 700324
rect 214616 700312 214622 700324
rect 559650 700312 559656 700324
rect 214616 700284 559656 700312
rect 214616 700272 214622 700284
rect 559650 700272 559656 700284
rect 559708 700272 559714 700324
rect 88334 699660 88340 699712
rect 88392 699700 88398 699712
rect 89162 699700 89168 699712
rect 88392 699672 89168 699700
rect 88392 699660 88398 699672
rect 89162 699660 89168 699672
rect 89220 699660 89226 699712
rect 104894 699660 104900 699712
rect 104952 699700 104958 699712
rect 105446 699700 105452 699712
rect 104952 699672 105452 699700
rect 104952 699660 104958 699672
rect 105446 699660 105452 699672
rect 105504 699660 105510 699712
rect 214650 699660 214656 699712
rect 214708 699700 214714 699712
rect 218974 699700 218980 699712
rect 214708 699672 218980 699700
rect 214708 699660 214714 699672
rect 218974 699660 218980 699672
rect 219032 699660 219038 699712
rect 360838 699660 360844 699712
rect 360896 699700 360902 699712
rect 364978 699700 364984 699712
rect 360896 699672 364984 699700
rect 360896 699660 360902 699672
rect 364978 699660 364984 699672
rect 365036 699660 365042 699712
rect 371878 696940 371884 696992
rect 371936 696980 371942 696992
rect 580166 696980 580172 696992
rect 371936 696952 580172 696980
rect 371936 696940 371942 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 138014 696872 138020 696924
rect 138072 696912 138078 696924
rect 140038 696912 140044 696924
rect 138072 696884 140044 696912
rect 138072 696872 138078 696884
rect 140038 696872 140044 696884
rect 140096 696872 140102 696924
rect 140038 689596 140044 689648
rect 140096 689636 140102 689648
rect 141142 689636 141148 689648
rect 140096 689608 141148 689636
rect 140096 689596 140102 689608
rect 141142 689596 141148 689608
rect 141200 689596 141206 689648
rect 141142 683612 141148 683664
rect 141200 683652 141206 683664
rect 143534 683652 143540 683664
rect 141200 683624 143540 683652
rect 141200 683612 141206 683624
rect 143534 683612 143540 683624
rect 143592 683612 143598 683664
rect 3418 683136 3424 683188
rect 3476 683176 3482 683188
rect 11698 683176 11704 683188
rect 3476 683148 11704 683176
rect 3476 683136 3482 683148
rect 11698 683136 11704 683148
rect 11756 683136 11762 683188
rect 385678 683136 385684 683188
rect 385736 683176 385742 683188
rect 580166 683176 580172 683188
rect 385736 683148 580172 683176
rect 385736 683136 385742 683148
rect 580166 683136 580172 683148
rect 580224 683136 580230 683188
rect 143534 680484 143540 680536
rect 143592 680524 143598 680536
rect 145558 680524 145564 680536
rect 143592 680496 145564 680524
rect 143592 680484 143598 680496
rect 145558 680484 145564 680496
rect 145616 680484 145622 680536
rect 3510 670692 3516 670744
rect 3568 670732 3574 670744
rect 36538 670732 36544 670744
rect 3568 670704 36544 670732
rect 3568 670692 3574 670704
rect 36538 670692 36544 670704
rect 36596 670692 36602 670744
rect 213362 670692 213368 670744
rect 213420 670732 213426 670744
rect 580166 670732 580172 670744
rect 213420 670704 580172 670732
rect 213420 670692 213426 670704
rect 580166 670692 580172 670704
rect 580224 670692 580230 670744
rect 145558 663212 145564 663264
rect 145616 663252 145622 663264
rect 149698 663252 149704 663264
rect 145616 663224 149704 663252
rect 145616 663212 145622 663224
rect 149698 663212 149704 663224
rect 149756 663212 149762 663264
rect 3418 656888 3424 656940
rect 3476 656928 3482 656940
rect 22738 656928 22744 656940
rect 3476 656900 22744 656928
rect 3476 656888 3482 656900
rect 22738 656888 22744 656900
rect 22796 656888 22802 656940
rect 149698 645872 149704 645924
rect 149756 645912 149762 645924
rect 149756 645884 151814 645912
rect 149756 645872 149762 645884
rect 151786 645844 151814 645884
rect 153194 645844 153200 645856
rect 151786 645816 153200 645844
rect 153194 645804 153200 645816
rect 153252 645804 153258 645856
rect 370498 643084 370504 643136
rect 370556 643124 370562 643136
rect 580166 643124 580172 643136
rect 370556 643096 580172 643124
rect 370556 643084 370562 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 153194 638868 153200 638920
rect 153252 638908 153258 638920
rect 155218 638908 155224 638920
rect 153252 638880 155224 638908
rect 153252 638868 153258 638880
rect 155218 638868 155224 638880
rect 155276 638868 155282 638920
rect 3418 632068 3424 632120
rect 3476 632108 3482 632120
rect 14458 632108 14464 632120
rect 3476 632080 14464 632108
rect 3476 632068 3482 632080
rect 14458 632068 14464 632080
rect 14516 632068 14522 632120
rect 382918 630640 382924 630692
rect 382976 630680 382982 630692
rect 580166 630680 580172 630692
rect 382976 630652 580172 630680
rect 382976 630640 382982 630652
rect 580166 630640 580172 630652
rect 580224 630640 580230 630692
rect 155218 627920 155224 627972
rect 155276 627960 155282 627972
rect 155276 627932 158760 627960
rect 155276 627920 155282 627932
rect 158732 627892 158760 627932
rect 160462 627892 160468 627904
rect 158732 627864 160468 627892
rect 160462 627852 160468 627864
rect 160520 627852 160526 627904
rect 160462 619624 160468 619676
rect 160520 619664 160526 619676
rect 160520 619636 161474 619664
rect 160520 619624 160526 619636
rect 161446 619596 161474 619636
rect 163498 619596 163504 619608
rect 161446 619568 163504 619596
rect 163498 619556 163504 619568
rect 163556 619556 163562 619608
rect 3142 618264 3148 618316
rect 3200 618304 3206 618316
rect 35158 618304 35164 618316
rect 3200 618276 35164 618304
rect 3200 618264 3206 618276
rect 35158 618264 35164 618276
rect 35216 618264 35222 618316
rect 209130 616836 209136 616888
rect 209188 616876 209194 616888
rect 580166 616876 580172 616888
rect 209188 616848 580172 616876
rect 209188 616836 209194 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 163498 611940 163504 611992
rect 163556 611980 163562 611992
rect 164878 611980 164884 611992
rect 163556 611952 164884 611980
rect 163556 611940 163562 611952
rect 164878 611940 164884 611952
rect 164936 611940 164942 611992
rect 3234 605820 3240 605872
rect 3292 605860 3298 605872
rect 25498 605860 25504 605872
rect 3292 605832 25504 605860
rect 3292 605820 3298 605832
rect 25498 605820 25504 605832
rect 25556 605820 25562 605872
rect 367738 590656 367744 590708
rect 367796 590696 367802 590708
rect 579798 590696 579804 590708
rect 367796 590668 579804 590696
rect 367796 590656 367802 590668
rect 579798 590656 579804 590668
rect 579856 590656 579862 590708
rect 164878 585692 164884 585744
rect 164936 585732 164942 585744
rect 167546 585732 167552 585744
rect 164936 585704 167552 585732
rect 164936 585692 164942 585704
rect 167546 585692 167552 585704
rect 167604 585692 167610 585744
rect 3326 579640 3332 579692
rect 3384 579680 3390 579692
rect 21358 579680 21364 579692
rect 3384 579652 21364 579680
rect 3384 579640 3390 579652
rect 21358 579640 21364 579652
rect 21416 579640 21422 579692
rect 167546 579572 167552 579624
rect 167604 579612 167610 579624
rect 170398 579612 170404 579624
rect 167604 579584 170404 579612
rect 167604 579572 167610 579584
rect 170398 579572 170404 579584
rect 170456 579572 170462 579624
rect 449158 576852 449164 576904
rect 449216 576892 449222 576904
rect 580166 576892 580172 576904
rect 449216 576864 580172 576892
rect 449216 576852 449222 576864
rect 580166 576852 580172 576864
rect 580224 576852 580230 576904
rect 170398 569100 170404 569152
rect 170456 569140 170462 569152
rect 172422 569140 172428 569152
rect 170456 569112 172428 569140
rect 170456 569100 170462 569112
rect 172422 569100 172428 569112
rect 172480 569100 172486 569152
rect 3418 565836 3424 565888
rect 3476 565876 3482 565888
rect 39298 565876 39304 565888
rect 3476 565848 39304 565876
rect 3476 565836 3482 565848
rect 39298 565836 39304 565848
rect 39356 565836 39362 565888
rect 172422 563048 172428 563100
rect 172480 563088 172486 563100
rect 172480 563060 172560 563088
rect 172480 563048 172486 563060
rect 172532 563020 172560 563060
rect 206278 563048 206284 563100
rect 206336 563088 206342 563100
rect 579798 563088 579804 563100
rect 206336 563060 579804 563088
rect 206336 563048 206342 563060
rect 579798 563048 579804 563060
rect 579856 563048 579862 563100
rect 178034 563020 178040 563032
rect 172532 562992 178040 563020
rect 178034 562980 178040 562992
rect 178092 562980 178098 563032
rect 178034 560192 178040 560244
rect 178092 560232 178098 560244
rect 180702 560232 180708 560244
rect 178092 560204 180708 560232
rect 178092 560192 178098 560204
rect 180702 560192 180708 560204
rect 180760 560192 180766 560244
rect 3418 553392 3424 553444
rect 3476 553432 3482 553444
rect 29638 553432 29644 553444
rect 3476 553404 29644 553432
rect 3476 553392 3482 553404
rect 29638 553392 29644 553404
rect 29696 553392 29702 553444
rect 180702 552032 180708 552084
rect 180760 552072 180766 552084
rect 180760 552032 180794 552072
rect 180766 552004 180794 552032
rect 182818 552004 182824 552016
rect 180766 551976 182824 552004
rect 182818 551964 182824 551976
rect 182876 551964 182882 552016
rect 182818 542308 182824 542360
rect 182876 542348 182882 542360
rect 184198 542348 184204 542360
rect 182876 542320 184204 542348
rect 182876 542308 182882 542320
rect 184198 542308 184204 542320
rect 184256 542308 184262 542360
rect 431218 536800 431224 536852
rect 431276 536840 431282 536852
rect 580166 536840 580172 536852
rect 431276 536812 580172 536840
rect 431276 536800 431282 536812
rect 580166 536800 580172 536812
rect 580224 536800 580230 536852
rect 184198 534080 184204 534132
rect 184256 534120 184262 534132
rect 186130 534120 186136 534132
rect 184256 534092 186136 534120
rect 184256 534080 184262 534092
rect 186130 534080 186136 534092
rect 186188 534080 186194 534132
rect 186130 531292 186136 531344
rect 186188 531332 186194 531344
rect 186188 531304 186360 531332
rect 186188 531292 186194 531304
rect 186332 531264 186360 531304
rect 187694 531264 187700 531276
rect 186332 531236 187700 531264
rect 187694 531224 187700 531236
rect 187752 531224 187758 531276
rect 187694 529184 187700 529236
rect 187752 529224 187758 529236
rect 196802 529224 196808 529236
rect 187752 529196 196808 529224
rect 187752 529184 187758 529196
rect 196802 529184 196808 529196
rect 196860 529184 196866 529236
rect 3418 527144 3424 527196
rect 3476 527184 3482 527196
rect 15838 527184 15844 527196
rect 3476 527156 15844 527184
rect 3476 527144 3482 527156
rect 15838 527144 15844 527156
rect 15896 527144 15902 527196
rect 381538 524424 381544 524476
rect 381596 524464 381602 524476
rect 580166 524464 580172 524476
rect 381596 524436 580172 524464
rect 381596 524424 381602 524436
rect 580166 524424 580172 524436
rect 580224 524424 580230 524476
rect 3418 514768 3424 514820
rect 3476 514808 3482 514820
rect 43438 514808 43444 514820
rect 3476 514780 43444 514808
rect 3476 514768 3482 514780
rect 43438 514768 43444 514780
rect 43496 514768 43502 514820
rect 204990 510620 204996 510672
rect 205048 510660 205054 510672
rect 580166 510660 580172 510672
rect 205048 510632 580172 510660
rect 205048 510620 205054 510632
rect 580166 510620 580172 510632
rect 580224 510620 580230 510672
rect 89622 505724 89628 505776
rect 89680 505764 89686 505776
rect 218882 505764 218888 505776
rect 89680 505736 218888 505764
rect 89680 505724 89686 505736
rect 218882 505724 218888 505736
rect 218940 505724 218946 505776
rect 114462 505656 114468 505708
rect 114520 505696 114526 505708
rect 218698 505696 218704 505708
rect 114520 505668 218704 505696
rect 114520 505656 114526 505668
rect 218698 505656 218704 505668
rect 218756 505656 218762 505708
rect 144822 505588 144828 505640
rect 144880 505628 144886 505640
rect 216306 505628 216312 505640
rect 144880 505600 216312 505628
rect 144880 505588 144886 505600
rect 216306 505588 216312 505600
rect 216364 505588 216370 505640
rect 142062 505520 142068 505572
rect 142120 505560 142126 505572
rect 216122 505560 216128 505572
rect 142120 505532 216128 505560
rect 142120 505520 142126 505532
rect 216122 505520 216128 505532
rect 216180 505520 216186 505572
rect 143350 505452 143356 505504
rect 143408 505492 143414 505504
rect 216490 505492 216496 505504
rect 143408 505464 216496 505492
rect 143408 505452 143414 505464
rect 216490 505452 216496 505464
rect 216548 505452 216554 505504
rect 219802 505452 219808 505504
rect 219860 505492 219866 505504
rect 260834 505492 260840 505504
rect 219860 505464 260840 505492
rect 219860 505452 219866 505464
rect 260834 505452 260840 505464
rect 260892 505452 260898 505504
rect 133782 505384 133788 505436
rect 133840 505424 133846 505436
rect 218790 505424 218796 505436
rect 133840 505396 218796 505424
rect 133840 505384 133846 505396
rect 218790 505384 218796 505396
rect 218848 505384 218854 505436
rect 219158 505384 219164 505436
rect 219216 505424 219222 505436
rect 288434 505424 288440 505436
rect 219216 505396 288440 505424
rect 219216 505384 219222 505396
rect 288434 505384 288440 505396
rect 288492 505384 288498 505436
rect 129642 505316 129648 505368
rect 129700 505356 129706 505368
rect 219250 505356 219256 505368
rect 129700 505328 219256 505356
rect 129700 505316 129706 505328
rect 219250 505316 219256 505328
rect 219308 505316 219314 505368
rect 219342 505316 219348 505368
rect 219400 505356 219406 505368
rect 298094 505356 298100 505368
rect 219400 505328 298100 505356
rect 219400 505316 219406 505328
rect 298094 505316 298100 505328
rect 298152 505316 298158 505368
rect 117222 505248 117228 505300
rect 117280 505288 117286 505300
rect 219066 505288 219072 505300
rect 117280 505260 219072 505288
rect 117280 505248 117286 505260
rect 219066 505248 219072 505260
rect 219124 505248 219130 505300
rect 219710 505248 219716 505300
rect 219768 505288 219774 505300
rect 300854 505288 300860 505300
rect 219768 505260 300860 505288
rect 219768 505248 219774 505260
rect 300854 505248 300860 505260
rect 300912 505248 300918 505300
rect 217778 505180 217784 505232
rect 217836 505220 217842 505232
rect 316034 505220 316040 505232
rect 217836 505192 316040 505220
rect 217836 505180 217842 505192
rect 316034 505180 316040 505192
rect 316092 505180 316098 505232
rect 218606 505112 218612 505164
rect 218664 505152 218670 505164
rect 325694 505152 325700 505164
rect 218664 505124 325700 505152
rect 218664 505112 218670 505124
rect 325694 505112 325700 505124
rect 325752 505112 325758 505164
rect 56502 505044 56508 505096
rect 56560 505084 56566 505096
rect 153194 505084 153200 505096
rect 56560 505056 153200 505084
rect 56560 505044 56566 505056
rect 153194 505044 153200 505056
rect 153252 505044 153258 505096
rect 158622 505044 158628 505096
rect 158680 505084 158686 505096
rect 219986 505084 219992 505096
rect 158680 505056 219992 505084
rect 158680 505044 158686 505056
rect 219986 505044 219992 505056
rect 220044 505044 220050 505096
rect 57606 504976 57612 505028
rect 57664 505016 57670 505028
rect 317414 505016 317420 505028
rect 57664 504988 317420 505016
rect 57664 504976 57670 504988
rect 317414 504976 317420 504988
rect 317472 504976 317478 505028
rect 53282 504908 53288 504960
rect 53340 504948 53346 504960
rect 128630 504948 128636 504960
rect 53340 504920 128636 504948
rect 53340 504908 53346 504920
rect 128630 504908 128636 504920
rect 128688 504908 128694 504960
rect 146297 504951 146355 504957
rect 142126 504920 146248 504948
rect 58342 504840 58348 504892
rect 58400 504880 58406 504892
rect 104894 504880 104900 504892
rect 58400 504852 104900 504880
rect 58400 504840 58406 504852
rect 104894 504840 104900 504852
rect 104952 504840 104958 504892
rect 108942 504840 108948 504892
rect 109000 504880 109006 504892
rect 142126 504880 142154 504920
rect 109000 504852 142154 504880
rect 146220 504880 146248 504920
rect 146297 504917 146309 504951
rect 146343 504948 146355 504951
rect 148502 504948 148508 504960
rect 146343 504920 148508 504948
rect 146343 504917 146355 504920
rect 146297 504911 146355 504917
rect 148502 504908 148508 504920
rect 148560 504908 148566 504960
rect 164050 504908 164056 504960
rect 164108 504948 164114 504960
rect 218974 504948 218980 504960
rect 164108 504920 218980 504948
rect 164108 504908 164114 504920
rect 218974 504908 218980 504920
rect 219032 504908 219038 504960
rect 219618 504908 219624 504960
rect 219676 504948 219682 504960
rect 273254 504948 273260 504960
rect 219676 504920 273260 504948
rect 219676 504908 219682 504920
rect 273254 504908 273260 504920
rect 273312 504908 273318 504960
rect 197446 504880 197452 504892
rect 146220 504852 197452 504880
rect 109000 504840 109006 504852
rect 197446 504840 197452 504852
rect 197504 504840 197510 504892
rect 219434 504840 219440 504892
rect 219492 504880 219498 504892
rect 277302 504880 277308 504892
rect 219492 504852 277308 504880
rect 219492 504840 219498 504852
rect 277302 504840 277308 504852
rect 277360 504840 277366 504892
rect 146570 504772 146576 504824
rect 146628 504812 146634 504824
rect 215754 504812 215760 504824
rect 146628 504784 215760 504812
rect 146628 504772 146634 504784
rect 215754 504772 215760 504784
rect 215812 504772 215818 504824
rect 218422 504772 218428 504824
rect 218480 504812 218486 504824
rect 277394 504812 277400 504824
rect 218480 504784 277400 504812
rect 218480 504772 218486 504784
rect 277394 504772 277400 504784
rect 277452 504772 277458 504824
rect 55030 504704 55036 504756
rect 55088 504744 55094 504756
rect 146297 504747 146355 504753
rect 146297 504744 146309 504747
rect 55088 504716 146309 504744
rect 55088 504704 55094 504716
rect 146297 504713 146309 504716
rect 146343 504713 146355 504747
rect 146297 504707 146355 504713
rect 149514 504704 149520 504756
rect 149572 504744 149578 504756
rect 215294 504744 215300 504756
rect 149572 504716 215300 504744
rect 149572 504704 149578 504716
rect 215294 504704 215300 504716
rect 215352 504704 215358 504756
rect 219526 504704 219532 504756
rect 219584 504744 219590 504756
rect 280154 504744 280160 504756
rect 219584 504716 280160 504744
rect 219584 504704 219590 504716
rect 280154 504704 280160 504716
rect 280212 504704 280218 504756
rect 98546 504636 98552 504688
rect 98604 504676 98610 504688
rect 197354 504676 197360 504688
rect 98604 504648 197360 504676
rect 98604 504636 98610 504648
rect 197354 504636 197360 504648
rect 197412 504636 197418 504688
rect 218330 504636 218336 504688
rect 218388 504676 218394 504688
rect 282914 504676 282920 504688
rect 218388 504648 282920 504676
rect 218388 504636 218394 504648
rect 282914 504636 282920 504648
rect 282972 504636 282978 504688
rect 57514 504568 57520 504620
rect 57572 504608 57578 504620
rect 155957 504611 156015 504617
rect 155957 504608 155969 504611
rect 57572 504580 155969 504608
rect 57572 504568 57578 504580
rect 155957 504577 155969 504580
rect 156003 504577 156015 504611
rect 155957 504571 156015 504577
rect 156046 504568 156052 504620
rect 156104 504608 156110 504620
rect 219894 504608 219900 504620
rect 156104 504580 219900 504608
rect 156104 504568 156110 504580
rect 219894 504568 219900 504580
rect 219952 504568 219958 504620
rect 111702 504500 111708 504552
rect 111760 504540 111766 504552
rect 215570 504540 215576 504552
rect 111760 504512 215576 504540
rect 111760 504500 111766 504512
rect 215570 504500 215576 504512
rect 215628 504500 215634 504552
rect 218514 504500 218520 504552
rect 218572 504540 218578 504552
rect 295334 504540 295340 504552
rect 218572 504512 295340 504540
rect 218572 504500 218578 504512
rect 295334 504500 295340 504512
rect 295392 504500 295398 504552
rect 56410 504432 56416 504484
rect 56468 504472 56474 504484
rect 165614 504472 165620 504484
rect 56468 504444 165620 504472
rect 56468 504432 56474 504444
rect 165614 504432 165620 504444
rect 165672 504432 165678 504484
rect 212442 504432 212448 504484
rect 212500 504472 212506 504484
rect 307754 504472 307760 504484
rect 212500 504444 307760 504472
rect 212500 504432 212506 504444
rect 307754 504432 307760 504444
rect 307812 504432 307818 504484
rect 59998 504364 60004 504416
rect 60056 504404 60062 504416
rect 88334 504404 88340 504416
rect 60056 504376 88340 504404
rect 60056 504364 60062 504376
rect 88334 504364 88340 504376
rect 88392 504364 88398 504416
rect 103882 504364 103888 504416
rect 103940 504404 103946 504416
rect 215478 504404 215484 504416
rect 103940 504376 215484 504404
rect 103940 504364 103946 504376
rect 215478 504364 215484 504376
rect 215536 504364 215542 504416
rect 216582 504364 216588 504416
rect 216640 504404 216646 504416
rect 313274 504404 313280 504416
rect 216640 504376 313280 504404
rect 216640 504364 216646 504376
rect 313274 504364 313280 504376
rect 313332 504364 313338 504416
rect 101306 504296 101312 504348
rect 101364 504336 101370 504348
rect 215846 504336 215852 504348
rect 101364 504308 215852 504336
rect 101364 504296 101370 504308
rect 215846 504296 215852 504308
rect 215904 504296 215910 504348
rect 216398 504296 216404 504348
rect 216456 504336 216462 504348
rect 320174 504336 320180 504348
rect 216456 504308 320180 504336
rect 216456 504296 216462 504308
rect 320174 504296 320180 504308
rect 320232 504296 320238 504348
rect 96522 504228 96528 504280
rect 96580 504268 96586 504280
rect 215662 504268 215668 504280
rect 96580 504240 215668 504268
rect 96580 504228 96586 504240
rect 215662 504228 215668 504240
rect 215720 504228 215726 504280
rect 216214 504228 216220 504280
rect 216272 504268 216278 504280
rect 322934 504268 322940 504280
rect 216272 504240 322940 504268
rect 216272 504228 216278 504240
rect 322934 504228 322940 504240
rect 322992 504228 322998 504280
rect 52270 504160 52276 504212
rect 52328 504200 52334 504212
rect 176838 504200 176844 504212
rect 52328 504172 176844 504200
rect 52328 504160 52334 504172
rect 176838 504160 176844 504172
rect 176896 504160 176902 504212
rect 206462 504160 206468 504212
rect 206520 504200 206526 504212
rect 339494 504200 339500 504212
rect 206520 504172 339500 504200
rect 206520 504160 206526 504172
rect 339494 504160 339500 504172
rect 339552 504160 339558 504212
rect 57790 504092 57796 504144
rect 57848 504132 57854 504144
rect 270494 504132 270500 504144
rect 57848 504104 270500 504132
rect 57848 504092 57854 504104
rect 270494 504092 270500 504104
rect 270552 504092 270558 504144
rect 50798 504024 50804 504076
rect 50856 504064 50862 504076
rect 265710 504064 265716 504076
rect 50856 504036 265716 504064
rect 50856 504024 50862 504036
rect 265710 504024 265716 504036
rect 265768 504024 265774 504076
rect 52178 503956 52184 504008
rect 52236 503996 52242 504008
rect 267734 503996 267740 504008
rect 52236 503968 267740 503996
rect 52236 503956 52242 503968
rect 267734 503956 267740 503968
rect 267792 503956 267798 504008
rect 50614 503888 50620 503940
rect 50672 503928 50678 503940
rect 302234 503928 302240 503940
rect 50672 503900 302240 503928
rect 50672 503888 50678 503900
rect 302234 503888 302240 503900
rect 302292 503888 302298 503940
rect 53190 503820 53196 503872
rect 53248 503860 53254 503872
rect 304994 503860 305000 503872
rect 53248 503832 305000 503860
rect 53248 503820 53254 503832
rect 304994 503820 305000 503832
rect 305052 503820 305058 503872
rect 55122 503752 55128 503804
rect 55180 503792 55186 503804
rect 310514 503792 310520 503804
rect 55180 503764 310520 503792
rect 55180 503752 55186 503764
rect 310514 503752 310520 503764
rect 310572 503752 310578 503804
rect 53374 503684 53380 503736
rect 53432 503724 53438 503736
rect 129734 503724 129740 503736
rect 53432 503696 129740 503724
rect 53432 503684 53438 503696
rect 129734 503684 129740 503696
rect 129792 503684 129798 503736
rect 155957 503727 156015 503733
rect 155957 503693 155969 503727
rect 156003 503724 156015 503727
rect 160094 503724 160100 503736
rect 156003 503696 160100 503724
rect 156003 503693 156015 503696
rect 155957 503687 156015 503693
rect 160094 503684 160100 503696
rect 160152 503684 160158 503736
rect 180702 503684 180708 503736
rect 180760 503724 180766 503736
rect 216030 503724 216036 503736
rect 180760 503696 216036 503724
rect 180760 503684 180766 503696
rect 216030 503684 216036 503696
rect 216088 503684 216094 503736
rect 218238 503684 218244 503736
rect 218296 503724 218302 503736
rect 292574 503724 292580 503736
rect 218296 503696 292580 503724
rect 218296 503684 218302 503696
rect 292574 503684 292580 503696
rect 292632 503684 292638 503736
rect 53466 503616 53472 503668
rect 53524 503656 53530 503668
rect 123754 503656 123760 503668
rect 53524 503628 123760 503656
rect 53524 503616 53530 503628
rect 123754 503616 123760 503628
rect 123812 503616 123818 503668
rect 220722 503616 220728 503668
rect 220780 503656 220786 503668
rect 245838 503656 245844 503668
rect 220780 503628 245844 503656
rect 220780 503616 220786 503628
rect 245838 503616 245844 503628
rect 245896 503616 245902 503668
rect 53650 503548 53656 503600
rect 53708 503588 53714 503600
rect 104066 503588 104072 503600
rect 53708 503560 104072 503588
rect 53708 503548 53714 503560
rect 104066 503548 104072 503560
rect 104124 503548 104130 503600
rect 201586 503588 201592 503600
rect 180766 503560 201592 503588
rect 93762 503480 93768 503532
rect 93820 503480 93826 503532
rect 123570 503480 123576 503532
rect 123628 503520 123634 503532
rect 180766 503520 180794 503560
rect 201586 503548 201592 503560
rect 201644 503548 201650 503600
rect 263594 503588 263600 503600
rect 209746 503560 263600 503588
rect 200206 503520 200212 503532
rect 123628 503492 180794 503520
rect 191668 503492 200212 503520
rect 123628 503480 123634 503492
rect 53558 503412 53564 503464
rect 53616 503452 53622 503464
rect 93673 503455 93731 503461
rect 93673 503452 93685 503455
rect 53616 503424 93685 503452
rect 53616 503412 53622 503424
rect 93673 503421 93685 503424
rect 93719 503421 93731 503455
rect 93673 503415 93731 503421
rect 93780 503384 93808 503480
rect 93857 503455 93915 503461
rect 93857 503421 93869 503455
rect 93903 503452 93915 503455
rect 113542 503452 113548 503464
rect 93903 503424 113548 503452
rect 93903 503421 93915 503424
rect 93857 503415 93915 503421
rect 113542 503412 113548 503424
rect 113600 503412 113606 503464
rect 121362 503412 121368 503464
rect 121420 503452 121426 503464
rect 191668 503452 191696 503492
rect 200206 503480 200212 503492
rect 200264 503480 200270 503532
rect 200758 503480 200764 503532
rect 200816 503520 200822 503532
rect 209746 503520 209774 503560
rect 263594 503548 263600 503560
rect 263652 503548 263658 503600
rect 200816 503492 209774 503520
rect 200816 503480 200822 503492
rect 218146 503480 218152 503532
rect 218204 503520 218210 503532
rect 285674 503520 285680 503532
rect 218204 503492 285680 503520
rect 218204 503480 218210 503492
rect 285674 503480 285680 503492
rect 285732 503480 285738 503532
rect 339402 503480 339408 503532
rect 339460 503520 339466 503532
rect 356514 503520 356520 503532
rect 339460 503492 356520 503520
rect 339460 503480 339466 503492
rect 356514 503480 356520 503492
rect 356572 503480 356578 503532
rect 121420 503424 191696 503452
rect 121420 503412 121426 503424
rect 191742 503412 191748 503464
rect 191800 503452 191806 503464
rect 196713 503455 196771 503461
rect 196713 503452 196725 503455
rect 191800 503424 196725 503452
rect 191800 503412 191806 503424
rect 196713 503421 196725 503424
rect 196759 503421 196771 503455
rect 196713 503415 196771 503421
rect 218054 503412 218060 503464
rect 218112 503452 218118 503464
rect 286870 503452 286876 503464
rect 218112 503424 286876 503452
rect 218112 503412 218118 503424
rect 286870 503412 286876 503424
rect 286928 503412 286934 503464
rect 350534 503412 350540 503464
rect 350592 503412 350598 503464
rect 93780 503356 196756 503384
rect 196728 503328 196756 503356
rect 213178 503344 213184 503396
rect 213236 503384 213242 503396
rect 350552 503384 350580 503412
rect 213236 503356 350580 503384
rect 213236 503344 213242 503356
rect 196710 503276 196716 503328
rect 196768 503276 196774 503328
rect 196713 502367 196771 502373
rect 196713 502333 196725 502367
rect 196759 502364 196771 502367
rect 213178 502364 213184 502376
rect 196759 502336 213184 502364
rect 196759 502333 196771 502336
rect 196713 502327 196771 502333
rect 213178 502324 213184 502336
rect 213236 502324 213242 502376
rect 2774 501032 2780 501084
rect 2832 501072 2838 501084
rect 4798 501072 4804 501084
rect 2832 501044 4804 501072
rect 2832 501032 2838 501044
rect 4798 501032 4804 501044
rect 4856 501032 4862 501084
rect 196710 487296 196716 487348
rect 196768 487336 196774 487348
rect 196768 487308 196813 487336
rect 196768 487296 196774 487308
rect 219713 486455 219771 486461
rect 219713 486421 219725 486455
rect 219759 486452 219771 486455
rect 219802 486452 219808 486464
rect 219759 486424 219808 486452
rect 219759 486421 219771 486424
rect 219713 486415 219771 486421
rect 219802 486412 219808 486424
rect 219860 486412 219866 486464
rect 196710 486344 196716 486396
rect 196768 486344 196774 486396
rect 196728 486192 196756 486344
rect 196710 486140 196716 486192
rect 196768 486140 196774 486192
rect 363598 484372 363604 484424
rect 363656 484412 363662 484424
rect 580166 484412 580172 484424
rect 363656 484384 580172 484412
rect 363656 484372 363662 484384
rect 580166 484372 580172 484384
rect 580224 484372 580230 484424
rect 196710 483828 196716 483880
rect 196768 483868 196774 483880
rect 196768 483840 196813 483868
rect 196768 483828 196774 483840
rect 219621 483395 219679 483401
rect 219621 483361 219633 483395
rect 219667 483392 219679 483395
rect 219802 483392 219808 483404
rect 219667 483364 219808 483392
rect 219667 483361 219679 483364
rect 219621 483355 219679 483361
rect 219802 483352 219808 483364
rect 219860 483352 219866 483404
rect 219802 483256 219808 483268
rect 219763 483228 219808 483256
rect 219802 483216 219808 483228
rect 219860 483216 219866 483268
rect 219621 481423 219679 481429
rect 219621 481389 219633 481423
rect 219667 481420 219679 481423
rect 219802 481420 219808 481432
rect 219667 481392 219808 481420
rect 219667 481389 219679 481392
rect 219621 481383 219679 481389
rect 219802 481380 219808 481392
rect 219860 481380 219866 481432
rect 219713 480743 219771 480749
rect 219713 480709 219725 480743
rect 219759 480740 219771 480743
rect 219802 480740 219808 480752
rect 219759 480712 219808 480740
rect 219759 480709 219771 480712
rect 219713 480703 219771 480709
rect 219802 480700 219808 480712
rect 219860 480700 219866 480752
rect 3418 474716 3424 474768
rect 3476 474756 3482 474768
rect 17218 474756 17224 474768
rect 3476 474728 17224 474756
rect 3476 474716 3482 474728
rect 17218 474716 17224 474728
rect 17276 474716 17282 474768
rect 219802 470676 219808 470688
rect 219763 470648 219808 470676
rect 219802 470636 219808 470648
rect 219860 470636 219866 470688
rect 443638 470568 443644 470620
rect 443696 470608 443702 470620
rect 579982 470608 579988 470620
rect 443696 470580 579988 470608
rect 443696 470568 443702 470580
rect 579982 470568 579988 470580
rect 580040 470568 580046 470620
rect 219802 470540 219808 470552
rect 219763 470512 219808 470540
rect 219802 470500 219808 470512
rect 219860 470500 219866 470552
rect 3234 462340 3240 462392
rect 3292 462380 3298 462392
rect 47578 462380 47584 462392
rect 3292 462352 47584 462380
rect 3292 462340 3298 462352
rect 47578 462340 47584 462352
rect 47636 462340 47642 462392
rect 358078 456764 358084 456816
rect 358136 456804 358142 456816
rect 580166 456804 580172 456816
rect 358136 456776 580172 456804
rect 358136 456764 358142 456776
rect 580166 456764 580172 456776
rect 580224 456764 580230 456816
rect 219802 451364 219808 451376
rect 219763 451336 219808 451364
rect 219802 451324 219808 451336
rect 219860 451324 219866 451376
rect 219802 451228 219808 451240
rect 219763 451200 219808 451228
rect 219802 451188 219808 451200
rect 219860 451188 219866 451240
rect 3142 448536 3148 448588
rect 3200 448576 3206 448588
rect 32398 448576 32404 448588
rect 3200 448548 32404 448576
rect 3200 448536 3206 448548
rect 32398 448536 32404 448548
rect 32456 448536 32462 448588
rect 219802 432052 219808 432064
rect 219763 432024 219808 432052
rect 219802 432012 219808 432024
rect 219860 432012 219866 432064
rect 219802 431916 219808 431928
rect 219763 431888 219808 431916
rect 219802 431876 219808 431888
rect 219860 431876 219866 431928
rect 210510 430584 210516 430636
rect 210568 430624 210574 430636
rect 216674 430624 216680 430636
rect 210568 430596 216680 430624
rect 210568 430584 210574 430596
rect 216674 430584 216680 430596
rect 216732 430584 216738 430636
rect 378778 430584 378784 430636
rect 378836 430624 378842 430636
rect 580166 430624 580172 430636
rect 378836 430596 580172 430624
rect 378836 430584 378842 430596
rect 580166 430584 580172 430596
rect 580224 430584 580230 430636
rect 50706 429156 50712 429208
rect 50764 429196 50770 429208
rect 57330 429196 57336 429208
rect 50764 429168 57336 429196
rect 50764 429156 50770 429168
rect 57330 429156 57336 429168
rect 57388 429156 57394 429208
rect 210602 429156 210608 429208
rect 210660 429196 210666 429208
rect 216674 429196 216680 429208
rect 210660 429168 216680 429196
rect 210660 429156 210666 429168
rect 216674 429156 216680 429168
rect 216732 429156 216738 429208
rect 57330 426640 57336 426692
rect 57388 426680 57394 426692
rect 57882 426680 57888 426692
rect 57388 426652 57888 426680
rect 57388 426640 57394 426652
rect 57882 426640 57888 426652
rect 57940 426640 57946 426692
rect 219713 422399 219771 422405
rect 219713 422365 219725 422399
rect 219759 422396 219771 422399
rect 219802 422396 219808 422408
rect 219759 422368 219808 422396
rect 219759 422365 219771 422368
rect 219713 422359 219771 422365
rect 219802 422356 219808 422368
rect 219860 422356 219866 422408
rect 3418 422288 3424 422340
rect 3476 422328 3482 422340
rect 18598 422328 18604 422340
rect 3476 422300 18604 422328
rect 3476 422288 3482 422300
rect 18598 422288 18604 422300
rect 18656 422288 18662 422340
rect 219713 422263 219771 422269
rect 219713 422229 219725 422263
rect 219759 422260 219771 422263
rect 219802 422260 219808 422272
rect 219759 422232 219808 422260
rect 219759 422229 219771 422232
rect 219713 422223 219771 422229
rect 219802 422220 219808 422232
rect 219860 422220 219866 422272
rect 219802 412740 219808 412752
rect 219763 412712 219808 412740
rect 219802 412700 219808 412712
rect 219860 412700 219866 412752
rect 219618 412632 219624 412684
rect 219676 412632 219682 412684
rect 219989 412675 220047 412681
rect 219989 412672 220001 412675
rect 219820 412646 220001 412672
rect 219529 412607 219587 412613
rect 219529 412573 219541 412607
rect 219575 412604 219587 412607
rect 219636 412604 219664 412632
rect 219575 412576 219664 412604
rect 219802 412594 219808 412646
rect 219860 412644 220001 412646
rect 219860 412594 219866 412644
rect 219989 412641 220001 412644
rect 220035 412641 220047 412675
rect 219989 412635 220047 412641
rect 219575 412573 219587 412576
rect 219529 412567 219587 412573
rect 219618 412496 219624 412548
rect 219676 412536 219682 412548
rect 219805 412539 219863 412545
rect 219805 412536 219817 412539
rect 219676 412508 219817 412536
rect 219676 412496 219682 412508
rect 219805 412505 219817 412508
rect 219851 412505 219863 412539
rect 219805 412499 219863 412505
rect 3142 409844 3148 409896
rect 3200 409884 3206 409896
rect 50338 409884 50344 409896
rect 3200 409856 50344 409884
rect 3200 409844 3206 409856
rect 50338 409844 50344 409856
rect 50396 409844 50402 409896
rect 210418 407872 210424 407924
rect 210476 407912 210482 407924
rect 213178 407912 213184 407924
rect 210476 407884 213184 407912
rect 210476 407872 210482 407884
rect 213178 407872 213184 407884
rect 213236 407912 213242 407924
rect 216674 407912 216680 407924
rect 213236 407884 216680 407912
rect 213236 407872 213242 407884
rect 216674 407872 216680 407884
rect 216732 407872 216738 407924
rect 210694 407124 210700 407176
rect 210752 407164 210758 407176
rect 216766 407164 216772 407176
rect 210752 407136 216772 407164
rect 210752 407124 210758 407136
rect 216766 407124 216772 407136
rect 216824 407124 216830 407176
rect 219618 405832 219624 405884
rect 219676 405832 219682 405884
rect 219636 405668 219664 405832
rect 219710 405668 219716 405680
rect 219636 405640 219716 405668
rect 219710 405628 219716 405640
rect 219768 405628 219774 405680
rect 425698 404336 425704 404388
rect 425756 404376 425762 404388
rect 580166 404376 580172 404388
rect 425756 404348 580172 404376
rect 425756 404336 425762 404348
rect 580166 404336 580172 404348
rect 580224 404336 580230 404388
rect 219434 403044 219440 403096
rect 219492 403084 219498 403096
rect 219492 403056 219537 403084
rect 219492 403044 219498 403056
rect 219526 402908 219532 402960
rect 219584 402948 219590 402960
rect 219621 402951 219679 402957
rect 219621 402948 219633 402951
rect 219584 402920 219633 402948
rect 219584 402908 219590 402920
rect 219621 402917 219633 402920
rect 219667 402917 219679 402951
rect 219621 402911 219679 402917
rect 219434 402840 219440 402892
rect 219492 402880 219498 402892
rect 219492 402852 219537 402880
rect 219492 402840 219498 402852
rect 219526 402812 219532 402824
rect 219487 402784 219532 402812
rect 219526 402772 219532 402784
rect 219584 402772 219590 402824
rect 197538 400092 197544 400104
rect 187620 400064 197544 400092
rect 187620 400036 187648 400064
rect 197538 400052 197544 400064
rect 197596 400052 197602 400104
rect 176562 399984 176568 400036
rect 176620 400024 176626 400036
rect 187513 400027 187571 400033
rect 187513 400024 187525 400027
rect 176620 399996 187525 400024
rect 176620 399984 176626 399996
rect 187513 399993 187525 399996
rect 187559 399993 187571 400027
rect 187513 399987 187571 399993
rect 187602 399984 187608 400036
rect 187660 399984 187666 400036
rect 187697 400027 187755 400033
rect 187697 399993 187709 400027
rect 187743 400024 187755 400027
rect 198826 400024 198832 400036
rect 187743 399996 198832 400024
rect 187743 399993 187755 399996
rect 187697 399987 187755 399993
rect 198826 399984 198832 399996
rect 198884 399984 198890 400036
rect 184198 399916 184204 399968
rect 184256 399956 184262 399968
rect 217410 399956 217416 399968
rect 184256 399928 217416 399956
rect 184256 399916 184262 399928
rect 217410 399916 217416 399928
rect 217468 399916 217474 399968
rect 115750 399848 115756 399900
rect 115808 399888 115814 399900
rect 206370 399888 206376 399900
rect 115808 399860 206376 399888
rect 115808 399848 115814 399860
rect 206370 399848 206376 399860
rect 206428 399848 206434 399900
rect 217594 399848 217600 399900
rect 217652 399888 217658 399900
rect 226334 399888 226340 399900
rect 217652 399860 226340 399888
rect 217652 399848 217658 399860
rect 226334 399848 226340 399860
rect 226392 399848 226398 399900
rect 119982 399780 119988 399832
rect 120040 399820 120046 399832
rect 214650 399820 214656 399832
rect 120040 399792 214656 399820
rect 120040 399780 120046 399792
rect 214650 399780 214656 399792
rect 214708 399780 214714 399832
rect 217686 399780 217692 399832
rect 217744 399820 217750 399832
rect 230474 399820 230480 399832
rect 217744 399792 230480 399820
rect 217744 399780 217750 399792
rect 230474 399780 230480 399792
rect 230532 399780 230538 399832
rect 113082 399712 113088 399764
rect 113140 399752 113146 399764
rect 215938 399752 215944 399764
rect 113140 399724 215944 399752
rect 113140 399712 113146 399724
rect 215938 399712 215944 399724
rect 215996 399712 216002 399764
rect 217870 399712 217876 399764
rect 217928 399752 217934 399764
rect 233234 399752 233240 399764
rect 217928 399724 233240 399752
rect 217928 399712 217934 399724
rect 233234 399712 233240 399724
rect 233292 399712 233298 399764
rect 52086 399644 52092 399696
rect 52144 399684 52150 399696
rect 198918 399684 198924 399696
rect 52144 399656 198924 399684
rect 52144 399644 52150 399656
rect 198918 399644 198924 399656
rect 198976 399644 198982 399696
rect 199470 399644 199476 399696
rect 199528 399684 199534 399696
rect 232038 399684 232044 399696
rect 199528 399656 232044 399684
rect 199528 399644 199534 399656
rect 232038 399644 232044 399656
rect 232096 399644 232102 399696
rect 56962 399576 56968 399628
rect 57020 399616 57026 399628
rect 231946 399616 231952 399628
rect 57020 399588 231952 399616
rect 57020 399576 57026 399588
rect 231946 399576 231952 399588
rect 232004 399576 232010 399628
rect 59262 399508 59268 399560
rect 59320 399548 59326 399560
rect 122926 399548 122932 399560
rect 59320 399520 122932 399548
rect 59320 399508 59326 399520
rect 122926 399508 122932 399520
rect 122984 399508 122990 399560
rect 180702 399508 180708 399560
rect 180760 399548 180766 399560
rect 357618 399548 357624 399560
rect 180760 399520 357624 399548
rect 180760 399508 180766 399520
rect 357618 399508 357624 399520
rect 357676 399508 357682 399560
rect 51994 399440 52000 399492
rect 52052 399480 52058 399492
rect 358998 399480 359004 399492
rect 52052 399452 359004 399480
rect 52052 399440 52058 399452
rect 358998 399440 359004 399452
rect 359056 399440 359062 399492
rect 57882 398760 57888 398812
rect 57940 398800 57946 398812
rect 210418 398800 210424 398812
rect 57940 398772 210424 398800
rect 57940 398760 57946 398772
rect 210418 398760 210424 398772
rect 210476 398760 210482 398812
rect 218514 398760 218520 398812
rect 218572 398800 218578 398812
rect 219437 398803 219495 398809
rect 219437 398800 219449 398803
rect 218572 398772 219449 398800
rect 218572 398760 218578 398772
rect 219437 398769 219449 398772
rect 219483 398769 219495 398803
rect 219437 398763 219495 398769
rect 219526 398760 219532 398812
rect 219584 398800 219590 398812
rect 224494 398800 224500 398812
rect 219584 398772 224500 398800
rect 219584 398760 219590 398772
rect 224494 398760 224500 398772
rect 224552 398760 224558 398812
rect 218146 398692 218152 398744
rect 218204 398732 218210 398744
rect 219621 398735 219679 398741
rect 218204 398704 219572 398732
rect 218204 398692 218210 398704
rect 219158 398556 219164 398608
rect 219216 398596 219222 398608
rect 219437 398599 219495 398605
rect 219437 398596 219449 398599
rect 219216 398568 219449 398596
rect 219216 398556 219222 398568
rect 219437 398565 219449 398568
rect 219483 398565 219495 398599
rect 219544 398596 219572 398704
rect 219621 398701 219633 398735
rect 219667 398732 219679 398735
rect 227714 398732 227720 398744
rect 219667 398704 227720 398732
rect 219667 398701 219679 398704
rect 219621 398695 219679 398701
rect 227714 398692 227720 398704
rect 227772 398692 227778 398744
rect 219802 398624 219808 398676
rect 219860 398664 219866 398676
rect 229278 398664 229284 398676
rect 219860 398636 229284 398664
rect 219860 398624 219866 398636
rect 229278 398624 229284 398636
rect 229336 398624 229342 398676
rect 226610 398596 226616 398608
rect 219544 398568 226616 398596
rect 219437 398559 219495 398565
rect 226610 398556 226616 398568
rect 226668 398556 226674 398608
rect 219342 398488 219348 398540
rect 219400 398528 219406 398540
rect 219529 398531 219587 398537
rect 219400 398488 219434 398528
rect 219529 398497 219541 398531
rect 219575 398528 219587 398531
rect 226702 398528 226708 398540
rect 219575 398500 226708 398528
rect 219575 398497 219587 398500
rect 219529 398491 219587 398497
rect 226702 398488 226708 398500
rect 226760 398488 226766 398540
rect 219406 398392 219434 398488
rect 219710 398420 219716 398472
rect 219768 398460 219774 398472
rect 229186 398460 229192 398472
rect 219768 398432 229192 398460
rect 219768 398420 219774 398432
rect 229186 398420 229192 398432
rect 229244 398420 229250 398472
rect 219529 398395 219587 398401
rect 219529 398392 219541 398395
rect 219406 398364 219541 398392
rect 219529 398361 219541 398364
rect 219575 398361 219587 398395
rect 219529 398355 219587 398361
rect 219618 398352 219624 398404
rect 219676 398392 219682 398404
rect 229094 398392 229100 398404
rect 219676 398364 229100 398392
rect 219676 398352 219682 398364
rect 229094 398352 229100 398364
rect 229152 398352 229158 398404
rect 185578 398284 185584 398336
rect 185636 398324 185642 398336
rect 196802 398324 196808 398336
rect 185636 398296 196808 398324
rect 185636 398284 185642 398296
rect 196802 398284 196808 398296
rect 196860 398284 196866 398336
rect 218330 398284 218336 398336
rect 218388 398324 218394 398336
rect 227806 398324 227812 398336
rect 218388 398296 227812 398324
rect 218388 398284 218394 398296
rect 227806 398284 227812 398296
rect 227864 398284 227870 398336
rect 177942 398216 177948 398268
rect 178000 398256 178006 398268
rect 210602 398256 210608 398268
rect 178000 398228 210608 398256
rect 178000 398216 178006 398228
rect 210602 398216 210608 398228
rect 210660 398216 210666 398268
rect 218238 398216 218244 398268
rect 218296 398256 218302 398268
rect 228358 398256 228364 398268
rect 218296 398228 228364 398256
rect 218296 398216 218302 398228
rect 228358 398216 228364 398228
rect 228416 398216 228422 398268
rect 169662 398148 169668 398200
rect 169720 398188 169726 398200
rect 210694 398188 210700 398200
rect 169720 398160 210700 398188
rect 169720 398148 169726 398160
rect 210694 398148 210700 398160
rect 210752 398148 210758 398200
rect 218054 398148 218060 398200
rect 218112 398188 218118 398200
rect 228266 398188 228272 398200
rect 218112 398160 228272 398188
rect 218112 398148 218118 398160
rect 228266 398148 228272 398160
rect 228324 398148 228330 398200
rect 122742 398080 122748 398132
rect 122800 398120 122806 398132
rect 196618 398120 196624 398132
rect 122800 398092 196624 398120
rect 122800 398080 122806 398092
rect 196618 398080 196624 398092
rect 196676 398080 196682 398132
rect 217778 398080 217784 398132
rect 217836 398120 217842 398132
rect 228634 398120 228640 398132
rect 217836 398092 228640 398120
rect 217836 398080 217842 398092
rect 228634 398080 228640 398092
rect 228692 398080 228698 398132
rect 219434 398012 219440 398064
rect 219492 398052 219498 398064
rect 226426 398052 226432 398064
rect 219492 398024 226432 398052
rect 219492 398012 219498 398024
rect 226426 398012 226432 398024
rect 226484 398012 226490 398064
rect 218422 397944 218428 397996
rect 218480 397984 218486 397996
rect 226518 397984 226524 397996
rect 218480 397956 226524 397984
rect 218480 397944 218486 397956
rect 226518 397944 226524 397956
rect 226576 397944 226582 397996
rect 219437 397919 219495 397925
rect 219437 397885 219449 397919
rect 219483 397916 219495 397919
rect 228082 397916 228088 397928
rect 219483 397888 228088 397916
rect 219483 397885 219495 397888
rect 219437 397879 219495 397885
rect 228082 397876 228088 397888
rect 228140 397876 228146 397928
rect 218606 397808 218612 397860
rect 218664 397848 218670 397860
rect 225414 397848 225420 397860
rect 218664 397820 225420 397848
rect 218664 397808 218670 397820
rect 225414 397808 225420 397820
rect 225472 397808 225478 397860
rect 219529 397783 219587 397789
rect 219529 397749 219541 397783
rect 219575 397780 219587 397783
rect 228450 397780 228456 397792
rect 219575 397752 228456 397780
rect 219575 397749 219587 397752
rect 219529 397743 219587 397749
rect 228450 397740 228456 397752
rect 228508 397740 228514 397792
rect 3418 397468 3424 397520
rect 3476 397508 3482 397520
rect 143534 397508 143540 397520
rect 3476 397480 143540 397508
rect 3476 397468 3482 397480
rect 143534 397468 143540 397480
rect 143592 397468 143598 397520
rect 81986 397400 81992 397452
rect 82044 397440 82050 397452
rect 224954 397440 224960 397452
rect 82044 397412 224960 397440
rect 82044 397400 82050 397412
rect 224954 397400 224960 397412
rect 225012 397400 225018 397452
rect 85482 397332 85488 397384
rect 85540 397372 85546 397384
rect 229370 397372 229376 397384
rect 85540 397344 229376 397372
rect 85540 397332 85546 397344
rect 229370 397332 229376 397344
rect 229428 397332 229434 397384
rect 61470 397264 61476 397316
rect 61528 397304 61534 397316
rect 278038 397304 278044 397316
rect 61528 397276 278044 397304
rect 61528 397264 61534 397276
rect 278038 397264 278044 397276
rect 278096 397264 278102 397316
rect 58802 397196 58808 397248
rect 58860 397236 58866 397248
rect 109494 397236 109500 397248
rect 58860 397208 109500 397236
rect 58860 397196 58866 397208
rect 109494 397196 109500 397208
rect 109552 397196 109558 397248
rect 111242 397196 111248 397248
rect 111300 397236 111306 397248
rect 137278 397236 137284 397248
rect 111300 397208 137284 397236
rect 111300 397196 111306 397208
rect 137278 397196 137284 397208
rect 137336 397196 137342 397248
rect 238018 397196 238024 397248
rect 238076 397236 238082 397248
rect 239214 397236 239220 397248
rect 238076 397208 239220 397236
rect 238076 397196 238082 397208
rect 239214 397196 239220 397208
rect 239272 397196 239278 397248
rect 291838 397196 291844 397248
rect 291896 397236 291902 397248
rect 298462 397236 298468 397248
rect 291896 397208 298468 397236
rect 291896 397196 291902 397208
rect 298462 397196 298468 397208
rect 298520 397196 298526 397248
rect 88794 397128 88800 397180
rect 88852 397168 88858 397180
rect 94498 397168 94504 397180
rect 88852 397140 94504 397168
rect 88852 397128 88858 397140
rect 94498 397128 94504 397140
rect 94556 397128 94562 397180
rect 106458 397128 106464 397180
rect 106516 397168 106522 397180
rect 134518 397168 134524 397180
rect 106516 397140 134524 397168
rect 106516 397128 106522 397140
rect 134518 397128 134524 397140
rect 134576 397128 134582 397180
rect 177298 397128 177304 397180
rect 177356 397168 177362 397180
rect 237006 397168 237012 397180
rect 177356 397140 237012 397168
rect 177356 397128 177362 397140
rect 237006 397128 237012 397140
rect 237064 397128 237070 397180
rect 58986 397060 58992 397112
rect 59044 397100 59050 397112
rect 99374 397100 99380 397112
rect 59044 397072 99380 397100
rect 59044 397060 59050 397072
rect 99374 397060 99380 397072
rect 99432 397060 99438 397112
rect 104066 397060 104072 397112
rect 104124 397100 104130 397112
rect 108393 397103 108451 397109
rect 108393 397100 108405 397103
rect 104124 397072 108405 397100
rect 104124 397060 104130 397072
rect 108393 397069 108405 397072
rect 108439 397069 108451 397103
rect 108393 397063 108451 397069
rect 113634 397060 113640 397112
rect 113692 397100 113698 397112
rect 170398 397100 170404 397112
rect 113692 397072 170404 397100
rect 113692 397060 113698 397072
rect 170398 397060 170404 397072
rect 170456 397060 170462 397112
rect 184290 397060 184296 397112
rect 184348 397100 184354 397112
rect 247678 397100 247684 397112
rect 184348 397072 247684 397100
rect 184348 397060 184354 397072
rect 247678 397060 247684 397072
rect 247736 397060 247742 397112
rect 80974 396992 80980 397044
rect 81032 397032 81038 397044
rect 142798 397032 142804 397044
rect 81032 397004 142804 397032
rect 81032 396992 81038 397004
rect 142798 396992 142804 397004
rect 142856 396992 142862 397044
rect 173802 396992 173808 397044
rect 173860 397032 173866 397044
rect 238110 397032 238116 397044
rect 173860 397004 238116 397032
rect 173860 396992 173866 397004
rect 238110 396992 238116 397004
rect 238168 396992 238174 397044
rect 90726 396924 90732 396976
rect 90784 396964 90790 396976
rect 187786 396964 187792 396976
rect 90784 396936 187792 396964
rect 90784 396924 90790 396936
rect 187786 396924 187792 396936
rect 187844 396924 187850 396976
rect 196618 396924 196624 396976
rect 196676 396964 196682 396976
rect 251266 396964 251272 396976
rect 196676 396936 251272 396964
rect 196676 396924 196682 396936
rect 251266 396924 251272 396936
rect 251324 396924 251330 396976
rect 58710 396856 58716 396908
rect 58768 396896 58774 396908
rect 112070 396896 112076 396908
rect 58768 396868 112076 396896
rect 58768 396856 58774 396868
rect 112070 396856 112076 396868
rect 112128 396856 112134 396908
rect 115842 396856 115848 396908
rect 115900 396896 115906 396908
rect 224770 396896 224776 396908
rect 115900 396868 224776 396896
rect 115900 396856 115906 396868
rect 224770 396856 224776 396868
rect 224828 396856 224834 396908
rect 58526 396788 58532 396840
rect 58584 396828 58590 396840
rect 113174 396828 113180 396840
rect 58584 396800 113180 396828
rect 58584 396788 58590 396800
rect 113174 396788 113180 396800
rect 113232 396788 113238 396840
rect 118326 396788 118332 396840
rect 118384 396828 118390 396840
rect 233418 396828 233424 396840
rect 118384 396800 233424 396828
rect 118384 396788 118390 396800
rect 233418 396788 233424 396800
rect 233476 396788 233482 396840
rect 58434 396720 58440 396772
rect 58492 396760 58498 396772
rect 113726 396760 113732 396772
rect 58492 396732 113732 396760
rect 58492 396720 58498 396732
rect 113726 396720 113732 396732
rect 113784 396720 113790 396772
rect 117130 396720 117136 396772
rect 117188 396760 117194 396772
rect 233326 396760 233332 396772
rect 117188 396732 233332 396760
rect 117188 396720 117194 396732
rect 233326 396720 233332 396732
rect 233384 396720 233390 396772
rect 240778 396720 240784 396772
rect 240836 396760 240842 396772
rect 242894 396760 242900 396772
rect 240836 396732 242900 396760
rect 240836 396720 240842 396732
rect 242894 396720 242900 396732
rect 242952 396720 242958 396772
rect 249058 396720 249064 396772
rect 249116 396760 249122 396772
rect 256878 396760 256884 396772
rect 249116 396732 256884 396760
rect 249116 396720 249122 396732
rect 256878 396720 256884 396732
rect 256936 396720 256942 396772
rect 268378 396720 268384 396772
rect 268436 396760 268442 396772
rect 273254 396760 273260 396772
rect 268436 396732 273260 396760
rect 268436 396720 268442 396732
rect 273254 396720 273260 396732
rect 273312 396720 273318 396772
rect 287698 396720 287704 396772
rect 287756 396760 287762 396772
rect 295886 396760 295892 396772
rect 287756 396732 295892 396760
rect 287756 396720 287762 396732
rect 295886 396720 295892 396732
rect 295944 396720 295950 396772
rect 307018 396720 307024 396772
rect 307076 396760 307082 396772
rect 307846 396760 307852 396772
rect 307076 396732 307852 396760
rect 307076 396720 307082 396732
rect 307846 396720 307852 396732
rect 307904 396720 307910 396772
rect 96338 396652 96344 396704
rect 96396 396692 96402 396704
rect 97258 396692 97264 396704
rect 96396 396664 97264 396692
rect 96396 396652 96402 396664
rect 97258 396652 97264 396664
rect 97316 396652 97322 396704
rect 105722 396652 105728 396704
rect 105780 396692 105786 396704
rect 108298 396692 108304 396704
rect 105780 396664 108304 396692
rect 105780 396652 105786 396664
rect 108298 396652 108304 396664
rect 108356 396652 108362 396704
rect 108393 396695 108451 396701
rect 108393 396661 108405 396695
rect 108439 396692 108451 396695
rect 231854 396692 231860 396704
rect 108439 396664 231860 396692
rect 108439 396661 108451 396664
rect 108393 396655 108451 396661
rect 231854 396652 231860 396664
rect 231912 396652 231918 396704
rect 253198 396652 253204 396704
rect 253256 396692 253262 396704
rect 254486 396692 254492 396704
rect 253256 396664 254492 396692
rect 253256 396652 253262 396664
rect 254486 396652 254492 396664
rect 254544 396652 254550 396704
rect 260098 396652 260104 396704
rect 260156 396692 260162 396704
rect 260926 396692 260932 396704
rect 260156 396664 260932 396692
rect 260156 396652 260162 396664
rect 260926 396652 260932 396664
rect 260984 396652 260990 396704
rect 291930 396652 291936 396704
rect 291988 396692 291994 396704
rect 292942 396692 292948 396704
rect 291988 396664 292948 396692
rect 291988 396652 291994 396664
rect 292942 396652 292948 396664
rect 293000 396652 293006 396704
rect 304258 396652 304264 396704
rect 304316 396692 304322 396704
rect 305270 396692 305276 396704
rect 304316 396664 305276 396692
rect 304316 396652 304322 396664
rect 305270 396652 305276 396664
rect 305328 396652 305334 396704
rect 309778 396652 309784 396704
rect 309836 396692 309842 396704
rect 315758 396692 315764 396704
rect 309836 396664 315764 396692
rect 309836 396652 309842 396664
rect 315758 396652 315764 396664
rect 315816 396652 315822 396704
rect 322198 396652 322204 396704
rect 322256 396692 322262 396704
rect 323118 396692 323124 396704
rect 322256 396664 323124 396692
rect 322256 396652 322262 396664
rect 323118 396652 323124 396664
rect 323176 396652 323182 396704
rect 58894 396584 58900 396636
rect 58952 396624 58958 396636
rect 95881 396627 95939 396633
rect 95881 396624 95893 396627
rect 58952 396596 95893 396624
rect 58952 396584 58958 396596
rect 95881 396593 95893 396596
rect 95927 396593 95939 396627
rect 95881 396587 95939 396593
rect 95970 396584 95976 396636
rect 96028 396624 96034 396636
rect 97350 396624 97356 396636
rect 96028 396596 97356 396624
rect 96028 396584 96034 396596
rect 97350 396584 97356 396596
rect 97408 396584 97414 396636
rect 102042 396584 102048 396636
rect 102100 396624 102106 396636
rect 229462 396624 229468 396636
rect 102100 396596 229468 396624
rect 102100 396584 102106 396596
rect 229462 396584 229468 396596
rect 229520 396584 229526 396636
rect 92382 396516 92388 396568
rect 92440 396556 92446 396568
rect 227898 396556 227904 396568
rect 92440 396528 227904 396556
rect 92440 396516 92446 396528
rect 227898 396516 227904 396528
rect 227956 396516 227962 396568
rect 246298 396516 246304 396568
rect 246356 396556 246362 396568
rect 262030 396556 262036 396568
rect 246356 396528 262036 396556
rect 246356 396516 246362 396528
rect 262030 396516 262036 396528
rect 262088 396516 262094 396568
rect 59262 396448 59268 396500
rect 59320 396488 59326 396500
rect 87598 396488 87604 396500
rect 59320 396460 87604 396488
rect 59320 396448 59326 396460
rect 87598 396448 87604 396460
rect 87656 396448 87662 396500
rect 95881 396491 95939 396497
rect 95881 396457 95893 396491
rect 95927 396488 95939 396491
rect 100754 396488 100760 396500
rect 95927 396460 100760 396488
rect 95927 396457 95939 396460
rect 95881 396451 95939 396457
rect 100754 396448 100760 396460
rect 100812 396448 100818 396500
rect 222102 396448 222108 396500
rect 222160 396488 222166 396500
rect 276382 396488 276388 396500
rect 222160 396460 276388 396488
rect 222160 396448 222166 396460
rect 276382 396448 276388 396460
rect 276440 396448 276446 396500
rect 59078 396380 59084 396432
rect 59136 396420 59142 396432
rect 94222 396420 94228 396432
rect 59136 396392 94228 396420
rect 59136 396380 59142 396392
rect 94222 396380 94228 396392
rect 94280 396380 94286 396432
rect 97626 396380 97632 396432
rect 97684 396420 97690 396432
rect 106918 396420 106924 396432
rect 97684 396392 106924 396420
rect 97684 396380 97690 396392
rect 106918 396380 106924 396392
rect 106976 396380 106982 396432
rect 220078 396380 220084 396432
rect 220136 396420 220142 396432
rect 273438 396420 273444 396432
rect 220136 396392 273444 396420
rect 220136 396380 220142 396392
rect 273438 396380 273444 396392
rect 273496 396380 273502 396432
rect 78306 396312 78312 396364
rect 78364 396352 78370 396364
rect 222838 396352 222844 396364
rect 78364 396324 222844 396352
rect 78364 396312 78370 396324
rect 222838 396312 222844 396324
rect 222896 396312 222902 396364
rect 224862 396312 224868 396364
rect 224920 396352 224926 396364
rect 278958 396352 278964 396364
rect 224920 396324 278964 396352
rect 224920 396312 224926 396324
rect 278958 396312 278964 396324
rect 279016 396312 279022 396364
rect 59722 396244 59728 396296
rect 59780 396284 59786 396296
rect 235994 396284 236000 396296
rect 59780 396256 236000 396284
rect 59780 396244 59786 396256
rect 235994 396244 236000 396256
rect 236052 396244 236058 396296
rect 238202 396244 238208 396296
rect 238260 396284 238266 396296
rect 272242 396284 272248 396296
rect 238260 396256 272248 396284
rect 238260 396244 238266 396256
rect 272242 396244 272248 396256
rect 272300 396244 272306 396296
rect 282178 396244 282184 396296
rect 282236 396284 282242 396296
rect 325878 396284 325884 396296
rect 282236 396256 325884 396284
rect 282236 396244 282242 396256
rect 325878 396244 325884 396256
rect 325936 396244 325942 396296
rect 59446 396176 59452 396228
rect 59504 396216 59510 396228
rect 240502 396216 240508 396228
rect 59504 396188 240508 396216
rect 59504 396176 59510 396188
rect 240502 396176 240508 396188
rect 240560 396176 240566 396228
rect 242250 396176 242256 396228
rect 242308 396216 242314 396228
rect 259822 396216 259828 396228
rect 242308 396188 259828 396216
rect 242308 396176 242314 396188
rect 259822 396176 259828 396188
rect 259880 396176 259886 396228
rect 284938 396176 284944 396228
rect 284996 396216 285002 396228
rect 289814 396216 289820 396228
rect 284996 396188 289820 396216
rect 284996 396176 285002 396188
rect 289814 396176 289820 396188
rect 289872 396176 289878 396228
rect 59538 396108 59544 396160
rect 59596 396148 59602 396160
rect 252738 396148 252744 396160
rect 59596 396120 252744 396148
rect 59596 396108 59602 396120
rect 252738 396108 252744 396120
rect 252796 396108 252802 396160
rect 316678 396108 316684 396160
rect 316736 396148 316742 396160
rect 343358 396148 343364 396160
rect 316736 396120 343364 396148
rect 316736 396108 316742 396120
rect 343358 396108 343364 396120
rect 343416 396108 343422 396160
rect 83366 396040 83372 396092
rect 83424 396080 83430 396092
rect 87598 396080 87604 396092
rect 83424 396052 87604 396080
rect 83424 396040 83430 396052
rect 87598 396040 87604 396052
rect 87656 396040 87662 396092
rect 242158 395972 242164 396024
rect 242216 396012 242222 396024
rect 247586 396012 247592 396024
rect 242216 395984 247592 396012
rect 242216 395972 242222 395984
rect 247586 395972 247592 395984
rect 247644 395972 247650 396024
rect 163866 395904 163872 395956
rect 163924 395944 163930 395956
rect 222194 395944 222200 395956
rect 163924 395916 222200 395944
rect 163924 395904 163930 395916
rect 222194 395904 222200 395916
rect 222252 395904 222258 395956
rect 156414 395836 156420 395888
rect 156472 395876 156478 395888
rect 215386 395876 215392 395888
rect 156472 395848 215392 395876
rect 156472 395836 156478 395848
rect 215386 395836 215392 395848
rect 215444 395836 215450 395888
rect 179322 395768 179328 395820
rect 179380 395808 179386 395820
rect 241606 395808 241612 395820
rect 179380 395780 241612 395808
rect 179380 395768 179386 395780
rect 241606 395768 241612 395780
rect 241664 395768 241670 395820
rect 146018 395700 146024 395752
rect 146076 395740 146082 395752
rect 209774 395740 209780 395752
rect 146076 395712 209780 395740
rect 146076 395700 146082 395712
rect 209774 395700 209780 395712
rect 209832 395700 209838 395752
rect 235258 395700 235264 395752
rect 235316 395740 235322 395752
rect 249978 395740 249984 395752
rect 235316 395712 249984 395740
rect 235316 395700 235322 395712
rect 249978 395700 249984 395712
rect 250036 395700 250042 395752
rect 191742 395632 191748 395684
rect 191800 395672 191806 395684
rect 268286 395672 268292 395684
rect 191800 395644 268292 395672
rect 191800 395632 191806 395644
rect 268286 395632 268292 395644
rect 268344 395632 268350 395684
rect 118602 395564 118608 395616
rect 118660 395604 118666 395616
rect 197538 395604 197544 395616
rect 118660 395576 197544 395604
rect 118660 395564 118666 395576
rect 197538 395564 197544 395576
rect 197596 395564 197602 395616
rect 231118 395564 231124 395616
rect 231176 395604 231182 395616
rect 265894 395604 265900 395616
rect 231176 395576 265900 395604
rect 231176 395564 231182 395576
rect 265894 395564 265900 395576
rect 265952 395564 265958 395616
rect 54846 395496 54852 395548
rect 54904 395536 54910 395548
rect 138382 395536 138388 395548
rect 54904 395508 138388 395536
rect 54904 395496 54910 395508
rect 138382 395496 138388 395508
rect 138440 395496 138446 395548
rect 183278 395496 183284 395548
rect 183336 395536 183342 395548
rect 185578 395536 185584 395548
rect 183336 395508 185584 395536
rect 183336 395496 183342 395508
rect 185578 395496 185584 395508
rect 185636 395496 185642 395548
rect 195882 395496 195888 395548
rect 195940 395536 195946 395548
rect 276198 395536 276204 395548
rect 195940 395508 276204 395536
rect 195940 395496 195946 395508
rect 276198 395496 276204 395508
rect 276256 395496 276262 395548
rect 51902 395428 51908 395480
rect 51960 395468 51966 395480
rect 91278 395468 91284 395480
rect 51960 395440 91284 395468
rect 51960 395428 51966 395440
rect 91278 395428 91284 395440
rect 91336 395428 91342 395480
rect 136266 395428 136272 395480
rect 136324 395468 136330 395480
rect 227990 395468 227996 395480
rect 136324 395440 227996 395468
rect 136324 395428 136330 395440
rect 227990 395428 227996 395440
rect 228048 395428 228054 395480
rect 238110 395428 238116 395480
rect 238168 395468 238174 395480
rect 273346 395468 273352 395480
rect 238168 395440 273352 395468
rect 238168 395428 238174 395440
rect 273346 395428 273352 395440
rect 273404 395428 273410 395480
rect 54938 395360 54944 395412
rect 54996 395400 55002 395412
rect 123478 395400 123484 395412
rect 54996 395372 123484 395400
rect 54996 395360 55002 395372
rect 123478 395360 123484 395372
rect 123536 395360 123542 395412
rect 125962 395360 125968 395412
rect 126020 395400 126026 395412
rect 228174 395400 228180 395412
rect 126020 395372 228180 395400
rect 126020 395360 126026 395372
rect 228174 395360 228180 395372
rect 228232 395360 228238 395412
rect 232498 395360 232504 395412
rect 232556 395400 232562 395412
rect 270862 395400 270868 395412
rect 232556 395372 270868 395400
rect 232556 395360 232562 395372
rect 270862 395360 270868 395372
rect 270920 395360 270926 395412
rect 85022 395292 85028 395344
rect 85080 395332 85086 395344
rect 233510 395332 233516 395344
rect 85080 395304 233516 395332
rect 85080 395292 85086 395304
rect 233510 395292 233516 395304
rect 233568 395292 233574 395344
rect 240870 395292 240876 395344
rect 240928 395332 240934 395344
rect 283190 395332 283196 395344
rect 240928 395304 283196 395332
rect 240928 395292 240934 395304
rect 283190 395292 283196 395304
rect 283248 395292 283254 395344
rect 180518 393320 180524 393372
rect 180576 393360 180582 393372
rect 183278 393360 183284 393372
rect 180576 393332 183284 393360
rect 180576 393320 180582 393332
rect 183278 393320 183284 393332
rect 183336 393320 183342 393372
rect 177390 388492 177396 388544
rect 177448 388532 177454 388544
rect 180518 388532 180524 388544
rect 177448 388504 180524 388532
rect 177448 388492 177454 388504
rect 180518 388492 180524 388504
rect 180576 388492 180582 388544
rect 85482 378156 85488 378208
rect 85540 378196 85546 378208
rect 580166 378196 580172 378208
rect 85540 378168 580172 378196
rect 85540 378156 85546 378168
rect 580166 378156 580172 378168
rect 580224 378156 580230 378208
rect 175274 377000 175280 377052
rect 175332 377040 175338 377052
rect 177390 377040 177396 377052
rect 175332 377012 177396 377040
rect 175332 377000 175338 377012
rect 177390 377000 177396 377012
rect 177448 377000 177454 377052
rect 171134 375096 171140 375148
rect 171192 375136 171198 375148
rect 175274 375136 175280 375148
rect 171192 375108 175280 375136
rect 171192 375096 171198 375108
rect 175274 375096 175280 375108
rect 175332 375096 175338 375148
rect 171134 372620 171140 372632
rect 171106 372580 171140 372620
rect 171192 372580 171198 372632
rect 164878 372512 164884 372564
rect 164936 372552 164942 372564
rect 171106 372552 171134 372580
rect 164936 372524 171134 372552
rect 164936 372512 164942 372524
rect 3418 371220 3424 371272
rect 3476 371260 3482 371272
rect 144914 371260 144920 371272
rect 3476 371232 144920 371260
rect 3476 371220 3482 371232
rect 144914 371220 144920 371232
rect 144972 371220 144978 371272
rect 154482 367752 154488 367804
rect 154540 367792 154546 367804
rect 228910 367792 228916 367804
rect 154540 367764 228916 367792
rect 154540 367752 154546 367764
rect 228910 367752 228916 367764
rect 228968 367752 228974 367804
rect 85390 364352 85396 364404
rect 85448 364392 85454 364404
rect 579614 364392 579620 364404
rect 85448 364364 579620 364392
rect 85448 364352 85454 364364
rect 579614 364352 579620 364364
rect 579672 364352 579678 364404
rect 160094 359456 160100 359508
rect 160152 359496 160158 359508
rect 164878 359496 164884 359508
rect 160152 359468 164884 359496
rect 160152 359456 160158 359468
rect 164878 359456 164884 359468
rect 164936 359456 164942 359508
rect 54754 358028 54760 358080
rect 54812 358068 54818 358080
rect 147674 358068 147680 358080
rect 54812 358040 147680 358068
rect 54812 358028 54818 358040
rect 147674 358028 147680 358040
rect 147732 358028 147738 358080
rect 3142 357416 3148 357468
rect 3200 357456 3206 357468
rect 147674 357456 147680 357468
rect 3200 357428 147680 357456
rect 3200 357416 3206 357428
rect 147674 357416 147680 357428
rect 147732 357416 147738 357468
rect 159358 357416 159364 357468
rect 159416 357456 159422 357468
rect 160094 357456 160100 357468
rect 159416 357428 160100 357456
rect 159416 357416 159422 357428
rect 160094 357416 160100 357428
rect 160152 357416 160158 357468
rect 84102 351908 84108 351960
rect 84160 351948 84166 351960
rect 580166 351948 580172 351960
rect 84160 351920 580172 351948
rect 84160 351908 84166 351920
rect 580166 351908 580172 351920
rect 580224 351908 580230 351960
rect 156598 346332 156604 346384
rect 156656 346372 156662 346384
rect 159358 346372 159364 346384
rect 156656 346344 159364 346372
rect 156656 346332 156662 346344
rect 159358 346332 159364 346344
rect 159416 346332 159422 346384
rect 3326 345040 3332 345092
rect 3384 345080 3390 345092
rect 146294 345080 146300 345092
rect 3384 345052 146300 345080
rect 3384 345040 3390 345052
rect 146294 345040 146300 345052
rect 146352 345040 146358 345092
rect 81342 324300 81348 324352
rect 81400 324340 81406 324352
rect 580166 324340 580172 324352
rect 81400 324312 580172 324340
rect 81400 324300 81406 324312
rect 580166 324300 580172 324312
rect 580224 324300 580230 324352
rect 3418 318792 3424 318844
rect 3476 318832 3482 318844
rect 147766 318832 147772 318844
rect 3476 318804 147772 318832
rect 3476 318792 3482 318804
rect 147766 318792 147772 318804
rect 147824 318792 147830 318844
rect 154574 311924 154580 311976
rect 154632 311964 154638 311976
rect 156598 311964 156604 311976
rect 154632 311936 156604 311964
rect 154632 311924 154638 311936
rect 156598 311924 156604 311936
rect 156656 311924 156662 311976
rect 82722 311856 82728 311908
rect 82780 311896 82786 311908
rect 579982 311896 579988 311908
rect 82780 311868 579988 311896
rect 82780 311856 82786 311868
rect 579982 311856 579988 311868
rect 580040 311856 580046 311908
rect 151078 306348 151084 306400
rect 151136 306388 151142 306400
rect 154482 306388 154488 306400
rect 151136 306360 154488 306388
rect 151136 306348 151142 306360
rect 154482 306348 154488 306360
rect 154540 306348 154546 306400
rect 3234 304988 3240 305040
rect 3292 305028 3298 305040
rect 150434 305028 150440 305040
rect 3292 305000 150440 305028
rect 3292 304988 3298 305000
rect 150434 304988 150440 305000
rect 150492 304988 150498 305040
rect 149698 299412 149704 299464
rect 149756 299452 149762 299464
rect 151078 299452 151084 299464
rect 149756 299424 151084 299452
rect 149756 299412 149762 299424
rect 151078 299412 151084 299424
rect 151136 299412 151142 299464
rect 81250 298120 81256 298172
rect 81308 298160 81314 298172
rect 580166 298160 580172 298172
rect 81308 298132 580172 298160
rect 81308 298120 81314 298132
rect 580166 298120 580172 298132
rect 580224 298120 580230 298172
rect 3418 292544 3424 292596
rect 3476 292584 3482 292596
rect 149054 292584 149060 292596
rect 3476 292556 149060 292584
rect 3476 292544 3482 292556
rect 149054 292544 149060 292556
rect 149112 292544 149118 292596
rect 148318 282888 148324 282940
rect 148376 282928 148382 282940
rect 149698 282928 149704 282940
rect 148376 282900 149704 282928
rect 148376 282888 148382 282900
rect 149698 282888 149704 282900
rect 149756 282888 149762 282940
rect 78582 271872 78588 271924
rect 78640 271912 78646 271924
rect 580166 271912 580172 271924
rect 78640 271884 580172 271912
rect 78640 271872 78646 271884
rect 580166 271872 580172 271884
rect 580224 271872 580230 271924
rect 146938 271192 146944 271244
rect 146996 271232 147002 271244
rect 148318 271232 148324 271244
rect 146996 271204 148324 271232
rect 146996 271192 147002 271204
rect 148318 271192 148324 271204
rect 148376 271192 148382 271244
rect 151722 266976 151728 267028
rect 151780 267016 151786 267028
rect 212534 267016 212540 267028
rect 151780 266988 212540 267016
rect 151780 266976 151786 266988
rect 212534 266976 212540 266988
rect 212592 266976 212598 267028
rect 150526 266472 150532 266484
rect 142126 266444 150532 266472
rect 3050 266364 3056 266416
rect 3108 266404 3114 266416
rect 142126 266404 142154 266444
rect 150526 266432 150532 266444
rect 150584 266432 150590 266484
rect 3108 266376 142154 266404
rect 3108 266364 3114 266376
rect 145558 266364 145564 266416
rect 145616 266404 145622 266416
rect 146938 266404 146944 266416
rect 145616 266376 146944 266404
rect 145616 266364 145622 266376
rect 146938 266364 146944 266376
rect 146996 266364 147002 266416
rect 144178 262896 144184 262948
rect 144236 262936 144242 262948
rect 145558 262936 145564 262948
rect 144236 262908 145564 262936
rect 144236 262896 144242 262908
rect 145558 262896 145564 262908
rect 145616 262896 145622 262948
rect 104710 261468 104716 261520
rect 104768 261508 104774 261520
rect 229646 261508 229652 261520
rect 104768 261480 229652 261508
rect 104768 261468 104774 261480
rect 229646 261468 229652 261480
rect 229704 261468 229710 261520
rect 112990 258748 112996 258800
rect 113048 258788 113054 258800
rect 360838 258788 360844 258800
rect 113048 258760 360844 258788
rect 113048 258748 113054 258760
rect 360838 258748 360844 258760
rect 360896 258748 360902 258800
rect 107470 258680 107476 258732
rect 107528 258720 107534 258732
rect 376018 258720 376024 258732
rect 107528 258692 376024 258720
rect 107528 258680 107534 258692
rect 376018 258680 376024 258692
rect 376076 258680 376082 258732
rect 79962 258068 79968 258120
rect 80020 258108 80026 258120
rect 580166 258108 580172 258120
rect 80020 258080 580172 258108
rect 80020 258068 80026 258080
rect 580166 258068 580172 258080
rect 580224 258068 580230 258120
rect 142798 256708 142804 256760
rect 142856 256748 142862 256760
rect 144178 256748 144184 256760
rect 142856 256720 144184 256748
rect 142856 256708 142862 256720
rect 144178 256708 144184 256720
rect 144236 256708 144242 256760
rect 3418 253920 3424 253972
rect 3476 253960 3482 253972
rect 153194 253960 153200 253972
rect 3476 253932 153200 253960
rect 3476 253920 3482 253932
rect 153194 253920 153200 253932
rect 153252 253920 153258 253972
rect 141418 251744 141424 251796
rect 141476 251784 141482 251796
rect 142798 251784 142804 251796
rect 141476 251756 142804 251784
rect 141476 251744 141482 251756
rect 142798 251744 142804 251756
rect 142856 251744 142862 251796
rect 232682 250452 232688 250504
rect 232740 250492 232746 250504
rect 317414 250492 317420 250504
rect 232740 250464 317420 250492
rect 232740 250452 232746 250464
rect 317414 250452 317420 250464
rect 317472 250452 317478 250504
rect 142890 249568 142896 249620
rect 142948 249608 142954 249620
rect 226886 249608 226892 249620
rect 142948 249580 226892 249608
rect 142948 249568 142954 249580
rect 226886 249568 226892 249580
rect 226944 249568 226950 249620
rect 94498 249500 94504 249552
rect 94556 249540 94562 249552
rect 180886 249540 180892 249552
rect 94556 249512 180892 249540
rect 94556 249500 94562 249512
rect 180886 249500 180892 249512
rect 180944 249500 180950 249552
rect 97350 249432 97356 249484
rect 97408 249472 97414 249484
rect 195974 249472 195980 249484
rect 97408 249444 195980 249472
rect 97408 249432 97414 249444
rect 195974 249432 195980 249444
rect 196032 249432 196038 249484
rect 108298 249364 108304 249416
rect 108356 249404 108362 249416
rect 207014 249404 207020 249416
rect 108356 249376 207020 249404
rect 108356 249364 108362 249376
rect 207014 249364 207020 249376
rect 207072 249364 207078 249416
rect 119890 249296 119896 249348
rect 119948 249336 119954 249348
rect 223666 249336 223672 249348
rect 119948 249308 223672 249336
rect 119948 249296 119954 249308
rect 223666 249296 223672 249308
rect 223724 249296 223730 249348
rect 99190 249228 99196 249280
rect 99248 249268 99254 249280
rect 225046 249268 225052 249280
rect 99248 249240 225052 249268
rect 99248 249228 99254 249240
rect 225046 249228 225052 249240
rect 225104 249228 225110 249280
rect 99282 249160 99288 249212
rect 99340 249200 99346 249212
rect 230658 249200 230664 249212
rect 99340 249172 230664 249200
rect 99340 249160 99346 249172
rect 230658 249160 230664 249172
rect 230716 249160 230722 249212
rect 77110 249092 77116 249144
rect 77168 249132 77174 249144
rect 233694 249132 233700 249144
rect 77168 249104 233700 249132
rect 77168 249092 77174 249104
rect 233694 249092 233700 249104
rect 233752 249092 233758 249144
rect 51810 249024 51816 249076
rect 51868 249064 51874 249076
rect 259546 249064 259552 249076
rect 51868 249036 259552 249064
rect 51868 249024 51874 249036
rect 259546 249024 259552 249036
rect 259604 249024 259610 249076
rect 54202 248344 54208 248396
rect 54260 248384 54266 248396
rect 129734 248384 129740 248396
rect 54260 248356 129740 248384
rect 54260 248344 54266 248356
rect 129734 248344 129740 248356
rect 129792 248344 129798 248396
rect 97258 248276 97264 248328
rect 97316 248316 97322 248328
rect 176010 248316 176016 248328
rect 97316 248288 176016 248316
rect 97316 248276 97322 248288
rect 176010 248276 176016 248288
rect 176068 248276 176074 248328
rect 111702 248208 111708 248260
rect 111760 248248 111766 248260
rect 193214 248248 193220 248260
rect 111760 248220 193220 248248
rect 111760 248208 111766 248220
rect 193214 248208 193220 248220
rect 193272 248208 193278 248260
rect 106918 248140 106924 248192
rect 106976 248180 106982 248192
rect 198826 248180 198832 248192
rect 106976 248152 198832 248180
rect 106976 248140 106982 248152
rect 198826 248140 198832 248152
rect 198884 248140 198890 248192
rect 87598 248072 87604 248124
rect 87656 248112 87662 248124
rect 171226 248112 171232 248124
rect 87656 248084 171232 248112
rect 87656 248072 87662 248084
rect 171226 248072 171232 248084
rect 171284 248072 171290 248124
rect 193122 248072 193128 248124
rect 193180 248112 193186 248124
rect 316678 248112 316684 248124
rect 193180 248084 316684 248112
rect 193180 248072 193186 248084
rect 316678 248072 316684 248084
rect 316736 248072 316742 248124
rect 101950 248004 101956 248056
rect 102008 248044 102014 248056
rect 229738 248044 229744 248056
rect 102008 248016 229744 248044
rect 102008 248004 102014 248016
rect 229738 248004 229744 248016
rect 229796 248004 229802 248056
rect 47578 247936 47584 247988
rect 47636 247976 47642 247988
rect 142154 247976 142160 247988
rect 47636 247948 142160 247976
rect 47636 247936 47642 247948
rect 142154 247936 142160 247948
rect 142212 247936 142218 247988
rect 188982 247936 188988 247988
rect 189040 247976 189046 247988
rect 342346 247976 342352 247988
rect 189040 247948 342352 247976
rect 189040 247936 189046 247948
rect 342346 247936 342352 247948
rect 342404 247936 342410 247988
rect 51718 247868 51724 247920
rect 51776 247908 51782 247920
rect 265066 247908 265072 247920
rect 51776 247880 265072 247908
rect 51776 247868 51782 247880
rect 265066 247868 265072 247880
rect 265124 247868 265130 247920
rect 54570 247800 54576 247852
rect 54628 247840 54634 247852
rect 277486 247840 277492 247852
rect 54628 247812 277492 247840
rect 54628 247800 54634 247812
rect 277486 247800 277492 247812
rect 277544 247800 277550 247852
rect 55858 247732 55864 247784
rect 55916 247772 55922 247784
rect 310514 247772 310520 247784
rect 55916 247744 310520 247772
rect 55916 247732 55922 247744
rect 310514 247732 310520 247744
rect 310572 247732 310578 247784
rect 88242 247664 88248 247716
rect 88300 247704 88306 247716
rect 580258 247704 580264 247716
rect 88300 247676 580264 247704
rect 88300 247664 88306 247676
rect 580258 247664 580264 247676
rect 580316 247664 580322 247716
rect 120718 247596 120724 247648
rect 120776 247636 120782 247648
rect 196526 247636 196532 247648
rect 120776 247608 196532 247636
rect 120776 247596 120782 247608
rect 196526 247596 196532 247608
rect 196584 247596 196590 247648
rect 32398 246984 32404 247036
rect 32456 247024 32462 247036
rect 140866 247024 140872 247036
rect 32456 246996 140872 247024
rect 32456 246984 32462 246996
rect 140866 246984 140872 246996
rect 140924 246984 140930 247036
rect 161382 246984 161388 247036
rect 161440 247024 161446 247036
rect 233602 247024 233608 247036
rect 161440 246996 233608 247024
rect 161440 246984 161446 246996
rect 233602 246984 233608 246996
rect 233660 246984 233666 247036
rect 108850 246916 108856 246968
rect 108908 246956 108914 246968
rect 229830 246956 229836 246968
rect 108908 246928 229836 246956
rect 108908 246916 108914 246928
rect 229830 246916 229836 246928
rect 229888 246916 229894 246968
rect 91002 246848 91008 246900
rect 91060 246888 91066 246900
rect 228818 246888 228824 246900
rect 91060 246860 228824 246888
rect 91060 246848 91066 246860
rect 228818 246848 228824 246860
rect 228876 246848 228882 246900
rect 54478 246780 54484 246832
rect 54536 246820 54542 246832
rect 280154 246820 280160 246832
rect 54536 246792 280160 246820
rect 54536 246780 54542 246792
rect 280154 246780 280160 246792
rect 280212 246780 280218 246832
rect 54294 246712 54300 246764
rect 54352 246752 54358 246764
rect 287054 246752 287060 246764
rect 54352 246724 287060 246752
rect 54352 246712 54358 246724
rect 287054 246712 287060 246724
rect 287112 246712 287118 246764
rect 108850 246644 108856 246696
rect 108908 246684 108914 246696
rect 388438 246684 388444 246696
rect 108908 246656 388444 246684
rect 108908 246644 108914 246656
rect 388438 246644 388444 246656
rect 388496 246644 388502 246696
rect 100662 246576 100668 246628
rect 100720 246616 100726 246628
rect 382918 246616 382924 246628
rect 100720 246588 382924 246616
rect 100720 246576 100726 246588
rect 382918 246576 382924 246588
rect 382976 246576 382982 246628
rect 103330 246508 103336 246560
rect 103388 246548 103394 246560
rect 385678 246548 385684 246560
rect 103388 246520 385684 246548
rect 103388 246508 103394 246520
rect 385678 246508 385684 246520
rect 385736 246508 385742 246560
rect 88150 246440 88156 246492
rect 88208 246480 88214 246492
rect 378778 246480 378784 246492
rect 88208 246452 378784 246480
rect 88208 246440 88214 246452
rect 378778 246440 378784 246452
rect 378836 246440 378842 246492
rect 111702 246372 111708 246424
rect 111760 246412 111766 246424
rect 412634 246412 412640 246424
rect 111760 246384 412640 246412
rect 111760 246372 111766 246384
rect 412634 246372 412640 246384
rect 412692 246372 412698 246424
rect 106182 246304 106188 246356
rect 106240 246344 106246 246356
rect 542354 246344 542360 246356
rect 106240 246316 542360 246344
rect 106240 246304 106246 246316
rect 542354 246304 542360 246316
rect 542412 246304 542418 246356
rect 35158 246236 35164 246288
rect 35216 246276 35222 246288
rect 132494 246276 132500 246288
rect 35216 246248 132500 246276
rect 35216 246236 35222 246248
rect 132494 246236 132500 246248
rect 132552 246236 132558 246288
rect 133782 246236 133788 246288
rect 133840 246276 133846 246288
rect 228542 246276 228548 246288
rect 133840 246248 228548 246276
rect 133840 246236 133846 246248
rect 228542 246236 228548 246248
rect 228600 246236 228606 246288
rect 33778 246168 33784 246220
rect 33836 246208 33842 246220
rect 126974 246208 126980 246220
rect 33836 246180 126980 246208
rect 33836 246168 33842 246180
rect 126974 246168 126980 246180
rect 127032 246168 127038 246220
rect 137278 246168 137284 246220
rect 137336 246208 137342 246220
rect 212626 246208 212632 246220
rect 137336 246180 212632 246208
rect 137336 246168 137342 246180
rect 212626 246168 212632 246180
rect 212684 246168 212690 246220
rect 36538 246100 36544 246152
rect 36596 246140 36602 246152
rect 129734 246140 129740 246152
rect 36596 246112 129740 246140
rect 36596 246100 36602 246112
rect 129734 246100 129740 246112
rect 129792 246100 129798 246152
rect 55950 246032 55956 246084
rect 56008 246072 56014 246084
rect 140774 246072 140780 246084
rect 56008 246044 140780 246072
rect 56008 246032 56014 246044
rect 140774 246032 140780 246044
rect 140832 246032 140838 246084
rect 56042 245964 56048 246016
rect 56100 246004 56106 246016
rect 120074 246004 120080 246016
rect 56100 245976 120080 246004
rect 56100 245964 56106 245976
rect 120074 245964 120080 245976
rect 120132 245964 120138 246016
rect 141418 245664 141424 245676
rect 139412 245636 141424 245664
rect 22738 245556 22744 245608
rect 22796 245596 22802 245608
rect 129826 245596 129832 245608
rect 22796 245568 129832 245596
rect 22796 245556 22802 245568
rect 129826 245556 129832 245568
rect 129884 245556 129890 245608
rect 138566 245556 138572 245608
rect 138624 245596 138630 245608
rect 139412 245596 139440 245636
rect 141418 245624 141424 245636
rect 141476 245624 141482 245676
rect 138624 245568 139440 245596
rect 138624 245556 138630 245568
rect 183462 245556 183468 245608
rect 183520 245596 183526 245608
rect 232314 245596 232320 245608
rect 183520 245568 232320 245596
rect 183520 245556 183526 245568
rect 232314 245556 232320 245568
rect 232372 245556 232378 245608
rect 8202 245488 8208 245540
rect 8260 245528 8266 245540
rect 127066 245528 127072 245540
rect 8260 245500 127072 245528
rect 8260 245488 8266 245500
rect 127066 245488 127072 245500
rect 127124 245488 127130 245540
rect 134518 245488 134524 245540
rect 134576 245528 134582 245540
rect 208486 245528 208492 245540
rect 134576 245500 208492 245528
rect 134576 245488 134582 245500
rect 208486 245488 208492 245500
rect 208544 245488 208550 245540
rect 106090 245420 106096 245472
rect 106148 245460 106154 245472
rect 228726 245460 228732 245472
rect 106148 245432 228732 245460
rect 106148 245420 106154 245432
rect 228726 245420 228732 245432
rect 228784 245420 228790 245472
rect 18598 245352 18604 245404
rect 18656 245392 18662 245404
rect 142706 245392 142712 245404
rect 18656 245364 142712 245392
rect 18656 245352 18662 245364
rect 142706 245352 142712 245364
rect 142764 245352 142770 245404
rect 206922 245352 206928 245404
rect 206980 245392 206986 245404
rect 287698 245392 287704 245404
rect 206980 245364 287704 245392
rect 206980 245352 206986 245364
rect 287698 245352 287704 245364
rect 287756 245352 287762 245404
rect 4798 245284 4804 245336
rect 4856 245324 4862 245336
rect 138106 245324 138112 245336
rect 4856 245296 138112 245324
rect 4856 245284 4862 245296
rect 138106 245284 138112 245296
rect 138164 245284 138170 245336
rect 186222 245284 186228 245336
rect 186280 245324 186286 245336
rect 357526 245324 357532 245336
rect 186280 245296 357532 245324
rect 186280 245284 186286 245296
rect 357526 245284 357532 245296
rect 357584 245284 357590 245336
rect 51626 245216 51632 245268
rect 51684 245256 51690 245268
rect 266446 245256 266452 245268
rect 51684 245228 266452 245256
rect 51684 245216 51690 245228
rect 266446 245216 266452 245228
rect 266504 245216 266510 245268
rect 110322 245148 110328 245200
rect 110380 245188 110386 245200
rect 377398 245188 377404 245200
rect 110380 245160 377404 245188
rect 110380 245148 110386 245160
rect 377398 245148 377404 245160
rect 377456 245148 377462 245200
rect 104802 245080 104808 245132
rect 104860 245120 104866 245132
rect 374638 245120 374644 245132
rect 104860 245092 374644 245120
rect 104860 245080 104866 245092
rect 374638 245080 374644 245092
rect 374696 245080 374702 245132
rect 99282 245012 99288 245064
rect 99340 245052 99346 245064
rect 370498 245052 370504 245064
rect 99340 245024 370504 245052
rect 99340 245012 99346 245024
rect 370498 245012 370504 245024
rect 370556 245012 370562 245064
rect 93578 244944 93584 244996
rect 93636 244984 93642 244996
rect 381538 244984 381544 244996
rect 93636 244956 381544 244984
rect 93636 244944 93642 244956
rect 381538 244944 381544 244956
rect 381596 244944 381602 244996
rect 91002 244876 91008 244928
rect 91060 244916 91066 244928
rect 443638 244916 443644 244928
rect 91060 244888 443644 244916
rect 91060 244876 91066 244888
rect 443638 244876 443644 244888
rect 443696 244876 443702 244928
rect 25498 244808 25504 244860
rect 25556 244848 25562 244860
rect 132586 244848 132592 244860
rect 25556 244820 132592 244848
rect 25556 244808 25562 244820
rect 132586 244808 132592 244820
rect 132644 244808 132650 244860
rect 199378 244808 199384 244860
rect 199436 244848 199442 244860
rect 232222 244848 232228 244860
rect 199436 244820 232228 244848
rect 199436 244808 199442 244820
rect 232222 244808 232228 244820
rect 232280 244808 232286 244860
rect 29638 244740 29644 244792
rect 29696 244780 29702 244792
rect 135254 244780 135260 244792
rect 29696 244752 135260 244780
rect 29696 244740 29702 244752
rect 135254 244740 135260 244752
rect 135312 244740 135318 244792
rect 117130 244672 117136 244724
rect 117188 244712 117194 244724
rect 213270 244712 213276 244724
rect 117188 244684 213276 244712
rect 117188 244672 117194 244684
rect 213270 244672 213276 244684
rect 213328 244672 213334 244724
rect 50338 244604 50344 244656
rect 50396 244644 50402 244656
rect 145006 244644 145012 244656
rect 50396 244616 145012 244644
rect 50396 244604 50402 244616
rect 145006 244604 145012 244616
rect 145064 244604 145070 244656
rect 43438 244536 43444 244588
rect 43496 244576 43502 244588
rect 138014 244576 138020 244588
rect 43496 244548 138020 244576
rect 43496 244536 43502 244548
rect 138014 244536 138020 244548
rect 138072 244536 138078 244588
rect 173710 244332 173716 244384
rect 173768 244372 173774 244384
rect 177298 244372 177304 244384
rect 173768 244344 177304 244372
rect 173768 244332 173774 244344
rect 177298 244332 177304 244344
rect 177356 244332 177362 244384
rect 78490 244264 78496 244316
rect 78548 244304 78554 244316
rect 579798 244304 579804 244316
rect 78548 244276 579804 244304
rect 78548 244264 78554 244276
rect 579798 244264 579804 244276
rect 579856 244264 579862 244316
rect 11698 244196 11704 244248
rect 11756 244236 11762 244248
rect 128538 244236 128544 244248
rect 11756 244208 128544 244236
rect 11756 244196 11762 244208
rect 128538 244196 128544 244208
rect 128596 244196 128602 244248
rect 158622 244196 158628 244248
rect 158680 244236 158686 244248
rect 218146 244236 218152 244248
rect 158680 244208 218152 244236
rect 158680 244196 158686 244208
rect 218146 244196 218152 244208
rect 218204 244196 218210 244248
rect 15838 244128 15844 244180
rect 15896 244168 15902 244180
rect 137002 244168 137008 244180
rect 15896 244140 137008 244168
rect 15896 244128 15902 244140
rect 137002 244128 137008 244140
rect 137060 244128 137066 244180
rect 205542 244128 205548 244180
rect 205600 244168 205606 244180
rect 291930 244168 291936 244180
rect 205600 244140 291936 244168
rect 205600 244128 205606 244140
rect 291930 244128 291936 244140
rect 291988 244128 291994 244180
rect 17218 244060 17224 244112
rect 17276 244100 17282 244112
rect 139946 244100 139952 244112
rect 17276 244072 139952 244100
rect 17276 244060 17282 244072
rect 139946 244060 139952 244072
rect 140004 244060 140010 244112
rect 209682 244060 209688 244112
rect 209740 244100 209746 244112
rect 302234 244100 302240 244112
rect 209740 244072 302240 244100
rect 209740 244060 209746 244072
rect 302234 244060 302240 244072
rect 302292 244060 302298 244112
rect 54386 243992 54392 244044
rect 54444 244032 54450 244044
rect 285674 244032 285680 244044
rect 54444 244004 285680 244032
rect 54444 243992 54450 244004
rect 285674 243992 285680 244004
rect 285732 243992 285738 244044
rect 102042 243924 102048 243976
rect 102100 243964 102106 243976
rect 371878 243964 371884 243976
rect 102100 243936 371884 243964
rect 102100 243924 102106 243936
rect 371878 243924 371884 243936
rect 371936 243924 371942 243976
rect 96522 243856 96528 243908
rect 96580 243896 96586 243908
rect 367738 243896 367744 243908
rect 96580 243868 367744 243896
rect 96580 243856 96586 243868
rect 367738 243856 367744 243868
rect 367796 243856 367802 243908
rect 90910 243788 90916 243840
rect 90968 243828 90974 243840
rect 363598 243828 363604 243840
rect 90968 243800 363604 243828
rect 90968 243788 90974 243800
rect 363598 243788 363604 243800
rect 363656 243788 363662 243840
rect 108758 243720 108764 243772
rect 108816 243760 108822 243772
rect 429194 243760 429200 243772
rect 108816 243732 429200 243760
rect 108816 243720 108822 243732
rect 429194 243720 429200 243732
rect 429252 243720 429258 243772
rect 93486 243652 93492 243704
rect 93544 243692 93550 243704
rect 431218 243692 431224 243704
rect 93544 243664 431224 243692
rect 93544 243652 93550 243664
rect 431218 243652 431224 243664
rect 431276 243652 431282 243704
rect 86770 243584 86776 243636
rect 86828 243624 86834 243636
rect 425698 243624 425704 243636
rect 86828 243596 425704 243624
rect 86828 243584 86834 243596
rect 425698 243584 425704 243596
rect 425756 243584 425762 243636
rect 96430 243516 96436 243568
rect 96488 243556 96494 243568
rect 449158 243556 449164 243568
rect 96488 243528 449164 243556
rect 96488 243516 96494 243528
rect 449158 243516 449164 243528
rect 449216 243516 449222 243568
rect 21358 243448 21364 243500
rect 21416 243488 21422 243500
rect 134242 243488 134248 243500
rect 21416 243460 134248 243488
rect 21416 243448 21422 243460
rect 134242 243448 134248 243460
rect 134300 243448 134306 243500
rect 135898 243448 135904 243500
rect 135956 243488 135962 243500
rect 138566 243488 138572 243500
rect 135956 243460 138572 243488
rect 135956 243448 135962 243460
rect 138566 243448 138572 243460
rect 138624 243448 138630 243500
rect 204162 243448 204168 243500
rect 204220 243488 204226 243500
rect 242250 243488 242256 243500
rect 204220 243460 242256 243488
rect 204220 243448 204226 243460
rect 242250 243448 242256 243460
rect 242308 243448 242314 243500
rect 97902 243380 97908 243432
rect 97960 243420 97966 243432
rect 209130 243420 209136 243432
rect 97960 243392 209136 243420
rect 97960 243380 97966 243392
rect 209130 243380 209136 243392
rect 209188 243380 209194 243432
rect 95142 243312 95148 243364
rect 95200 243352 95206 243364
rect 206278 243352 206284 243364
rect 95200 243324 206284 243352
rect 95200 243312 95206 243324
rect 206278 243312 206284 243324
rect 206336 243312 206342 243364
rect 56318 243244 56324 243296
rect 56376 243284 56382 243296
rect 165614 243284 165620 243296
rect 56376 243256 165620 243284
rect 56376 243244 56382 243256
rect 165614 243244 165620 243256
rect 165672 243244 165678 243296
rect 39298 243176 39304 243228
rect 39356 243216 39362 243228
rect 135346 243216 135352 243228
rect 39356 243188 135352 243216
rect 39356 243176 39362 243188
rect 135346 243176 135352 243188
rect 135404 243176 135410 243228
rect 41322 243108 41328 243160
rect 41380 243148 41386 243160
rect 125594 243148 125600 243160
rect 41380 243120 125600 243148
rect 41380 243108 41386 243120
rect 125594 243108 125600 243120
rect 125652 243108 125658 243160
rect 118602 243040 118608 243092
rect 118660 243080 118666 243092
rect 201494 243080 201500 243092
rect 118660 243052 201500 243080
rect 118660 243040 118666 243052
rect 201494 243040 201500 243052
rect 201552 243040 201558 243092
rect 115750 242972 115756 243024
rect 115808 243012 115814 243024
rect 197998 243012 198004 243024
rect 115808 242984 198004 243012
rect 115808 242972 115814 242984
rect 197998 242972 198004 242984
rect 198056 242972 198062 243024
rect 117038 242836 117044 242888
rect 117096 242876 117102 242888
rect 226058 242876 226064 242888
rect 117096 242848 226064 242876
rect 117096 242836 117102 242848
rect 226058 242836 226064 242848
rect 226116 242836 226122 242888
rect 103238 242768 103244 242820
rect 103296 242808 103302 242820
rect 214558 242808 214564 242820
rect 103296 242780 214564 242808
rect 103296 242768 103302 242780
rect 214558 242768 214564 242780
rect 214616 242768 214622 242820
rect 92382 242700 92388 242752
rect 92440 242740 92446 242752
rect 204990 242740 204996 242752
rect 92440 242712 204996 242740
rect 92440 242700 92446 242712
rect 204990 242700 204996 242712
rect 205048 242700 205054 242752
rect 57054 242632 57060 242684
rect 57112 242672 57118 242684
rect 169754 242672 169760 242684
rect 57112 242644 169760 242672
rect 57112 242632 57118 242644
rect 169754 242632 169760 242644
rect 169812 242632 169818 242684
rect 206830 242632 206836 242684
rect 206888 242672 206894 242684
rect 263686 242672 263692 242684
rect 206888 242644 263692 242672
rect 206888 242632 206894 242644
rect 263686 242632 263692 242644
rect 263744 242632 263750 242684
rect 100570 242564 100576 242616
rect 100628 242604 100634 242616
rect 213362 242604 213368 242616
rect 100628 242576 213368 242604
rect 100628 242564 100634 242576
rect 213362 242564 213368 242576
rect 213420 242564 213426 242616
rect 14458 242496 14464 242548
rect 14516 242536 14522 242548
rect 131298 242536 131304 242548
rect 14516 242508 131304 242536
rect 14516 242496 14522 242508
rect 131298 242496 131304 242508
rect 131356 242496 131362 242548
rect 170398 242496 170404 242548
rect 170456 242536 170462 242548
rect 194042 242536 194048 242548
rect 170456 242508 194048 242536
rect 170456 242496 170462 242508
rect 194042 242496 194048 242508
rect 194100 242496 194106 242548
rect 204070 242496 204076 242548
rect 204128 242536 204134 242548
rect 284938 242536 284944 242548
rect 204128 242508 284944 242536
rect 204128 242496 204134 242508
rect 284938 242496 284944 242508
rect 284996 242496 285002 242548
rect 57146 242428 57152 242480
rect 57204 242468 57210 242480
rect 183554 242468 183560 242480
rect 57204 242440 183560 242468
rect 57204 242428 57210 242440
rect 183554 242428 183560 242440
rect 183612 242428 183618 242480
rect 219342 242428 219348 242480
rect 219400 242468 219406 242480
rect 320174 242468 320180 242480
rect 219400 242440 320180 242468
rect 219400 242428 219406 242440
rect 320174 242428 320180 242440
rect 320232 242428 320238 242480
rect 93670 242360 93676 242412
rect 93728 242400 93734 242412
rect 230566 242400 230572 242412
rect 93728 242372 230572 242400
rect 93728 242360 93734 242372
rect 230566 242360 230572 242372
rect 230624 242360 230630 242412
rect 58158 242292 58164 242344
rect 58216 242332 58222 242344
rect 266354 242332 266360 242344
rect 58216 242304 266360 242332
rect 58216 242292 58222 242304
rect 266354 242292 266360 242304
rect 266412 242292 266418 242344
rect 89622 242224 89628 242276
rect 89680 242264 89686 242276
rect 358078 242264 358084 242276
rect 89680 242236 358084 242264
rect 89680 242224 89686 242236
rect 358078 242224 358084 242236
rect 358136 242224 358142 242276
rect 56226 242156 56232 242208
rect 56284 242196 56290 242208
rect 88334 242196 88340 242208
rect 56284 242168 88340 242196
rect 56284 242156 56290 242168
rect 88334 242156 88340 242168
rect 88392 242156 88398 242208
rect 106090 242156 106096 242208
rect 106148 242196 106154 242208
rect 446398 242196 446404 242208
rect 106148 242168 446404 242196
rect 106148 242156 106154 242168
rect 446398 242156 446404 242168
rect 446456 242156 446462 242208
rect 129642 242088 129648 242140
rect 129700 242128 129706 242140
rect 225230 242128 225236 242140
rect 129700 242100 225236 242128
rect 129700 242088 129706 242100
rect 225230 242088 225236 242100
rect 225288 242088 225294 242140
rect 114462 242020 114468 242072
rect 114520 242060 114526 242072
rect 209038 242060 209044 242072
rect 114520 242032 209044 242060
rect 114520 242020 114526 242032
rect 209038 242020 209044 242032
rect 209096 242020 209102 242072
rect 118510 241952 118516 242004
rect 118568 241992 118574 242004
rect 204898 241992 204904 242004
rect 118568 241964 204904 241992
rect 118568 241952 118574 241964
rect 204898 241952 204904 241964
rect 204956 241952 204962 242004
rect 144822 241884 144828 241936
rect 144880 241924 144886 241936
rect 225138 241924 225144 241936
rect 144880 241896 225144 241924
rect 144880 241884 144886 241896
rect 225138 241884 225144 241896
rect 225196 241884 225202 241936
rect 75822 241544 75828 241596
rect 75880 241584 75886 241596
rect 242250 241584 242256 241596
rect 75880 241556 242256 241584
rect 75880 241544 75886 241556
rect 242250 241544 242256 241556
rect 242308 241544 242314 241596
rect 72326 241476 72332 241528
rect 72384 241516 72390 241528
rect 240962 241516 240968 241528
rect 72384 241488 240968 241516
rect 72384 241476 72390 241488
rect 240962 241476 240968 241488
rect 241020 241476 241026 241528
rect 57882 241408 57888 241460
rect 57940 241448 57946 241460
rect 58618 241448 58624 241460
rect 57940 241420 58624 241448
rect 57940 241408 57946 241420
rect 58618 241408 58624 241420
rect 58676 241408 58682 241460
rect 107562 241408 107568 241460
rect 107620 241448 107626 241460
rect 230750 241448 230756 241460
rect 107620 241420 230756 241448
rect 107620 241408 107626 241420
rect 230750 241408 230756 241420
rect 230808 241408 230814 241460
rect 58250 241340 58256 241392
rect 58308 241380 58314 241392
rect 181990 241380 181996 241392
rect 58308 241352 181996 241380
rect 58308 241340 58314 241352
rect 181990 241340 181996 241352
rect 182048 241340 182054 241392
rect 182082 241340 182088 241392
rect 182140 241380 182146 241392
rect 184290 241380 184296 241392
rect 182140 241352 184296 241380
rect 182140 241340 182146 241352
rect 184290 241340 184296 241352
rect 184348 241340 184354 241392
rect 190362 241340 190368 241392
rect 190420 241380 190426 241392
rect 196618 241380 196624 241392
rect 190420 241352 196624 241380
rect 190420 241340 190426 241352
rect 196618 241340 196624 241352
rect 196676 241340 196682 241392
rect 198642 241340 198648 241392
rect 198700 241380 198706 241392
rect 249058 241380 249064 241392
rect 198700 241352 249064 241380
rect 198700 241340 198706 241352
rect 249058 241340 249064 241352
rect 249116 241340 249122 241392
rect 103422 241272 103428 241324
rect 103480 241312 103486 241324
rect 229002 241312 229008 241324
rect 103480 241284 229008 241312
rect 103480 241272 103486 241284
rect 229002 241272 229008 241284
rect 229060 241272 229066 241324
rect 93762 241204 93768 241256
rect 93820 241244 93826 241256
rect 225966 241244 225972 241256
rect 93820 241216 225972 241244
rect 93820 241204 93826 241216
rect 225966 241204 225972 241216
rect 226024 241204 226030 241256
rect 59170 241136 59176 241188
rect 59228 241176 59234 241188
rect 198734 241176 198740 241188
rect 59228 241148 198740 241176
rect 59228 241136 59234 241148
rect 198734 241136 198740 241148
rect 198792 241136 198798 241188
rect 201402 241136 201408 241188
rect 201460 241176 201466 241188
rect 258166 241176 258172 241188
rect 201460 241148 258172 241176
rect 201460 241136 201466 241148
rect 258166 241136 258172 241148
rect 258224 241136 258230 241188
rect 86862 241068 86868 241120
rect 86920 241108 86926 241120
rect 232130 241108 232136 241120
rect 86920 241080 232136 241108
rect 86920 241068 86926 241080
rect 232130 241068 232136 241080
rect 232188 241068 232194 241120
rect 77202 241000 77208 241052
rect 77260 241040 77266 241052
rect 226978 241040 226984 241052
rect 77260 241012 226984 241040
rect 77260 241000 77266 241012
rect 226978 241000 226984 241012
rect 227036 241000 227042 241052
rect 57146 240932 57152 240984
rect 57204 240972 57210 240984
rect 210510 240972 210516 240984
rect 57204 240944 210516 240972
rect 57204 240932 57210 240944
rect 210510 240932 210516 240944
rect 210568 240932 210574 240984
rect 235350 240932 235356 240984
rect 235408 240972 235414 240984
rect 270586 240972 270592 240984
rect 235408 240944 270592 240972
rect 235408 240932 235414 240944
rect 270586 240932 270592 240944
rect 270644 240932 270650 240984
rect 54662 240864 54668 240916
rect 54720 240904 54726 240916
rect 244366 240904 244372 240916
rect 54720 240876 244372 240904
rect 54720 240864 54726 240876
rect 244366 240864 244372 240876
rect 244424 240864 244430 240916
rect 53098 240796 53104 240848
rect 53156 240836 53162 240848
rect 249794 240836 249800 240848
rect 53156 240808 249800 240836
rect 53156 240796 53162 240808
rect 249794 240796 249800 240808
rect 249852 240796 249858 240848
rect 59630 240728 59636 240780
rect 59688 240768 59694 240780
rect 274634 240768 274640 240780
rect 59688 240740 274640 240768
rect 59688 240728 59694 240740
rect 274634 240728 274640 240740
rect 274692 240728 274698 240780
rect 108942 240660 108948 240712
rect 109000 240700 109006 240712
rect 226150 240700 226156 240712
rect 109000 240672 226156 240700
rect 109000 240660 109006 240672
rect 226150 240660 226156 240672
rect 226208 240660 226214 240712
rect 215202 240592 215208 240644
rect 215260 240632 215266 240644
rect 238202 240632 238208 240644
rect 215260 240604 238208 240632
rect 215260 240592 215266 240604
rect 238202 240592 238208 240604
rect 238260 240592 238266 240644
rect 3418 240116 3424 240168
rect 3476 240156 3482 240168
rect 106918 240156 106924 240168
rect 3476 240128 106924 240156
rect 3476 240116 3482 240128
rect 106918 240116 106924 240128
rect 106976 240116 106982 240168
rect 217226 240116 217232 240168
rect 217284 240116 217290 240168
rect 226794 240116 226800 240168
rect 226852 240116 226858 240168
rect 217244 240088 217272 240116
rect 226812 240088 226840 240116
rect 217244 240060 226840 240088
rect 56134 227740 56140 227792
rect 56192 227780 56198 227792
rect 59814 227780 59820 227792
rect 56192 227752 59820 227780
rect 56192 227740 56198 227752
rect 59814 227740 59820 227752
rect 59872 227740 59878 227792
rect 244918 225564 244924 225616
rect 244976 225604 244982 225616
rect 255406 225604 255412 225616
rect 244976 225576 255412 225604
rect 244976 225564 244982 225576
rect 255406 225564 255412 225576
rect 255464 225564 255470 225616
rect 3510 215092 3516 215144
rect 3568 215132 3574 215144
rect 7558 215132 7564 215144
rect 3568 215104 7564 215132
rect 3568 215092 3574 215104
rect 7558 215092 7564 215104
rect 7616 215092 7622 215144
rect 242250 206932 242256 206984
rect 242308 206972 242314 206984
rect 580166 206972 580172 206984
rect 242308 206944 580172 206972
rect 242308 206932 242314 206944
rect 580166 206932 580172 206944
rect 580224 206932 580230 206984
rect 3050 202784 3056 202836
rect 3108 202824 3114 202836
rect 29638 202824 29644 202836
rect 3108 202796 29644 202824
rect 3108 202784 3114 202796
rect 29638 202784 29644 202796
rect 29696 202784 29702 202836
rect 57330 201424 57336 201476
rect 57388 201464 57394 201476
rect 58526 201464 58532 201476
rect 57388 201436 58532 201464
rect 57388 201424 57394 201436
rect 58526 201424 58532 201436
rect 58584 201424 58590 201476
rect 55030 198636 55036 198688
rect 55088 198676 55094 198688
rect 57606 198676 57612 198688
rect 55088 198648 57612 198676
rect 55088 198636 55094 198648
rect 57606 198636 57612 198648
rect 57664 198636 57670 198688
rect 55122 195916 55128 195968
rect 55180 195956 55186 195968
rect 57606 195956 57612 195968
rect 55180 195928 57612 195956
rect 55180 195916 55186 195928
rect 57606 195916 57612 195928
rect 57664 195916 57670 195968
rect 278038 193128 278044 193180
rect 278096 193168 278102 193180
rect 580166 193168 580172 193180
rect 278096 193140 580172 193168
rect 278096 193128 278102 193140
rect 580166 193128 580172 193140
rect 580224 193128 580230 193180
rect 54754 190408 54760 190460
rect 54812 190448 54818 190460
rect 57606 190448 57612 190460
rect 54812 190420 57612 190448
rect 54812 190408 54818 190420
rect 57606 190408 57612 190420
rect 57664 190408 57670 190460
rect 2774 188844 2780 188896
rect 2832 188884 2838 188896
rect 4798 188884 4804 188896
rect 2832 188856 4804 188884
rect 2832 188844 2838 188856
rect 4798 188844 4804 188856
rect 4856 188844 4862 188896
rect 53190 184832 53196 184884
rect 53248 184872 53254 184884
rect 57606 184872 57612 184884
rect 53248 184844 57612 184872
rect 53248 184832 53254 184844
rect 57606 184832 57612 184844
rect 57664 184832 57670 184884
rect 50614 183268 50620 183320
rect 50672 183308 50678 183320
rect 57606 183308 57612 183320
rect 50672 183280 57612 183308
rect 50672 183268 50678 183280
rect 57606 183268 57612 183280
rect 57664 183268 57670 183320
rect 51626 180752 51632 180804
rect 51684 180792 51690 180804
rect 56870 180792 56876 180804
rect 51684 180764 56876 180792
rect 51684 180752 51690 180764
rect 56870 180752 56876 180764
rect 56928 180752 56934 180804
rect 54846 172456 54852 172508
rect 54904 172496 54910 172508
rect 57606 172496 57612 172508
rect 54904 172468 57612 172496
rect 54904 172456 54910 172468
rect 57606 172456 57612 172468
rect 57664 172456 57670 172508
rect 51718 169668 51724 169720
rect 51776 169708 51782 169720
rect 57606 169708 57612 169720
rect 51776 169680 57612 169708
rect 51776 169668 51782 169680
rect 57606 169668 57612 169680
rect 57664 169668 57670 169720
rect 53282 166948 53288 167000
rect 53340 166988 53346 167000
rect 57606 166988 57612 167000
rect 53340 166960 57612 166988
rect 53340 166948 53346 166960
rect 57606 166948 57612 166960
rect 57664 166948 57670 167000
rect 240962 166948 240968 167000
rect 241020 166988 241026 167000
rect 580166 166988 580172 167000
rect 241020 166960 580172 166988
rect 241020 166948 241026 166960
rect 580166 166948 580172 166960
rect 580224 166948 580230 167000
rect 3234 164160 3240 164212
rect 3292 164200 3298 164212
rect 11698 164200 11704 164212
rect 3292 164172 11704 164200
rect 3292 164160 3298 164172
rect 11698 164160 11704 164172
rect 11756 164160 11762 164212
rect 53374 163480 53380 163532
rect 53432 163520 53438 163532
rect 57606 163520 57612 163532
rect 53432 163492 57612 163520
rect 53432 163480 53438 163492
rect 57606 163480 57612 163492
rect 57664 163480 57670 163532
rect 54202 161372 54208 161424
rect 54260 161412 54266 161424
rect 57238 161412 57244 161424
rect 54260 161384 57244 161412
rect 54260 161372 54266 161384
rect 57238 161372 57244 161384
rect 57296 161372 57302 161424
rect 54294 158652 54300 158704
rect 54352 158692 54358 158704
rect 57606 158692 57612 158704
rect 54352 158664 57612 158692
rect 54352 158652 54358 158664
rect 57606 158652 57612 158664
rect 57664 158652 57670 158704
rect 57422 155864 57428 155916
rect 57480 155904 57486 155916
rect 58710 155904 58716 155916
rect 57480 155876 58716 155904
rect 57480 155864 57486 155876
rect 58710 155864 58716 155876
rect 58768 155864 58774 155916
rect 53466 153144 53472 153196
rect 53524 153184 53530 153196
rect 57606 153184 57612 153196
rect 53524 153156 57612 153184
rect 53524 153144 53530 153156
rect 57606 153144 57612 153156
rect 57664 153144 57670 153196
rect 3510 150356 3516 150408
rect 3568 150396 3574 150408
rect 18598 150396 18604 150408
rect 3568 150368 18604 150396
rect 3568 150356 3574 150368
rect 18598 150356 18604 150368
rect 18656 150356 18662 150408
rect 54386 150356 54392 150408
rect 54444 150396 54450 150408
rect 57606 150396 57612 150408
rect 54444 150368 57612 150396
rect 54444 150356 54450 150368
rect 57606 150356 57612 150368
rect 57664 150356 57670 150408
rect 51810 144168 51816 144220
rect 51868 144208 51874 144220
rect 57606 144208 57612 144220
rect 51868 144180 57612 144208
rect 51868 144168 51874 144180
rect 57606 144168 57612 144180
rect 57664 144168 57670 144220
rect 54938 142060 54944 142112
rect 54996 142100 55002 142112
rect 57606 142100 57612 142112
rect 54996 142072 57612 142100
rect 54996 142060 55002 142072
rect 57606 142060 57612 142072
rect 57664 142060 57670 142112
rect 410518 139340 410524 139392
rect 410576 139380 410582 139392
rect 580166 139380 580172 139392
rect 410576 139352 580172 139380
rect 410576 139340 410582 139352
rect 580166 139340 580172 139352
rect 580224 139340 580230 139392
rect 3510 137912 3516 137964
rect 3568 137952 3574 137964
rect 15838 137952 15844 137964
rect 3568 137924 15844 137952
rect 3568 137912 3574 137924
rect 15838 137912 15844 137924
rect 15896 137912 15902 137964
rect 54478 136552 54484 136604
rect 54536 136592 54542 136604
rect 57606 136592 57612 136604
rect 54536 136564 57612 136592
rect 54536 136552 54542 136564
rect 57606 136552 57612 136564
rect 57664 136552 57670 136604
rect 53558 133832 53564 133884
rect 53616 133872 53622 133884
rect 57606 133872 57612 133884
rect 53616 133844 57612 133872
rect 53616 133832 53622 133844
rect 57606 133832 57612 133844
rect 57664 133832 57670 133884
rect 54570 132404 54576 132456
rect 54628 132444 54634 132456
rect 57606 132444 57612 132456
rect 54628 132416 57612 132444
rect 54628 132404 54634 132416
rect 57606 132404 57612 132416
rect 57664 132404 57670 132456
rect 271138 126896 271144 126948
rect 271196 126936 271202 126948
rect 580166 126936 580172 126948
rect 271196 126908 580172 126936
rect 271196 126896 271202 126908
rect 580166 126896 580172 126908
rect 580224 126896 580230 126948
rect 52178 118600 52184 118652
rect 52236 118640 52242 118652
rect 57606 118640 57612 118652
rect 52236 118612 57612 118640
rect 52236 118600 52242 118612
rect 57606 118600 57612 118612
rect 57664 118600 57670 118652
rect 51902 115540 51908 115592
rect 51960 115580 51966 115592
rect 57606 115580 57612 115592
rect 51960 115552 57612 115580
rect 51960 115540 51966 115552
rect 57606 115540 57612 115552
rect 57664 115540 57670 115592
rect 3142 111732 3148 111784
rect 3200 111772 3206 111784
rect 14458 111772 14464 111784
rect 3200 111744 14464 111772
rect 3200 111732 3206 111744
rect 14458 111732 14464 111744
rect 14516 111732 14522 111784
rect 53650 110372 53656 110424
rect 53708 110412 53714 110424
rect 57606 110412 57612 110424
rect 53708 110384 57612 110412
rect 53708 110372 53714 110384
rect 57606 110372 57612 110384
rect 57664 110372 57670 110424
rect 50798 107584 50804 107636
rect 50856 107624 50862 107636
rect 57606 107624 57612 107636
rect 50856 107596 57612 107624
rect 50856 107584 50862 107596
rect 57606 107584 57612 107596
rect 57664 107584 57670 107636
rect 53098 104796 53104 104848
rect 53156 104836 53162 104848
rect 57606 104836 57612 104848
rect 53156 104808 57612 104836
rect 53156 104796 53162 104808
rect 57606 104796 57612 104808
rect 57664 104796 57670 104848
rect 51994 102076 52000 102128
rect 52052 102116 52058 102128
rect 57606 102116 57612 102128
rect 52052 102088 57612 102116
rect 52052 102076 52058 102088
rect 57606 102076 57612 102088
rect 57664 102076 57670 102128
rect 302878 100648 302884 100700
rect 302936 100688 302942 100700
rect 580166 100688 580172 100700
rect 302936 100660 580172 100688
rect 302936 100648 302942 100660
rect 580166 100648 580172 100660
rect 580224 100648 580230 100700
rect 3510 97928 3516 97980
rect 3568 97968 3574 97980
rect 25498 97968 25504 97980
rect 3568 97940 25504 97968
rect 3568 97928 3574 97940
rect 25498 97928 25504 97940
rect 25556 97928 25562 97980
rect 53742 90992 53748 91044
rect 53800 91032 53806 91044
rect 57606 91032 57612 91044
rect 53800 91004 57612 91032
rect 53800 90992 53806 91004
rect 57606 90992 57612 91004
rect 57664 90992 57670 91044
rect 52086 88272 52092 88324
rect 52144 88312 52150 88324
rect 57606 88312 57612 88324
rect 52144 88284 57612 88312
rect 52144 88272 52150 88284
rect 57606 88272 57612 88284
rect 57664 88272 57670 88324
rect 3510 85484 3516 85536
rect 3568 85524 3574 85536
rect 17218 85524 17224 85536
rect 3568 85496 17224 85524
rect 3568 85484 3574 85496
rect 17218 85484 17224 85496
rect 17276 85484 17282 85536
rect 50890 85484 50896 85536
rect 50948 85524 50954 85536
rect 57606 85524 57612 85536
rect 50948 85496 57612 85524
rect 50948 85484 50954 85496
rect 57606 85484 57612 85496
rect 57664 85484 57670 85536
rect 50982 79976 50988 80028
rect 51040 80016 51046 80028
rect 57606 80016 57612 80028
rect 51040 79988 57612 80016
rect 51040 79976 51046 79988
rect 57606 79976 57612 79988
rect 57664 79976 57670 80028
rect 54662 78616 54668 78668
rect 54720 78656 54726 78668
rect 57606 78656 57612 78668
rect 54720 78628 57612 78656
rect 54720 78616 54726 78628
rect 57606 78616 57612 78628
rect 57664 78616 57670 78668
rect 52270 75828 52276 75880
rect 52328 75868 52334 75880
rect 57606 75868 57612 75880
rect 52328 75840 57612 75868
rect 52328 75828 52334 75840
rect 57606 75828 57612 75840
rect 57664 75828 57670 75880
rect 3510 71680 3516 71732
rect 3568 71720 3574 71732
rect 21358 71720 21364 71732
rect 3568 71692 21364 71720
rect 3568 71680 3574 71692
rect 21358 71680 21364 71692
rect 21416 71680 21422 71732
rect 52362 70320 52368 70372
rect 52420 70360 52426 70372
rect 57606 70360 57612 70372
rect 52420 70332 57612 70360
rect 52420 70320 52426 70332
rect 57606 70320 57612 70332
rect 57664 70320 57670 70372
rect 295978 60664 295984 60716
rect 296036 60704 296042 60716
rect 580166 60704 580172 60716
rect 296036 60676 580172 60704
rect 296036 60664 296042 60676
rect 580166 60664 580172 60676
rect 580224 60664 580230 60716
rect 58618 60256 58624 60308
rect 58676 60296 58682 60308
rect 59814 60296 59820 60308
rect 58676 60268 59820 60296
rect 58676 60256 58682 60268
rect 59814 60256 59820 60268
rect 59872 60256 59878 60308
rect 223684 59928 233372 59956
rect 223684 59900 223712 59928
rect 233344 59900 233372 59928
rect 223666 59848 223672 59900
rect 223724 59848 223730 59900
rect 224218 59848 224224 59900
rect 224276 59888 224282 59900
rect 233234 59888 233240 59900
rect 224276 59860 233240 59888
rect 224276 59848 224282 59860
rect 233234 59848 233240 59860
rect 233292 59848 233298 59900
rect 233326 59848 233332 59900
rect 233384 59848 233390 59900
rect 209682 59780 209688 59832
rect 209740 59820 209746 59832
rect 252646 59820 252652 59832
rect 209740 59792 252652 59820
rect 209740 59780 209746 59792
rect 252646 59780 252652 59792
rect 252704 59780 252710 59832
rect 212626 59712 212632 59764
rect 212684 59752 212690 59764
rect 258074 59752 258080 59764
rect 212684 59724 258080 59752
rect 212684 59712 212690 59724
rect 258074 59712 258080 59724
rect 258132 59712 258138 59764
rect 219158 59644 219164 59696
rect 219216 59684 219222 59696
rect 291838 59684 291844 59696
rect 219216 59656 291844 59684
rect 219216 59644 219222 59656
rect 291838 59644 291844 59656
rect 291896 59644 291902 59696
rect 220998 59576 221004 59628
rect 221056 59616 221062 59628
rect 304258 59616 304264 59628
rect 221056 59588 304264 59616
rect 221056 59576 221062 59588
rect 304258 59576 304264 59588
rect 304316 59576 304322 59628
rect 222470 59508 222476 59560
rect 222528 59548 222534 59560
rect 309778 59548 309784 59560
rect 222528 59520 309784 59548
rect 222528 59508 222534 59520
rect 309778 59508 309784 59520
rect 309836 59508 309842 59560
rect 221826 59440 221832 59492
rect 221884 59480 221890 59492
rect 313274 59480 313280 59492
rect 221884 59452 313280 59480
rect 221884 59440 221890 59452
rect 313274 59440 313280 59452
rect 313332 59440 313338 59492
rect 223942 59372 223948 59424
rect 224000 59412 224006 59424
rect 322198 59412 322204 59424
rect 224000 59384 322204 59412
rect 224000 59372 224006 59384
rect 322198 59372 322204 59384
rect 322256 59372 322262 59424
rect 3050 59304 3056 59356
rect 3108 59344 3114 59356
rect 36538 59344 36544 59356
rect 3108 59316 36544 59344
rect 3108 59304 3114 59316
rect 36538 59304 36544 59316
rect 36596 59304 36602 59356
rect 50706 59304 50712 59356
rect 50764 59344 50770 59356
rect 211982 59344 211988 59356
rect 50764 59316 211988 59344
rect 50764 59304 50770 59316
rect 211982 59304 211988 59316
rect 212040 59304 212046 59356
rect 215938 59304 215944 59356
rect 215996 59344 216002 59356
rect 227898 59344 227904 59356
rect 215996 59316 227904 59344
rect 215996 59304 216002 59316
rect 227898 59304 227904 59316
rect 227956 59304 227962 59356
rect 217134 59236 217140 59288
rect 217192 59276 217198 59288
rect 227806 59276 227812 59288
rect 217192 59248 227812 59276
rect 217192 59236 217198 59248
rect 227806 59236 227812 59248
rect 227864 59236 227870 59288
rect 213178 59168 213184 59220
rect 213236 59208 213242 59220
rect 221185 59211 221243 59217
rect 221185 59208 221197 59211
rect 213236 59180 221197 59208
rect 213236 59168 213242 59180
rect 221185 59177 221197 59180
rect 221231 59177 221243 59211
rect 221185 59171 221243 59177
rect 221274 59168 221280 59220
rect 221332 59208 221338 59220
rect 269114 59208 269120 59220
rect 221332 59180 269120 59208
rect 221332 59168 221338 59180
rect 269114 59168 269120 59180
rect 269172 59168 269178 59220
rect 218606 59100 218612 59152
rect 218664 59140 218670 59152
rect 231854 59140 231860 59152
rect 218664 59112 231860 59140
rect 218664 59100 218670 59112
rect 231854 59100 231860 59112
rect 231912 59100 231918 59152
rect 222194 59032 222200 59084
rect 222252 59072 222258 59084
rect 268378 59072 268384 59084
rect 222252 59044 268384 59072
rect 222252 59032 222258 59044
rect 268378 59032 268384 59044
rect 268436 59032 268442 59084
rect 219802 58964 219808 59016
rect 219860 59004 219866 59016
rect 229094 59004 229100 59016
rect 219860 58976 229100 59004
rect 219860 58964 219866 58976
rect 229094 58964 229100 58976
rect 229152 58964 229158 59016
rect 214098 58896 214104 58948
rect 214156 58936 214162 58948
rect 248414 58936 248420 58948
rect 214156 58908 248420 58936
rect 214156 58896 214162 58908
rect 248414 58896 248420 58908
rect 248472 58896 248478 58948
rect 211706 58828 211712 58880
rect 211764 58868 211770 58880
rect 245654 58868 245660 58880
rect 211764 58840 245660 58868
rect 211764 58828 211770 58840
rect 245654 58828 245660 58840
rect 245712 58828 245718 58880
rect 207842 58760 207848 58812
rect 207900 58800 207906 58812
rect 240778 58800 240784 58812
rect 207900 58772 240784 58800
rect 207900 58760 207906 58772
rect 240778 58760 240784 58772
rect 240836 58760 240842 58812
rect 217686 58692 217692 58744
rect 217744 58732 217750 58744
rect 229462 58732 229468 58744
rect 217744 58704 229468 58732
rect 217744 58692 217750 58704
rect 229462 58692 229468 58704
rect 229520 58692 229526 58744
rect 211430 58624 211436 58676
rect 211488 58664 211494 58676
rect 358906 58664 358912 58676
rect 211488 58636 358912 58664
rect 211488 58624 211494 58636
rect 358906 58624 358912 58636
rect 358964 58624 358970 58676
rect 209038 58556 209044 58608
rect 209096 58596 209102 58608
rect 238018 58596 238024 58608
rect 209096 58568 238024 58596
rect 209096 58556 209102 58568
rect 238018 58556 238024 58568
rect 238076 58556 238082 58608
rect 208118 58488 208124 58540
rect 208176 58528 208182 58540
rect 229278 58528 229284 58540
rect 208176 58500 229284 58528
rect 208176 58488 208182 58500
rect 229278 58488 229284 58500
rect 229336 58488 229342 58540
rect 210510 58420 210516 58472
rect 210568 58460 210574 58472
rect 229370 58460 229376 58472
rect 210568 58432 229376 58460
rect 210568 58420 210574 58432
rect 229370 58420 229376 58432
rect 229428 58420 229434 58472
rect 221185 58395 221243 58401
rect 221185 58361 221197 58395
rect 221231 58392 221243 58395
rect 260098 58392 260104 58404
rect 221231 58364 260104 58392
rect 221231 58361 221243 58364
rect 221185 58355 221243 58361
rect 260098 58352 260104 58364
rect 260156 58352 260162 58404
rect 213546 58284 213552 58336
rect 213604 58324 213610 58336
rect 229186 58324 229192 58336
rect 213604 58296 229192 58324
rect 213604 58284 213610 58296
rect 229186 58284 229192 58296
rect 229244 58284 229250 58336
rect 214374 58216 214380 58268
rect 214432 58256 214438 58268
rect 263594 58256 263600 58268
rect 214432 58228 263600 58256
rect 214432 58216 214438 58228
rect 263594 58216 263600 58228
rect 263652 58216 263658 58268
rect 215570 58148 215576 58200
rect 215628 58188 215634 58200
rect 251174 58188 251180 58200
rect 215628 58160 251180 58188
rect 215628 58148 215634 58160
rect 251174 58148 251180 58160
rect 251232 58148 251238 58200
rect 216766 58080 216772 58132
rect 216824 58120 216830 58132
rect 227714 58120 227720 58132
rect 216824 58092 227720 58120
rect 216824 58080 216830 58092
rect 227714 58080 227720 58092
rect 227772 58080 227778 58132
rect 216214 58012 216220 58064
rect 216272 58052 216278 58064
rect 224494 58052 224500 58064
rect 216272 58024 224500 58052
rect 216272 58012 216278 58024
rect 224494 58012 224500 58024
rect 224552 58012 224558 58064
rect 64506 57984 64512 57996
rect 64467 57956 64512 57984
rect 64506 57944 64512 57956
rect 64564 57944 64570 57996
rect 70857 57987 70915 57993
rect 70857 57984 70869 57987
rect 68204 57956 70869 57984
rect 66898 57916 66904 57928
rect 45526 57888 66904 57916
rect 28902 57808 28908 57860
rect 28960 57848 28966 57860
rect 45526 57848 45554 57888
rect 66898 57876 66904 57888
rect 66956 57876 66962 57928
rect 66993 57919 67051 57925
rect 66993 57885 67005 57919
rect 67039 57916 67051 57919
rect 68204 57916 68232 57956
rect 70857 57953 70869 57956
rect 70903 57953 70915 57987
rect 70857 57947 70915 57953
rect 67039 57888 68232 57916
rect 67039 57885 67051 57888
rect 66993 57879 67051 57885
rect 68278 57876 68284 57928
rect 68336 57916 68342 57928
rect 74074 57916 74080 57928
rect 68336 57888 74080 57916
rect 68336 57876 68342 57888
rect 74074 57876 74080 57888
rect 74132 57876 74138 57928
rect 209314 57916 209320 57928
rect 74506 57888 209320 57916
rect 28960 57820 45554 57848
rect 28960 57808 28966 57820
rect 58342 57808 58348 57860
rect 58400 57848 58406 57860
rect 74506 57848 74534 57888
rect 209314 57876 209320 57888
rect 209372 57876 209378 57928
rect 220078 57876 220084 57928
rect 220136 57916 220142 57928
rect 224678 57916 224684 57928
rect 220136 57888 224684 57916
rect 220136 57876 220142 57888
rect 224678 57876 224684 57888
rect 224736 57876 224742 57928
rect 58400 57820 74534 57848
rect 58400 57808 58406 57820
rect 87138 57808 87144 57860
rect 87196 57848 87202 57860
rect 105446 57848 105452 57860
rect 87196 57820 105452 57848
rect 87196 57808 87202 57820
rect 105446 57808 105452 57820
rect 105504 57808 105510 57860
rect 106274 57808 106280 57860
rect 106332 57848 106338 57860
rect 107562 57848 107568 57860
rect 106332 57820 107568 57848
rect 106332 57808 106338 57820
rect 107562 57808 107568 57820
rect 107620 57808 107626 57860
rect 109494 57808 109500 57860
rect 109552 57848 109558 57860
rect 110322 57848 110328 57860
rect 109552 57820 110328 57848
rect 109552 57808 109558 57820
rect 110322 57808 110328 57820
rect 110380 57808 110386 57860
rect 110509 57851 110567 57857
rect 110509 57817 110521 57851
rect 110555 57848 110567 57851
rect 133138 57848 133144 57860
rect 110555 57820 133144 57848
rect 110555 57817 110567 57820
rect 110509 57811 110567 57817
rect 133138 57808 133144 57820
rect 133196 57808 133202 57860
rect 136726 57848 136732 57860
rect 135180 57820 136732 57848
rect 26142 57740 26148 57792
rect 26200 57780 26206 57792
rect 66346 57780 66352 57792
rect 26200 57752 66352 57780
rect 26200 57740 26206 57752
rect 66346 57740 66352 57752
rect 66404 57740 66410 57792
rect 67082 57740 67088 57792
rect 67140 57780 67146 57792
rect 70762 57780 70768 57792
rect 67140 57752 70768 57780
rect 67140 57740 67146 57752
rect 70762 57740 70768 57752
rect 70820 57740 70826 57792
rect 70857 57783 70915 57789
rect 70857 57749 70869 57783
rect 70903 57780 70915 57783
rect 74350 57780 74356 57792
rect 70903 57752 74356 57780
rect 70903 57749 70915 57752
rect 70857 57743 70915 57749
rect 74350 57740 74356 57752
rect 74408 57740 74414 57792
rect 101490 57740 101496 57792
rect 101548 57780 101554 57792
rect 102873 57783 102931 57789
rect 101548 57752 102824 57780
rect 101548 57740 101554 57752
rect 24762 57672 24768 57724
rect 24820 57712 24826 57724
rect 65978 57712 65984 57724
rect 24820 57684 65984 57712
rect 24820 57672 24826 57684
rect 65978 57672 65984 57684
rect 66036 57672 66042 57724
rect 66070 57672 66076 57724
rect 66128 57712 66134 57724
rect 66622 57712 66628 57724
rect 66128 57684 66628 57712
rect 66128 57672 66134 57684
rect 66622 57672 66628 57684
rect 66680 57672 66686 57724
rect 66717 57715 66775 57721
rect 66717 57681 66729 57715
rect 66763 57712 66775 57715
rect 69109 57715 69167 57721
rect 69109 57712 69121 57715
rect 66763 57684 69121 57712
rect 66763 57681 66775 57684
rect 66717 57675 66775 57681
rect 69109 57681 69121 57684
rect 69155 57681 69167 57715
rect 69109 57675 69167 57681
rect 70302 57672 70308 57724
rect 70360 57712 70366 57724
rect 77662 57712 77668 57724
rect 70360 57684 77668 57712
rect 70360 57672 70366 57684
rect 77662 57672 77668 57684
rect 77720 57672 77726 57724
rect 90542 57672 90548 57724
rect 90600 57712 90606 57724
rect 91002 57712 91008 57724
rect 90600 57684 91008 57712
rect 90600 57672 90606 57684
rect 91002 57672 91008 57684
rect 91060 57672 91066 57724
rect 91646 57672 91652 57724
rect 91704 57712 91710 57724
rect 91704 57684 93854 57712
rect 91704 57672 91710 57684
rect 19242 57604 19248 57656
rect 19300 57644 19306 57656
rect 64509 57647 64567 57653
rect 64509 57644 64521 57647
rect 19300 57616 64521 57644
rect 19300 57604 19306 57616
rect 64509 57613 64521 57616
rect 64555 57613 64567 57647
rect 69566 57644 69572 57656
rect 64509 57607 64567 57613
rect 64846 57616 69572 57644
rect 16482 57536 16488 57588
rect 16540 57576 16546 57588
rect 63586 57576 63592 57588
rect 16540 57548 63592 57576
rect 16540 57536 16546 57548
rect 63586 57536 63592 57548
rect 63644 57536 63650 57588
rect 64846 57576 64874 57616
rect 69566 57604 69572 57616
rect 69624 57604 69630 57656
rect 70210 57604 70216 57656
rect 70268 57644 70274 57656
rect 77294 57644 77300 57656
rect 70268 57616 77300 57644
rect 70268 57604 70274 57616
rect 77294 57604 77300 57616
rect 77352 57604 77358 57656
rect 78766 57604 78772 57656
rect 78824 57644 78830 57656
rect 79502 57644 79508 57656
rect 78824 57616 79508 57644
rect 78824 57604 78830 57616
rect 79502 57604 79508 57616
rect 79560 57604 79566 57656
rect 92842 57604 92848 57656
rect 92900 57644 92906 57656
rect 93578 57644 93584 57656
rect 92900 57616 93584 57644
rect 92900 57604 92906 57616
rect 93578 57604 93584 57616
rect 93636 57604 93642 57656
rect 93826 57644 93854 57684
rect 94314 57672 94320 57724
rect 94372 57712 94378 57724
rect 95142 57712 95148 57724
rect 94372 57684 95148 57712
rect 94372 57672 94378 57684
rect 95142 57672 95148 57684
rect 95200 57672 95206 57724
rect 95786 57672 95792 57724
rect 95844 57712 95850 57724
rect 97534 57712 97540 57724
rect 95844 57684 97540 57712
rect 95844 57672 95850 57684
rect 97534 57672 97540 57684
rect 97592 57672 97598 57724
rect 99650 57672 99656 57724
rect 99708 57712 99714 57724
rect 100570 57712 100576 57724
rect 99708 57684 100576 57712
rect 99708 57672 99714 57684
rect 100570 57672 100576 57684
rect 100628 57672 100634 57724
rect 101214 57672 101220 57724
rect 101272 57712 101278 57724
rect 101858 57712 101864 57724
rect 101272 57684 101864 57712
rect 101272 57672 101278 57684
rect 101858 57672 101864 57684
rect 101916 57672 101922 57724
rect 102796 57712 102824 57752
rect 102873 57749 102885 57783
rect 102919 57780 102931 57783
rect 123297 57783 123355 57789
rect 123297 57780 123309 57783
rect 102919 57752 123309 57780
rect 102919 57749 102931 57752
rect 102873 57743 102931 57749
rect 123297 57749 123309 57752
rect 123343 57749 123355 57783
rect 124858 57780 124864 57792
rect 123297 57743 123355 57749
rect 123404 57752 124864 57780
rect 122837 57715 122895 57721
rect 122837 57712 122849 57715
rect 102796 57684 122849 57712
rect 122837 57681 122849 57684
rect 122883 57681 122895 57715
rect 122837 57675 122895 57681
rect 123404 57644 123432 57752
rect 124858 57740 124864 57752
rect 124916 57740 124922 57792
rect 125594 57740 125600 57792
rect 125652 57780 125658 57792
rect 126882 57780 126888 57792
rect 125652 57752 126888 57780
rect 125652 57740 125658 57752
rect 126882 57740 126888 57752
rect 126940 57740 126946 57792
rect 127434 57740 127440 57792
rect 127492 57780 127498 57792
rect 128170 57780 128176 57792
rect 127492 57752 128176 57780
rect 127492 57740 127498 57752
rect 128170 57740 128176 57752
rect 128228 57740 128234 57792
rect 131574 57740 131580 57792
rect 131632 57780 131638 57792
rect 135180 57780 135208 57820
rect 136726 57808 136732 57820
rect 136784 57808 136790 57860
rect 138106 57808 138112 57860
rect 138164 57848 138170 57860
rect 138164 57820 138704 57848
rect 138164 57808 138170 57820
rect 131632 57752 135208 57780
rect 131632 57740 131638 57752
rect 135990 57740 135996 57792
rect 136048 57780 136054 57792
rect 138676 57780 138704 57820
rect 138750 57808 138756 57860
rect 138808 57848 138814 57860
rect 149333 57851 149391 57857
rect 149333 57848 149345 57851
rect 138808 57820 149345 57848
rect 138808 57808 138814 57820
rect 149333 57817 149345 57820
rect 149379 57817 149391 57851
rect 149333 57811 149391 57817
rect 149422 57808 149428 57860
rect 149480 57848 149486 57860
rect 152369 57851 152427 57857
rect 152369 57848 152381 57851
rect 149480 57820 152381 57848
rect 149480 57808 149486 57820
rect 152369 57817 152381 57820
rect 152415 57817 152427 57851
rect 152369 57811 152427 57817
rect 152461 57851 152519 57857
rect 152461 57817 152473 57851
rect 152507 57848 152519 57851
rect 161566 57848 161572 57860
rect 152507 57820 161572 57848
rect 152507 57817 152519 57820
rect 152461 57811 152519 57817
rect 161566 57808 161572 57820
rect 161624 57808 161630 57860
rect 161934 57808 161940 57860
rect 161992 57848 161998 57860
rect 168285 57851 168343 57857
rect 168285 57848 168297 57851
rect 161992 57820 168297 57848
rect 161992 57808 161998 57820
rect 168285 57817 168297 57820
rect 168331 57817 168343 57851
rect 168285 57811 168343 57817
rect 170306 57808 170312 57860
rect 170364 57848 170370 57860
rect 170950 57848 170956 57860
rect 170364 57820 170956 57848
rect 170364 57808 170370 57820
rect 170950 57808 170956 57820
rect 171008 57808 171014 57860
rect 171045 57851 171103 57857
rect 171045 57817 171057 57851
rect 171091 57848 171103 57851
rect 201773 57851 201831 57857
rect 201773 57848 201785 57851
rect 171091 57820 201785 57848
rect 171091 57817 171103 57820
rect 171045 57811 171103 57817
rect 201773 57817 201785 57820
rect 201819 57817 201831 57851
rect 201773 57811 201831 57817
rect 201862 57808 201868 57860
rect 201920 57848 201926 57860
rect 202598 57848 202604 57860
rect 201920 57820 202604 57848
rect 201920 57808 201926 57820
rect 202598 57808 202604 57820
rect 202656 57808 202662 57860
rect 203702 57808 203708 57860
rect 203760 57848 203766 57860
rect 204070 57848 204076 57860
rect 203760 57820 204076 57848
rect 203760 57808 203766 57820
rect 204070 57808 204076 57820
rect 204128 57808 204134 57860
rect 204530 57808 204536 57860
rect 204588 57848 204594 57860
rect 205358 57848 205364 57860
rect 204588 57820 205364 57848
rect 204588 57808 204594 57820
rect 205358 57808 205364 57820
rect 205416 57808 205422 57860
rect 206094 57808 206100 57860
rect 206152 57848 206158 57860
rect 206922 57848 206928 57860
rect 206152 57820 206928 57848
rect 206152 57808 206158 57820
rect 206922 57808 206928 57820
rect 206980 57808 206986 57860
rect 220354 57808 220360 57860
rect 220412 57848 220418 57860
rect 225138 57848 225144 57860
rect 220412 57820 225144 57848
rect 220412 57808 220418 57820
rect 225138 57808 225144 57820
rect 225196 57808 225202 57860
rect 140314 57780 140320 57792
rect 136048 57752 138336 57780
rect 138676 57752 140320 57780
rect 136048 57740 136054 57752
rect 125870 57672 125876 57724
rect 125928 57712 125934 57724
rect 126698 57712 126704 57724
rect 125928 57684 126704 57712
rect 125928 57672 125934 57684
rect 126698 57672 126704 57684
rect 126756 57672 126762 57724
rect 127710 57672 127716 57724
rect 127768 57712 127774 57724
rect 128078 57712 128084 57724
rect 127768 57684 128084 57712
rect 127768 57672 127774 57684
rect 128078 57672 128084 57684
rect 128136 57672 128142 57724
rect 130102 57672 130108 57724
rect 130160 57712 130166 57724
rect 130930 57712 130936 57724
rect 130160 57684 130936 57712
rect 130160 57672 130166 57684
rect 130930 57672 130936 57684
rect 130988 57672 130994 57724
rect 131298 57672 131304 57724
rect 131356 57712 131362 57724
rect 132218 57712 132224 57724
rect 131356 57684 132224 57712
rect 131356 57672 131362 57684
rect 132218 57672 132224 57684
rect 132276 57672 132282 57724
rect 132494 57672 132500 57724
rect 132552 57712 132558 57724
rect 132552 57684 136588 57712
rect 132552 57672 132558 57684
rect 93826 57616 123432 57644
rect 123478 57604 123484 57656
rect 123536 57644 123542 57656
rect 123938 57644 123944 57656
rect 123536 57616 123944 57644
rect 123536 57604 123542 57616
rect 123938 57604 123944 57616
rect 123996 57604 124002 57656
rect 126514 57604 126520 57656
rect 126572 57644 126578 57656
rect 126790 57644 126796 57656
rect 126572 57616 126796 57644
rect 126572 57604 126578 57616
rect 126790 57604 126796 57616
rect 126848 57604 126854 57656
rect 127066 57604 127072 57656
rect 127124 57644 127130 57656
rect 127894 57644 127900 57656
rect 127124 57616 127900 57644
rect 127124 57604 127130 57616
rect 127894 57604 127900 57616
rect 127952 57604 127958 57656
rect 128630 57604 128636 57656
rect 128688 57644 128694 57656
rect 129550 57644 129556 57656
rect 128688 57616 129556 57644
rect 128688 57604 128694 57616
rect 129550 57604 129556 57616
rect 129608 57604 129614 57656
rect 130378 57604 130384 57656
rect 130436 57644 130442 57656
rect 130838 57644 130844 57656
rect 130436 57616 130844 57644
rect 130436 57604 130442 57616
rect 130838 57604 130844 57616
rect 130896 57604 130902 57656
rect 131850 57604 131856 57656
rect 131908 57644 131914 57656
rect 132402 57644 132408 57656
rect 131908 57616 132408 57644
rect 131908 57604 131914 57616
rect 132402 57604 132408 57616
rect 132460 57604 132466 57656
rect 132770 57604 132776 57656
rect 132828 57644 132834 57656
rect 133690 57644 133696 57656
rect 132828 57616 133696 57644
rect 132828 57604 132834 57616
rect 133690 57604 133696 57616
rect 133748 57604 133754 57656
rect 135073 57647 135131 57653
rect 135073 57644 135085 57647
rect 134444 57616 135085 57644
rect 64156 57548 64874 57576
rect 64156 57520 64184 57548
rect 65610 57536 65616 57588
rect 65668 57576 65674 57588
rect 66993 57579 67051 57585
rect 66993 57576 67005 57579
rect 65668 57548 67005 57576
rect 65668 57536 65674 57548
rect 66993 57545 67005 57548
rect 67039 57545 67051 57579
rect 66993 57539 67051 57545
rect 67542 57536 67548 57588
rect 67600 57576 67606 57588
rect 67600 57548 74534 57576
rect 67600 57536 67606 57548
rect 13722 57468 13728 57520
rect 13780 57508 13786 57520
rect 63310 57508 63316 57520
rect 13780 57480 63316 57508
rect 13780 57468 13786 57480
rect 63310 57468 63316 57480
rect 63368 57468 63374 57520
rect 64138 57468 64144 57520
rect 64196 57468 64202 57520
rect 66809 57511 66867 57517
rect 66809 57508 66821 57511
rect 64248 57480 66821 57508
rect 15102 57400 15108 57452
rect 15160 57440 15166 57452
rect 63494 57440 63500 57452
rect 15160 57412 63500 57440
rect 15160 57400 15166 57412
rect 63494 57400 63500 57412
rect 63552 57400 63558 57452
rect 6822 57332 6828 57384
rect 6880 57372 6886 57384
rect 61562 57372 61568 57384
rect 6880 57344 61568 57372
rect 6880 57332 6886 57344
rect 61562 57332 61568 57344
rect 61620 57332 61626 57384
rect 62758 57332 62764 57384
rect 62816 57372 62822 57384
rect 64248 57372 64276 57480
rect 66809 57477 66821 57480
rect 66855 57477 66867 57511
rect 66809 57471 66867 57477
rect 66898 57468 66904 57520
rect 66956 57508 66962 57520
rect 69014 57508 69020 57520
rect 66956 57480 69020 57508
rect 66956 57468 66962 57480
rect 69014 57468 69020 57480
rect 69072 57468 69078 57520
rect 69109 57511 69167 57517
rect 69109 57477 69121 57511
rect 69155 57508 69167 57511
rect 72234 57508 72240 57520
rect 69155 57480 72240 57508
rect 69155 57477 69167 57480
rect 69109 57471 69167 57477
rect 72234 57468 72240 57480
rect 72292 57468 72298 57520
rect 74506 57508 74534 57548
rect 74718 57536 74724 57588
rect 74776 57576 74782 57588
rect 75638 57576 75644 57588
rect 74776 57548 75644 57576
rect 74776 57536 74782 57548
rect 75638 57536 75644 57548
rect 75696 57536 75702 57588
rect 77202 57536 77208 57588
rect 77260 57576 77266 57588
rect 79134 57576 79140 57588
rect 77260 57548 79140 57576
rect 77260 57536 77266 57548
rect 79134 57536 79140 57548
rect 79192 57536 79198 57588
rect 92566 57536 92572 57588
rect 92624 57576 92630 57588
rect 93670 57576 93676 57588
rect 92624 57548 93676 57576
rect 92624 57536 92630 57548
rect 93670 57536 93676 57548
rect 93728 57536 93734 57588
rect 94038 57536 94044 57588
rect 94096 57576 94102 57588
rect 94866 57576 94872 57588
rect 94096 57548 94872 57576
rect 94096 57536 94102 57548
rect 94866 57536 94872 57548
rect 94924 57536 94930 57588
rect 95234 57536 95240 57588
rect 95292 57576 95298 57588
rect 96522 57576 96528 57588
rect 95292 57548 96528 57576
rect 95292 57536 95298 57548
rect 96522 57536 96528 57548
rect 96580 57536 96586 57588
rect 96706 57536 96712 57588
rect 96764 57576 96770 57588
rect 97718 57576 97724 57588
rect 96764 57548 97724 57576
rect 96764 57536 96770 57548
rect 97718 57536 97724 57548
rect 97776 57536 97782 57588
rect 98178 57536 98184 57588
rect 98236 57576 98242 57588
rect 99098 57576 99104 57588
rect 98236 57548 99104 57576
rect 98236 57536 98242 57548
rect 99098 57536 99104 57548
rect 99156 57536 99162 57588
rect 100018 57536 100024 57588
rect 100076 57576 100082 57588
rect 100478 57576 100484 57588
rect 100076 57548 100484 57576
rect 100076 57536 100082 57548
rect 100478 57536 100484 57548
rect 100536 57536 100542 57588
rect 101766 57536 101772 57588
rect 101824 57576 101830 57588
rect 102042 57576 102048 57588
rect 101824 57548 102048 57576
rect 101824 57536 101830 57548
rect 102042 57536 102048 57548
rect 102100 57536 102106 57588
rect 102686 57536 102692 57588
rect 102744 57576 102750 57588
rect 103422 57576 103428 57588
rect 102744 57548 103428 57576
rect 102744 57536 102750 57548
rect 103422 57536 103428 57548
rect 103480 57536 103486 57588
rect 103882 57536 103888 57588
rect 103940 57576 103946 57588
rect 104710 57576 104716 57588
rect 103940 57548 104716 57576
rect 103940 57536 103946 57548
rect 104710 57536 104716 57548
rect 104768 57536 104774 57588
rect 105354 57536 105360 57588
rect 105412 57576 105418 57588
rect 106182 57576 106188 57588
rect 105412 57548 106188 57576
rect 105412 57536 105418 57548
rect 106182 57536 106188 57548
rect 106240 57536 106246 57588
rect 106550 57536 106556 57588
rect 106608 57576 106614 57588
rect 107470 57576 107476 57588
rect 106608 57548 107476 57576
rect 106608 57536 106614 57548
rect 107470 57536 107476 57548
rect 107528 57536 107534 57588
rect 109770 57536 109776 57588
rect 109828 57576 109834 57588
rect 110138 57576 110144 57588
rect 109828 57548 110144 57576
rect 109828 57536 109834 57548
rect 110138 57536 110144 57548
rect 110196 57536 110202 57588
rect 111886 57536 111892 57588
rect 111944 57576 111950 57588
rect 112990 57576 112996 57588
rect 111944 57548 112996 57576
rect 111944 57536 111950 57548
rect 112990 57536 112996 57548
rect 113048 57536 113054 57588
rect 113085 57579 113143 57585
rect 113085 57545 113097 57579
rect 113131 57576 113143 57579
rect 134444 57576 134472 57616
rect 135073 57613 135085 57616
rect 135119 57613 135131 57647
rect 135073 57607 135131 57613
rect 135254 57604 135260 57656
rect 135312 57644 135318 57656
rect 136361 57647 136419 57653
rect 136361 57644 136373 57647
rect 135312 57616 136373 57644
rect 135312 57604 135318 57616
rect 136361 57613 136373 57616
rect 136407 57613 136419 57647
rect 136361 57607 136419 57613
rect 113131 57548 134472 57576
rect 113131 57545 113143 57548
rect 113085 57539 113143 57545
rect 134518 57536 134524 57588
rect 134576 57576 134582 57588
rect 135162 57576 135168 57588
rect 134576 57548 135168 57576
rect 134576 57536 134582 57548
rect 135162 57536 135168 57548
rect 135220 57536 135226 57588
rect 135714 57536 135720 57588
rect 135772 57576 135778 57588
rect 136450 57576 136456 57588
rect 135772 57548 136456 57576
rect 135772 57536 135778 57548
rect 136450 57536 136456 57548
rect 136508 57536 136514 57588
rect 136560 57576 136588 57684
rect 136634 57672 136640 57724
rect 136692 57712 136698 57724
rect 137830 57712 137836 57724
rect 136692 57684 137836 57712
rect 136692 57672 136698 57684
rect 137830 57672 137836 57684
rect 137888 57672 137894 57724
rect 136729 57647 136787 57653
rect 136729 57613 136741 57647
rect 136775 57644 136787 57647
rect 138201 57647 138259 57653
rect 138201 57644 138213 57647
rect 136775 57616 138213 57644
rect 136775 57613 136787 57616
rect 136729 57607 136787 57613
rect 138201 57613 138213 57616
rect 138247 57613 138259 57647
rect 138201 57607 138259 57613
rect 138308 57576 138336 57752
rect 140314 57740 140320 57752
rect 140372 57740 140378 57792
rect 140498 57740 140504 57792
rect 140556 57780 140562 57792
rect 140556 57752 162256 57780
rect 140556 57740 140562 57752
rect 141329 57715 141387 57721
rect 141329 57681 141341 57715
rect 141375 57712 141387 57715
rect 141375 57684 143028 57712
rect 141375 57681 141387 57684
rect 141329 57675 141387 57681
rect 138385 57647 138443 57653
rect 138385 57613 138397 57647
rect 138431 57644 138443 57647
rect 143000 57644 143028 57684
rect 145834 57672 145840 57724
rect 145892 57712 145898 57724
rect 152553 57715 152611 57721
rect 152553 57712 152565 57715
rect 145892 57684 152565 57712
rect 145892 57672 145898 57684
rect 152553 57681 152565 57684
rect 152599 57681 152611 57715
rect 152553 57675 152611 57681
rect 152645 57715 152703 57721
rect 152645 57681 152657 57715
rect 152691 57712 152703 57715
rect 156877 57715 156935 57721
rect 156877 57712 156889 57715
rect 152691 57684 156889 57712
rect 152691 57681 152703 57684
rect 152645 57675 152703 57681
rect 156877 57681 156889 57684
rect 156923 57681 156935 57715
rect 162118 57712 162124 57724
rect 156877 57675 156935 57681
rect 157306 57684 162124 57712
rect 147214 57644 147220 57656
rect 138431 57616 142936 57644
rect 143000 57616 147220 57644
rect 138431 57613 138443 57616
rect 138385 57607 138443 57613
rect 142798 57576 142804 57588
rect 136560 57548 138014 57576
rect 138308 57548 142804 57576
rect 76742 57508 76748 57520
rect 74506 57480 76748 57508
rect 76742 57468 76748 57480
rect 76800 57468 76806 57520
rect 90174 57468 90180 57520
rect 90232 57508 90238 57520
rect 90910 57508 90916 57520
rect 90232 57480 90916 57508
rect 90232 57468 90238 57480
rect 90910 57468 90916 57480
rect 90968 57468 90974 57520
rect 95421 57511 95479 57517
rect 95421 57508 95433 57511
rect 93826 57480 95433 57508
rect 64414 57400 64420 57452
rect 64472 57440 64478 57452
rect 67818 57440 67824 57452
rect 64472 57412 67824 57440
rect 64472 57400 64478 57412
rect 67818 57400 67824 57412
rect 67876 57400 67882 57452
rect 67913 57443 67971 57449
rect 67913 57409 67925 57443
rect 67959 57440 67971 57443
rect 71038 57440 71044 57452
rect 67959 57412 71044 57440
rect 67959 57409 67971 57412
rect 67913 57403 67971 57409
rect 71038 57400 71044 57412
rect 71096 57400 71102 57452
rect 73062 57400 73068 57452
rect 73120 57440 73126 57452
rect 73120 57412 75132 57440
rect 73120 57400 73126 57412
rect 62816 57344 64276 57372
rect 62816 57332 62822 57344
rect 65518 57332 65524 57384
rect 65576 57372 65582 57384
rect 74994 57372 75000 57384
rect 65576 57344 75000 57372
rect 65576 57332 65582 57344
rect 74994 57332 75000 57344
rect 75052 57332 75058 57384
rect 75104 57372 75132 57412
rect 75178 57400 75184 57452
rect 75236 57440 75242 57452
rect 78490 57440 78496 57452
rect 75236 57412 78496 57440
rect 75236 57400 75242 57412
rect 78490 57400 78496 57412
rect 78548 57400 78554 57452
rect 88610 57400 88616 57452
rect 88668 57440 88674 57452
rect 93826 57440 93854 57480
rect 95421 57477 95433 57480
rect 95467 57477 95479 57511
rect 95421 57471 95479 57477
rect 95510 57468 95516 57520
rect 95568 57508 95574 57520
rect 96338 57508 96344 57520
rect 95568 57480 96344 57508
rect 95568 57468 95574 57480
rect 96338 57468 96344 57480
rect 96396 57468 96402 57520
rect 97258 57468 97264 57520
rect 97316 57508 97322 57520
rect 97316 57480 102272 57508
rect 97316 57468 97322 57480
rect 88668 57412 93854 57440
rect 88668 57400 88674 57412
rect 100846 57400 100852 57452
rect 100904 57440 100910 57452
rect 102042 57440 102048 57452
rect 100904 57412 102048 57440
rect 100904 57400 100910 57412
rect 102042 57400 102048 57412
rect 102100 57400 102106 57452
rect 102244 57440 102272 57480
rect 102318 57468 102324 57520
rect 102376 57508 102382 57520
rect 134889 57511 134947 57517
rect 134889 57508 134901 57511
rect 102376 57480 134901 57508
rect 102376 57468 102382 57480
rect 134889 57477 134901 57480
rect 134935 57477 134947 57511
rect 134889 57471 134947 57477
rect 135438 57468 135444 57520
rect 135496 57508 135502 57520
rect 136542 57508 136548 57520
rect 135496 57480 136548 57508
rect 135496 57468 135502 57480
rect 136542 57468 136548 57480
rect 136600 57468 136606 57520
rect 137986 57508 138014 57548
rect 142798 57536 142804 57548
rect 142856 57536 142862 57588
rect 142908 57576 142936 57616
rect 147214 57604 147220 57616
rect 147272 57604 147278 57656
rect 148594 57604 148600 57656
rect 148652 57644 148658 57656
rect 157153 57647 157211 57653
rect 157153 57644 157165 57647
rect 148652 57616 157165 57644
rect 148652 57604 148658 57616
rect 157153 57613 157165 57616
rect 157199 57613 157211 57647
rect 157153 57607 157211 57613
rect 143077 57579 143135 57585
rect 143077 57576 143089 57579
rect 142908 57548 143089 57576
rect 143077 57545 143089 57548
rect 143123 57545 143135 57579
rect 143077 57539 143135 57545
rect 152461 57579 152519 57585
rect 152461 57545 152473 57579
rect 152507 57576 152519 57579
rect 157306 57576 157334 57684
rect 162118 57672 162124 57684
rect 162176 57672 162182 57724
rect 162228 57712 162256 57752
rect 164602 57740 164608 57792
rect 164660 57780 164666 57792
rect 170769 57783 170827 57789
rect 170769 57780 170781 57783
rect 164660 57752 170781 57780
rect 164660 57740 164666 57752
rect 170769 57749 170781 57752
rect 170815 57749 170827 57783
rect 170769 57743 170827 57749
rect 170858 57740 170864 57792
rect 170916 57780 170922 57792
rect 214558 57780 214564 57792
rect 170916 57752 214564 57780
rect 170916 57740 170922 57752
rect 214558 57740 214564 57752
rect 214616 57740 214622 57792
rect 220630 57740 220636 57792
rect 220688 57780 220694 57792
rect 225690 57780 225696 57792
rect 220688 57752 225696 57780
rect 220688 57740 220694 57752
rect 225690 57740 225696 57752
rect 225748 57740 225754 57792
rect 166258 57712 166264 57724
rect 162228 57684 166264 57712
rect 166258 57672 166264 57684
rect 166316 57672 166322 57724
rect 166442 57672 166448 57724
rect 166500 57712 166506 57724
rect 213178 57712 213184 57724
rect 166500 57684 213184 57712
rect 166500 57672 166506 57684
rect 213178 57672 213184 57684
rect 213236 57672 213242 57724
rect 217410 57672 217416 57724
rect 217468 57712 217474 57724
rect 225230 57712 225236 57724
rect 217468 57684 225236 57712
rect 217468 57672 217474 57684
rect 225230 57672 225236 57684
rect 225288 57672 225294 57724
rect 157518 57604 157524 57656
rect 157576 57644 157582 57656
rect 162213 57647 162271 57653
rect 162213 57644 162225 57647
rect 157576 57616 162225 57644
rect 157576 57604 157582 57616
rect 162213 57613 162225 57616
rect 162259 57613 162271 57647
rect 162213 57607 162271 57613
rect 166994 57604 167000 57656
rect 167052 57644 167058 57656
rect 168190 57644 168196 57656
rect 167052 57616 168196 57644
rect 167052 57604 167058 57616
rect 168190 57604 168196 57616
rect 168248 57604 168254 57656
rect 168285 57647 168343 57653
rect 168285 57613 168297 57647
rect 168331 57644 168343 57647
rect 213270 57644 213276 57656
rect 168331 57616 213276 57644
rect 168331 57613 168343 57616
rect 168285 57607 168343 57613
rect 213270 57604 213276 57616
rect 213328 57604 213334 57656
rect 215294 57604 215300 57656
rect 215352 57644 215358 57656
rect 223117 57647 223175 57653
rect 223117 57644 223129 57647
rect 215352 57616 223129 57644
rect 215352 57604 215358 57616
rect 223117 57613 223129 57616
rect 223163 57613 223175 57647
rect 223117 57607 223175 57613
rect 152507 57548 157334 57576
rect 157981 57579 158039 57585
rect 152507 57545 152519 57548
rect 152461 57539 152519 57545
rect 157981 57545 157993 57579
rect 158027 57576 158039 57579
rect 158027 57548 166948 57576
rect 158027 57545 158039 57548
rect 157981 57539 158039 57545
rect 147030 57508 147036 57520
rect 137986 57480 147036 57508
rect 147030 57468 147036 57480
rect 147088 57468 147094 57520
rect 150342 57468 150348 57520
rect 150400 57508 150406 57520
rect 150400 57480 155632 57508
rect 150400 57468 150406 57480
rect 102873 57443 102931 57449
rect 102873 57440 102885 57443
rect 102244 57412 102885 57440
rect 102873 57409 102885 57412
rect 102919 57409 102931 57443
rect 102873 57403 102931 57409
rect 103238 57400 103244 57452
rect 103296 57440 103302 57452
rect 142614 57440 142620 57452
rect 103296 57412 142620 57440
rect 103296 57400 103302 57412
rect 142614 57400 142620 57412
rect 142672 57400 142678 57452
rect 143166 57400 143172 57452
rect 143224 57440 143230 57452
rect 152277 57443 152335 57449
rect 152277 57440 152289 57443
rect 143224 57412 152289 57440
rect 143224 57400 143230 57412
rect 152277 57409 152289 57412
rect 152323 57409 152335 57443
rect 152277 57403 152335 57409
rect 78214 57372 78220 57384
rect 75104 57344 78220 57372
rect 78214 57332 78220 57344
rect 78272 57332 78278 57384
rect 101398 57372 101404 57384
rect 89732 57344 101404 57372
rect 10962 57264 10968 57316
rect 11020 57304 11026 57316
rect 62390 57304 62396 57316
rect 11020 57276 62396 57304
rect 11020 57264 11026 57276
rect 62390 57264 62396 57276
rect 62448 57264 62454 57316
rect 63678 57264 63684 57316
rect 63736 57304 63742 57316
rect 64598 57304 64604 57316
rect 63736 57276 64604 57304
rect 63736 57264 63742 57276
rect 64598 57264 64604 57276
rect 64656 57264 64662 57316
rect 64877 57307 64935 57313
rect 64877 57273 64889 57307
rect 64923 57304 64935 57307
rect 66717 57307 66775 57313
rect 66717 57304 66729 57307
rect 64923 57276 66729 57304
rect 64923 57273 64935 57276
rect 64877 57267 64935 57273
rect 66717 57273 66729 57276
rect 66763 57273 66775 57307
rect 66717 57267 66775 57273
rect 66809 57307 66867 57313
rect 66809 57273 66821 57307
rect 66855 57304 66867 57307
rect 73154 57304 73160 57316
rect 66855 57276 73160 57304
rect 66855 57273 66867 57276
rect 66809 57267 66867 57273
rect 73154 57264 73160 57276
rect 73212 57264 73218 57316
rect 86862 57264 86868 57316
rect 86920 57304 86926 57316
rect 89732 57304 89760 57344
rect 101398 57332 101404 57344
rect 101456 57332 101462 57384
rect 103514 57332 103520 57384
rect 103572 57372 103578 57384
rect 104802 57372 104808 57384
rect 103572 57344 104808 57372
rect 103572 57332 103578 57344
rect 104802 57332 104808 57344
rect 104860 57332 104866 57384
rect 108574 57332 108580 57384
rect 108632 57372 108638 57384
rect 108942 57372 108948 57384
rect 108632 57344 108948 57372
rect 108632 57332 108638 57344
rect 108942 57332 108948 57344
rect 109000 57332 109006 57384
rect 109218 57332 109224 57384
rect 109276 57372 109282 57384
rect 110230 57372 110236 57384
rect 109276 57344 110236 57372
rect 109276 57332 109282 57344
rect 110230 57332 110236 57344
rect 110288 57332 110294 57384
rect 110690 57332 110696 57384
rect 110748 57372 110754 57384
rect 111426 57372 111432 57384
rect 110748 57344 111432 57372
rect 110748 57332 110754 57344
rect 111426 57332 111432 57344
rect 111484 57332 111490 57384
rect 111981 57375 112039 57381
rect 111981 57341 111993 57375
rect 112027 57372 112039 57375
rect 140133 57375 140191 57381
rect 140133 57372 140145 57375
rect 112027 57344 140145 57372
rect 112027 57341 112039 57344
rect 111981 57335 112039 57341
rect 140133 57341 140145 57344
rect 140179 57341 140191 57375
rect 144178 57372 144184 57384
rect 140133 57335 140191 57341
rect 143092 57344 144184 57372
rect 86920 57276 89760 57304
rect 86920 57264 86926 57276
rect 89806 57264 89812 57316
rect 89864 57304 89870 57316
rect 90726 57304 90732 57316
rect 89864 57276 90732 57304
rect 89864 57264 89870 57276
rect 90726 57264 90732 57276
rect 90784 57264 90790 57316
rect 98638 57304 98644 57316
rect 90836 57276 98644 57304
rect 4062 57196 4068 57248
rect 4120 57236 4126 57248
rect 60918 57236 60924 57248
rect 4120 57208 60924 57236
rect 4120 57196 4126 57208
rect 60918 57196 60924 57208
rect 60976 57196 60982 57248
rect 64230 57196 64236 57248
rect 64288 57236 64294 57248
rect 68833 57239 68891 57245
rect 64288 57208 68784 57236
rect 64288 57196 64294 57208
rect 33042 57128 33048 57180
rect 33100 57168 33106 57180
rect 68094 57168 68100 57180
rect 33100 57140 68100 57168
rect 33100 57128 33106 57140
rect 68094 57128 68100 57140
rect 68152 57128 68158 57180
rect 68756 57168 68784 57208
rect 68833 57205 68845 57239
rect 68879 57236 68891 57239
rect 70486 57236 70492 57248
rect 68879 57208 70492 57236
rect 68879 57205 68891 57208
rect 68833 57199 68891 57205
rect 70486 57196 70492 57208
rect 70544 57196 70550 57248
rect 71682 57196 71688 57248
rect 71740 57236 71746 57248
rect 77938 57236 77944 57248
rect 71740 57208 77944 57236
rect 71740 57196 71746 57208
rect 77938 57196 77944 57208
rect 77996 57196 78002 57248
rect 72602 57168 72608 57180
rect 68756 57140 72608 57168
rect 72602 57128 72608 57140
rect 72660 57128 72666 57180
rect 75822 57128 75828 57180
rect 75880 57168 75886 57180
rect 78858 57168 78864 57180
rect 75880 57140 78864 57168
rect 75880 57128 75886 57140
rect 78858 57128 78864 57140
rect 78916 57128 78922 57180
rect 85390 57128 85396 57180
rect 85448 57168 85454 57180
rect 90836 57168 90864 57276
rect 98638 57264 98644 57276
rect 98696 57264 98702 57316
rect 100662 57264 100668 57316
rect 100720 57304 100726 57316
rect 143092 57304 143120 57344
rect 144178 57332 144184 57344
rect 144236 57332 144242 57384
rect 145006 57332 145012 57384
rect 145064 57372 145070 57384
rect 152645 57375 152703 57381
rect 145064 57344 152504 57372
rect 145064 57332 145070 57344
rect 100720 57276 137324 57304
rect 100720 57264 100726 57276
rect 94222 57236 94228 57248
rect 85448 57140 90864 57168
rect 90928 57208 94228 57236
rect 85448 57128 85454 57140
rect 35802 57060 35808 57112
rect 35860 57100 35866 57112
rect 68646 57100 68652 57112
rect 35860 57072 68652 57100
rect 35860 57060 35866 57072
rect 68646 57060 68652 57072
rect 68704 57060 68710 57112
rect 68922 57060 68928 57112
rect 68980 57100 68986 57112
rect 77018 57100 77024 57112
rect 68980 57072 77024 57100
rect 68980 57060 68986 57072
rect 77018 57060 77024 57072
rect 77076 57060 77082 57112
rect 80238 57060 80244 57112
rect 80296 57100 80302 57112
rect 80422 57100 80428 57112
rect 80296 57072 80428 57100
rect 80296 57060 80302 57072
rect 80422 57060 80428 57072
rect 80480 57060 80486 57112
rect 83550 57060 83556 57112
rect 83608 57100 83614 57112
rect 90928 57100 90956 57208
rect 94222 57196 94228 57208
rect 94280 57196 94286 57248
rect 96614 57196 96620 57248
rect 96672 57236 96678 57248
rect 137189 57239 137247 57245
rect 137189 57236 137201 57239
rect 96672 57208 137201 57236
rect 96672 57196 96678 57208
rect 137189 57205 137201 57208
rect 137235 57205 137247 57239
rect 137296 57236 137324 57276
rect 137986 57276 143120 57304
rect 137986 57236 138014 57276
rect 144086 57264 144092 57316
rect 144144 57304 144150 57316
rect 152369 57307 152427 57313
rect 152369 57304 152381 57307
rect 144144 57276 152381 57304
rect 144144 57264 144150 57276
rect 152369 57273 152381 57276
rect 152415 57273 152427 57307
rect 152476 57304 152504 57344
rect 152645 57341 152657 57375
rect 152691 57372 152703 57375
rect 155494 57372 155500 57384
rect 152691 57344 155500 57372
rect 152691 57341 152703 57344
rect 152645 57335 152703 57341
rect 155494 57332 155500 57344
rect 155552 57332 155558 57384
rect 155604 57372 155632 57480
rect 156046 57468 156052 57520
rect 156104 57508 156110 57520
rect 157150 57508 157156 57520
rect 156104 57480 157156 57508
rect 156104 57468 156110 57480
rect 157150 57468 157156 57480
rect 157208 57468 157214 57520
rect 158809 57511 158867 57517
rect 158809 57477 158821 57511
rect 158855 57508 158867 57511
rect 166920 57508 166948 57548
rect 167362 57536 167368 57588
rect 167420 57576 167426 57588
rect 167420 57548 216076 57576
rect 167420 57536 167426 57548
rect 200945 57511 201003 57517
rect 200945 57508 200957 57511
rect 158855 57480 166856 57508
rect 166920 57480 200957 57508
rect 158855 57477 158867 57480
rect 158809 57471 158867 57477
rect 156874 57400 156880 57452
rect 156932 57440 156938 57452
rect 157242 57440 157248 57452
rect 156932 57412 157248 57440
rect 156932 57400 156938 57412
rect 157242 57400 157248 57412
rect 157300 57400 157306 57452
rect 158993 57443 159051 57449
rect 158993 57409 159005 57443
rect 159039 57440 159051 57443
rect 166721 57443 166779 57449
rect 166721 57440 166733 57443
rect 159039 57412 166733 57440
rect 159039 57409 159051 57412
rect 158993 57403 159051 57409
rect 166721 57409 166733 57412
rect 166767 57409 166779 57443
rect 166828 57440 166856 57480
rect 200945 57477 200957 57480
rect 200991 57477 201003 57511
rect 200945 57471 201003 57477
rect 201034 57468 201040 57520
rect 201092 57508 201098 57520
rect 201310 57508 201316 57520
rect 201092 57480 201316 57508
rect 201092 57468 201098 57480
rect 201310 57468 201316 57480
rect 201368 57468 201374 57520
rect 202506 57468 202512 57520
rect 202564 57508 202570 57520
rect 202782 57508 202788 57520
rect 202564 57480 202788 57508
rect 202564 57468 202570 57480
rect 202782 57468 202788 57480
rect 202840 57468 202846 57520
rect 203058 57468 203064 57520
rect 203116 57508 203122 57520
rect 203886 57508 203892 57520
rect 203116 57480 203892 57508
rect 203116 57468 203122 57480
rect 203886 57468 203892 57480
rect 203944 57468 203950 57520
rect 205174 57468 205180 57520
rect 205232 57508 205238 57520
rect 205450 57508 205456 57520
rect 205232 57480 205456 57508
rect 205232 57468 205238 57480
rect 205450 57468 205456 57480
rect 205508 57468 205514 57520
rect 205726 57468 205732 57520
rect 205784 57508 205790 57520
rect 206738 57508 206744 57520
rect 205784 57480 206744 57508
rect 205784 57468 205790 57480
rect 206738 57468 206744 57480
rect 206796 57468 206802 57520
rect 215938 57508 215944 57520
rect 209746 57480 215944 57508
rect 209746 57440 209774 57480
rect 215938 57468 215944 57480
rect 215996 57468 216002 57520
rect 166828 57412 209774 57440
rect 216048 57440 216076 57548
rect 218882 57536 218888 57588
rect 218940 57576 218946 57588
rect 227990 57576 227996 57588
rect 218940 57548 227996 57576
rect 218940 57536 218946 57548
rect 227990 57536 227996 57548
rect 228048 57536 228054 57588
rect 217962 57468 217968 57520
rect 218020 57508 218026 57520
rect 228542 57508 228548 57520
rect 218020 57480 228548 57508
rect 218020 57468 218026 57480
rect 228542 57468 228548 57480
rect 228600 57468 228606 57520
rect 220078 57440 220084 57452
rect 216048 57412 220084 57440
rect 166721 57403 166779 57409
rect 220078 57400 220084 57412
rect 220136 57400 220142 57452
rect 182453 57375 182511 57381
rect 182453 57372 182465 57375
rect 155604 57344 182465 57372
rect 182453 57341 182465 57344
rect 182499 57341 182511 57375
rect 182453 57335 182511 57341
rect 182542 57332 182548 57384
rect 182600 57372 182606 57384
rect 183278 57372 183284 57384
rect 182600 57344 183284 57372
rect 182600 57332 182606 57344
rect 183278 57332 183284 57344
rect 183336 57332 183342 57384
rect 184014 57332 184020 57384
rect 184072 57372 184078 57384
rect 184658 57372 184664 57384
rect 184072 57344 184664 57372
rect 184072 57332 184078 57344
rect 184658 57332 184664 57344
rect 184716 57332 184722 57384
rect 184934 57332 184940 57384
rect 184992 57372 184998 57384
rect 185854 57372 185860 57384
rect 184992 57344 185860 57372
rect 184992 57332 184998 57344
rect 185854 57332 185860 57344
rect 185912 57332 185918 57384
rect 186498 57332 186504 57384
rect 186556 57372 186562 57384
rect 187602 57372 187608 57384
rect 186556 57344 187608 57372
rect 186556 57332 186562 57344
rect 187602 57332 187608 57344
rect 187660 57332 187666 57384
rect 187786 57332 187792 57384
rect 187844 57372 187850 57384
rect 188522 57372 188528 57384
rect 187844 57344 188528 57372
rect 187844 57332 187850 57344
rect 188522 57332 188528 57344
rect 188580 57332 188586 57384
rect 189074 57332 189080 57384
rect 189132 57372 189138 57384
rect 190086 57372 190092 57384
rect 189132 57344 190092 57372
rect 189132 57332 189138 57344
rect 190086 57332 190092 57344
rect 190144 57332 190150 57384
rect 190546 57332 190552 57384
rect 190604 57372 190610 57384
rect 191558 57372 191564 57384
rect 190604 57344 191564 57372
rect 190604 57332 190610 57344
rect 191558 57332 191564 57344
rect 191616 57332 191622 57384
rect 192386 57332 192392 57384
rect 192444 57372 192450 57384
rect 193030 57372 193036 57384
rect 192444 57344 193036 57372
rect 192444 57332 192450 57344
rect 193030 57332 193036 57344
rect 193088 57332 193094 57384
rect 193214 57332 193220 57384
rect 193272 57372 193278 57384
rect 193674 57372 193680 57384
rect 193272 57344 193680 57372
rect 193272 57332 193278 57344
rect 193674 57332 193680 57344
rect 193732 57332 193738 57384
rect 195330 57332 195336 57384
rect 195388 57372 195394 57384
rect 195882 57372 195888 57384
rect 195388 57344 195888 57372
rect 195388 57332 195394 57344
rect 195882 57332 195888 57344
rect 195940 57332 195946 57384
rect 196526 57332 196532 57384
rect 196584 57372 196590 57384
rect 197078 57372 197084 57384
rect 196584 57344 197084 57372
rect 196584 57332 196590 57344
rect 197078 57332 197084 57344
rect 197136 57332 197142 57384
rect 197446 57332 197452 57384
rect 197504 57372 197510 57384
rect 198458 57372 198464 57384
rect 197504 57344 198464 57372
rect 197504 57332 197510 57344
rect 198458 57332 198464 57344
rect 198516 57332 198522 57384
rect 199194 57332 199200 57384
rect 199252 57372 199258 57384
rect 199838 57372 199844 57384
rect 199252 57344 199844 57372
rect 199252 57332 199258 57344
rect 199838 57332 199844 57344
rect 199896 57332 199902 57384
rect 200114 57332 200120 57384
rect 200172 57372 200178 57384
rect 201218 57372 201224 57384
rect 200172 57344 201224 57372
rect 200172 57332 200178 57344
rect 201218 57332 201224 57344
rect 201276 57332 201282 57384
rect 201586 57332 201592 57384
rect 201644 57372 201650 57384
rect 202782 57372 202788 57384
rect 201644 57344 202788 57372
rect 201644 57332 201650 57344
rect 202782 57332 202788 57344
rect 202840 57332 202846 57384
rect 203426 57332 203432 57384
rect 203484 57372 203490 57384
rect 204162 57372 204168 57384
rect 203484 57344 204168 57372
rect 203484 57332 203490 57344
rect 204162 57332 204168 57344
rect 204220 57332 204226 57384
rect 204254 57332 204260 57384
rect 204312 57372 204318 57384
rect 205542 57372 205548 57384
rect 204312 57344 205548 57372
rect 204312 57332 204318 57344
rect 205542 57332 205548 57344
rect 205600 57332 205606 57384
rect 206370 57332 206376 57384
rect 206428 57372 206434 57384
rect 391198 57372 391204 57384
rect 206428 57344 391204 57372
rect 206428 57332 206434 57344
rect 391198 57332 391204 57344
rect 391256 57332 391262 57384
rect 171137 57307 171195 57313
rect 171137 57304 171149 57307
rect 152476 57276 171149 57304
rect 152369 57267 152427 57273
rect 171137 57273 171149 57276
rect 171183 57273 171195 57307
rect 171137 57267 171195 57273
rect 171226 57264 171232 57316
rect 171284 57304 171290 57316
rect 172238 57304 172244 57316
rect 171284 57276 172244 57304
rect 171284 57264 171290 57276
rect 172238 57264 172244 57276
rect 172296 57264 172302 57316
rect 173986 57264 173992 57316
rect 174044 57304 174050 57316
rect 174906 57304 174912 57316
rect 174044 57276 174912 57304
rect 174044 57264 174050 57276
rect 174906 57264 174912 57276
rect 174964 57264 174970 57316
rect 175366 57264 175372 57316
rect 175424 57304 175430 57316
rect 176562 57304 176568 57316
rect 175424 57276 176568 57304
rect 175424 57264 175430 57276
rect 176562 57264 176568 57276
rect 176620 57264 176626 57316
rect 176838 57264 176844 57316
rect 176896 57304 176902 57316
rect 177666 57304 177672 57316
rect 176896 57276 177672 57304
rect 176896 57264 176902 57276
rect 177666 57264 177672 57276
rect 177724 57264 177730 57316
rect 178954 57264 178960 57316
rect 179012 57304 179018 57316
rect 179322 57304 179328 57316
rect 179012 57276 179328 57304
rect 179012 57264 179018 57276
rect 179322 57264 179328 57276
rect 179380 57264 179386 57316
rect 382918 57304 382924 57316
rect 180628 57276 382924 57304
rect 137296 57208 138014 57236
rect 138109 57239 138167 57245
rect 137189 57199 137247 57205
rect 138109 57205 138121 57239
rect 138155 57236 138167 57239
rect 142246 57236 142252 57248
rect 138155 57208 142252 57236
rect 138155 57205 138167 57208
rect 138109 57199 138167 57205
rect 142246 57196 142252 57208
rect 142304 57196 142310 57248
rect 142338 57196 142344 57248
rect 142396 57236 142402 57248
rect 152553 57239 152611 57245
rect 142396 57208 152504 57236
rect 142396 57196 142402 57208
rect 92198 57128 92204 57180
rect 92256 57168 92262 57180
rect 105538 57168 105544 57180
rect 92256 57140 105544 57168
rect 92256 57128 92262 57140
rect 105538 57128 105544 57140
rect 105596 57128 105602 57180
rect 107746 57128 107752 57180
rect 107804 57168 107810 57180
rect 108942 57168 108948 57180
rect 107804 57140 108948 57168
rect 107804 57128 107810 57140
rect 108942 57128 108948 57140
rect 109000 57128 109006 57180
rect 111334 57128 111340 57180
rect 111392 57168 111398 57180
rect 111702 57168 111708 57180
rect 111392 57140 111708 57168
rect 111392 57128 111398 57140
rect 111702 57128 111708 57140
rect 111760 57128 111766 57180
rect 113358 57128 113364 57180
rect 113416 57168 113422 57180
rect 114462 57168 114468 57180
rect 113416 57140 114468 57168
rect 113416 57128 113422 57140
rect 114462 57128 114468 57140
rect 114520 57128 114526 57180
rect 115474 57128 115480 57180
rect 115532 57168 115538 57180
rect 115750 57168 115756 57180
rect 115532 57140 115756 57168
rect 115532 57128 115538 57140
rect 115750 57128 115756 57140
rect 115808 57128 115814 57180
rect 116026 57128 116032 57180
rect 116084 57168 116090 57180
rect 116854 57168 116860 57180
rect 116084 57140 116860 57168
rect 116084 57128 116090 57140
rect 116854 57128 116860 57140
rect 116912 57128 116918 57180
rect 119246 57128 119252 57180
rect 119304 57168 119310 57180
rect 119614 57168 119620 57180
rect 119304 57140 119620 57168
rect 119304 57128 119310 57140
rect 119614 57128 119620 57140
rect 119672 57128 119678 57180
rect 121730 57128 121736 57180
rect 121788 57168 121794 57180
rect 122558 57168 122564 57180
rect 121788 57140 122564 57168
rect 121788 57128 121794 57140
rect 122558 57128 122564 57140
rect 122616 57128 122622 57180
rect 122653 57171 122711 57177
rect 122653 57137 122665 57171
rect 122699 57168 122711 57171
rect 124769 57171 124827 57177
rect 124769 57168 124781 57171
rect 122699 57140 124781 57168
rect 122699 57137 122711 57140
rect 122653 57131 122711 57137
rect 124769 57137 124781 57140
rect 124815 57137 124827 57171
rect 124769 57131 124827 57137
rect 124861 57171 124919 57177
rect 124861 57137 124873 57171
rect 124907 57168 124919 57171
rect 134058 57168 134064 57180
rect 124907 57140 134064 57168
rect 124907 57137 124919 57140
rect 124861 57131 124919 57137
rect 134058 57128 134064 57140
rect 134116 57128 134122 57180
rect 136910 57128 136916 57180
rect 136968 57168 136974 57180
rect 146389 57171 146447 57177
rect 146389 57168 146401 57171
rect 136968 57140 146401 57168
rect 136968 57128 136974 57140
rect 146389 57137 146401 57140
rect 146435 57137 146447 57171
rect 146389 57131 146447 57137
rect 149333 57171 149391 57177
rect 149333 57137 149345 57171
rect 149379 57168 149391 57171
rect 152369 57171 152427 57177
rect 152369 57168 152381 57171
rect 149379 57140 152381 57168
rect 149379 57137 149391 57140
rect 149333 57131 149391 57137
rect 152369 57137 152381 57140
rect 152415 57137 152427 57171
rect 152476 57168 152504 57208
rect 152553 57205 152565 57239
rect 152599 57236 152611 57239
rect 162121 57239 162179 57245
rect 162121 57236 162133 57239
rect 152599 57208 162133 57236
rect 152599 57205 152611 57208
rect 152553 57199 152611 57205
rect 162121 57205 162133 57208
rect 162167 57205 162179 57239
rect 162121 57199 162179 57205
rect 163774 57196 163780 57248
rect 163832 57236 163838 57248
rect 170585 57239 170643 57245
rect 170585 57236 170597 57239
rect 163832 57208 170597 57236
rect 163832 57196 163838 57208
rect 170585 57205 170597 57208
rect 170631 57205 170643 57239
rect 170585 57199 170643 57205
rect 171318 57196 171324 57248
rect 171376 57236 171382 57248
rect 172422 57236 172428 57248
rect 171376 57208 172428 57236
rect 171376 57196 171382 57208
rect 172422 57196 172428 57208
rect 172480 57196 172486 57248
rect 173894 57196 173900 57248
rect 173952 57236 173958 57248
rect 175090 57236 175096 57248
rect 173952 57208 175096 57236
rect 173952 57196 173958 57208
rect 175090 57196 175096 57208
rect 175148 57196 175154 57248
rect 177482 57196 177488 57248
rect 177540 57236 177546 57248
rect 177850 57236 177856 57248
rect 177540 57208 177856 57236
rect 177540 57196 177546 57208
rect 177850 57196 177856 57208
rect 177908 57196 177914 57248
rect 178310 57196 178316 57248
rect 178368 57236 178374 57248
rect 179230 57236 179236 57248
rect 178368 57208 179236 57236
rect 178368 57196 178374 57208
rect 179230 57196 179236 57208
rect 179288 57196 179294 57248
rect 179874 57196 179880 57248
rect 179932 57236 179938 57248
rect 180628 57236 180656 57276
rect 382918 57264 382924 57276
rect 382976 57264 382982 57316
rect 179932 57208 180656 57236
rect 179932 57196 179938 57208
rect 180702 57196 180708 57248
rect 180760 57236 180766 57248
rect 387058 57236 387064 57248
rect 180760 57208 387064 57236
rect 180760 57196 180766 57208
rect 387058 57196 387064 57208
rect 387116 57196 387122 57248
rect 158993 57171 159051 57177
rect 158993 57168 159005 57171
rect 152476 57140 159005 57168
rect 152369 57131 152427 57137
rect 158993 57137 159005 57140
rect 159039 57137 159051 57171
rect 173158 57168 173164 57180
rect 158993 57131 159051 57137
rect 159100 57140 159312 57168
rect 83608 57072 90956 57100
rect 83608 57060 83614 57072
rect 91370 57060 91376 57112
rect 91428 57100 91434 57112
rect 92382 57100 92388 57112
rect 91428 57072 92388 57100
rect 91428 57060 91434 57072
rect 92382 57060 92388 57072
rect 92440 57060 92446 57112
rect 98822 57060 98828 57112
rect 98880 57100 98886 57112
rect 99282 57100 99288 57112
rect 98880 57072 99288 57100
rect 98880 57060 98886 57072
rect 99282 57060 99288 57072
rect 99340 57060 99346 57112
rect 108022 57060 108028 57112
rect 108080 57100 108086 57112
rect 108666 57100 108672 57112
rect 108080 57072 108672 57100
rect 108080 57060 108086 57072
rect 108666 57060 108672 57072
rect 108724 57060 108730 57112
rect 110509 57103 110567 57109
rect 110509 57100 110521 57103
rect 110340 57072 110521 57100
rect 39942 56992 39948 57044
rect 40000 57032 40006 57044
rect 40000 57004 66944 57032
rect 40000 56992 40006 57004
rect 43438 56924 43444 56976
rect 43496 56964 43502 56976
rect 66916 56964 66944 57004
rect 66990 56992 66996 57044
rect 67048 57032 67054 57044
rect 76098 57032 76104 57044
rect 67048 57004 76104 57032
rect 67048 56992 67054 57004
rect 76098 56992 76104 57004
rect 76156 56992 76162 57044
rect 94590 56992 94596 57044
rect 94648 57032 94654 57044
rect 95050 57032 95056 57044
rect 94648 57004 95056 57032
rect 94648 56992 94654 57004
rect 95050 56992 95056 57004
rect 95108 56992 95114 57044
rect 95421 57035 95479 57041
rect 95421 57001 95433 57035
rect 95467 57032 95479 57035
rect 102870 57032 102876 57044
rect 95467 57004 102876 57032
rect 95467 57001 95479 57004
rect 95421 56995 95479 57001
rect 102870 56992 102876 57004
rect 102928 56992 102934 57044
rect 105078 56992 105084 57044
rect 105136 57032 105142 57044
rect 105136 57004 106780 57032
rect 105136 56992 105142 57004
rect 69842 56964 69848 56976
rect 43496 56936 66852 56964
rect 66916 56936 69848 56964
rect 43496 56924 43502 56936
rect 53742 56856 53748 56908
rect 53800 56896 53806 56908
rect 66717 56899 66775 56905
rect 66717 56896 66729 56899
rect 53800 56868 66729 56896
rect 53800 56856 53806 56868
rect 66717 56865 66729 56868
rect 66763 56865 66775 56899
rect 66824 56896 66852 56936
rect 69842 56924 69848 56936
rect 69900 56924 69906 56976
rect 73430 56964 73436 56976
rect 69952 56936 73436 56964
rect 68833 56899 68891 56905
rect 68833 56896 68845 56899
rect 66824 56868 68845 56896
rect 66717 56859 66775 56865
rect 68833 56865 68845 56868
rect 68879 56865 68891 56899
rect 68833 56859 68891 56865
rect 50338 56788 50344 56840
rect 50396 56828 50402 56840
rect 68465 56831 68523 56837
rect 50396 56800 68324 56828
rect 50396 56788 50402 56800
rect 62942 56720 62948 56772
rect 63000 56760 63006 56772
rect 64693 56763 64751 56769
rect 64693 56760 64705 56763
rect 63000 56732 64705 56760
rect 63000 56720 63006 56732
rect 64693 56729 64705 56732
rect 64739 56729 64751 56763
rect 64693 56723 64751 56729
rect 64782 56720 64788 56772
rect 64840 56760 64846 56772
rect 64877 56763 64935 56769
rect 64877 56760 64889 56763
rect 64840 56732 64889 56760
rect 64840 56720 64846 56732
rect 64877 56729 64889 56732
rect 64923 56729 64935 56763
rect 64877 56723 64935 56729
rect 64969 56763 65027 56769
rect 64969 56729 64981 56763
rect 65015 56760 65027 56763
rect 67913 56763 67971 56769
rect 67913 56760 67925 56763
rect 65015 56732 67925 56760
rect 65015 56729 65027 56732
rect 64969 56723 65027 56729
rect 67913 56729 67925 56732
rect 67959 56729 67971 56763
rect 67913 56723 67971 56729
rect 57238 56652 57244 56704
rect 57296 56692 57302 56704
rect 64233 56695 64291 56701
rect 64233 56692 64245 56695
rect 57296 56664 64245 56692
rect 57296 56652 57302 56664
rect 64233 56661 64245 56664
rect 64279 56661 64291 56695
rect 64233 56655 64291 56661
rect 64322 56652 64328 56704
rect 64380 56692 64386 56704
rect 68296 56692 68324 56800
rect 68465 56797 68477 56831
rect 68511 56828 68523 56831
rect 69952 56828 69980 56936
rect 73430 56924 73436 56936
rect 73488 56924 73494 56976
rect 82722 56924 82728 56976
rect 82780 56964 82786 56976
rect 87690 56964 87696 56976
rect 82780 56936 87696 56964
rect 82780 56924 82786 56936
rect 87690 56924 87696 56936
rect 87748 56924 87754 56976
rect 87782 56924 87788 56976
rect 87840 56964 87846 56976
rect 102778 56964 102784 56976
rect 87840 56936 102784 56964
rect 87840 56924 87846 56936
rect 102778 56924 102784 56936
rect 102836 56924 102842 56976
rect 105630 56924 105636 56976
rect 105688 56964 105694 56976
rect 106090 56964 106096 56976
rect 105688 56936 106096 56964
rect 105688 56924 105694 56936
rect 106090 56924 106096 56936
rect 106148 56924 106154 56976
rect 106752 56964 106780 57004
rect 106826 56992 106832 57044
rect 106884 57032 106890 57044
rect 110340 57032 110368 57072
rect 110509 57069 110521 57072
rect 110555 57069 110567 57103
rect 110509 57063 110567 57069
rect 114554 57060 114560 57112
rect 114612 57100 114618 57112
rect 115658 57100 115664 57112
rect 114612 57072 115664 57100
rect 114612 57060 114618 57072
rect 115658 57060 115664 57072
rect 115716 57060 115722 57112
rect 119062 57060 119068 57112
rect 119120 57100 119126 57112
rect 119890 57100 119896 57112
rect 119120 57072 119896 57100
rect 119120 57060 119126 57072
rect 119890 57060 119896 57072
rect 119948 57060 119954 57112
rect 120534 57060 120540 57112
rect 120592 57100 120598 57112
rect 133877 57103 133935 57109
rect 133877 57100 133889 57103
rect 120592 57072 133889 57100
rect 120592 57060 120598 57072
rect 133877 57069 133889 57072
rect 133923 57069 133935 57103
rect 133877 57063 133935 57069
rect 134889 57103 134947 57109
rect 134889 57069 134901 57103
rect 134935 57100 134947 57103
rect 137278 57100 137284 57112
rect 134935 57072 137284 57100
rect 134935 57069 134947 57072
rect 134889 57063 134947 57069
rect 137278 57060 137284 57072
rect 137336 57060 137342 57112
rect 137373 57103 137431 57109
rect 137373 57069 137385 57103
rect 137419 57100 137431 57103
rect 141326 57100 141332 57112
rect 137419 57072 141332 57100
rect 137419 57069 137431 57072
rect 137373 57063 137431 57069
rect 141326 57060 141332 57072
rect 141384 57060 141390 57112
rect 143074 57060 143080 57112
rect 143132 57100 143138 57112
rect 144362 57100 144368 57112
rect 143132 57072 144368 57100
rect 143132 57060 143138 57072
rect 144362 57060 144368 57072
rect 144420 57060 144426 57112
rect 146754 57060 146760 57112
rect 146812 57100 146818 57112
rect 159100 57100 159128 57140
rect 146812 57072 159128 57100
rect 146812 57060 146818 57072
rect 106884 57004 110368 57032
rect 106884 56992 106890 57004
rect 110414 56992 110420 57044
rect 110472 57032 110478 57044
rect 111702 57032 111708 57044
rect 110472 57004 111708 57032
rect 110472 56992 110478 57004
rect 111702 56992 111708 57004
rect 111760 56992 111766 57044
rect 116946 56992 116952 57044
rect 117004 57032 117010 57044
rect 117130 57032 117136 57044
rect 117004 57004 117136 57032
rect 117004 56992 117010 57004
rect 117130 56992 117136 57004
rect 117188 56992 117194 57044
rect 120258 56992 120264 57044
rect 120316 57032 120322 57044
rect 121270 57032 121276 57044
rect 120316 57004 121276 57032
rect 120316 56992 120322 57004
rect 121270 56992 121276 57004
rect 121328 56992 121334 57044
rect 121454 56992 121460 57044
rect 121512 57032 121518 57044
rect 142706 57032 142712 57044
rect 121512 57004 142712 57032
rect 121512 56992 121518 57004
rect 142706 56992 142712 57004
rect 142764 56992 142770 57044
rect 152090 56992 152096 57044
rect 152148 57032 152154 57044
rect 157061 57035 157119 57041
rect 157061 57032 157073 57035
rect 152148 57004 157073 57032
rect 152148 56992 152154 57004
rect 157061 57001 157073 57004
rect 157107 57001 157119 57035
rect 157061 56995 157119 57001
rect 157153 57035 157211 57041
rect 157153 57001 157165 57035
rect 157199 57032 157211 57035
rect 157199 57004 159220 57032
rect 157199 57001 157211 57004
rect 157153 56995 157211 57001
rect 113085 56967 113143 56973
rect 113085 56964 113097 56967
rect 106752 56936 113097 56964
rect 113085 56933 113097 56936
rect 113131 56933 113143 56967
rect 113085 56927 113143 56933
rect 117590 56924 117596 56976
rect 117648 56964 117654 56976
rect 133506 56964 133512 56976
rect 117648 56936 133512 56964
rect 117648 56924 117654 56936
rect 133506 56924 133512 56936
rect 133564 56924 133570 56976
rect 141329 56967 141387 56973
rect 141329 56964 141341 56967
rect 137296 56936 141341 56964
rect 84470 56856 84476 56908
rect 84528 56896 84534 56908
rect 88886 56896 88892 56908
rect 84528 56868 88892 56896
rect 84528 56856 84534 56868
rect 88886 56856 88892 56868
rect 88944 56856 88950 56908
rect 96982 56856 96988 56908
rect 97040 56896 97046 56908
rect 97902 56896 97908 56908
rect 97040 56868 97908 56896
rect 97040 56856 97046 56868
rect 97902 56856 97908 56868
rect 97960 56856 97966 56908
rect 104158 56856 104164 56908
rect 104216 56896 104222 56908
rect 111981 56899 112039 56905
rect 111981 56896 111993 56899
rect 104216 56868 111993 56896
rect 104216 56856 104222 56868
rect 111981 56865 111993 56868
rect 112027 56865 112039 56899
rect 111981 56859 112039 56865
rect 116394 56856 116400 56908
rect 116452 56896 116458 56908
rect 116946 56896 116952 56908
rect 116452 56868 116952 56896
rect 116452 56856 116458 56868
rect 116946 56856 116952 56868
rect 117004 56856 117010 56908
rect 118418 56856 118424 56908
rect 118476 56896 118482 56908
rect 124861 56899 124919 56905
rect 124861 56896 124873 56899
rect 118476 56868 124873 56896
rect 118476 56856 118482 56868
rect 124861 56865 124873 56868
rect 124907 56865 124919 56899
rect 124861 56859 124919 56865
rect 124953 56899 125011 56905
rect 124953 56865 124965 56899
rect 124999 56896 125011 56899
rect 128998 56896 129004 56908
rect 124999 56868 129004 56896
rect 124999 56865 125011 56868
rect 124953 56859 125011 56865
rect 128998 56856 129004 56868
rect 129056 56856 129062 56908
rect 130010 56856 130016 56908
rect 130068 56896 130074 56908
rect 137296 56896 137324 56936
rect 141329 56933 141341 56936
rect 141375 56933 141387 56967
rect 141329 56927 141387 56933
rect 141418 56924 141424 56976
rect 141476 56964 141482 56976
rect 150894 56964 150900 56976
rect 141476 56936 150900 56964
rect 141476 56924 141482 56936
rect 150894 56924 150900 56936
rect 150952 56924 150958 56976
rect 151262 56924 151268 56976
rect 151320 56964 151326 56976
rect 159085 56967 159143 56973
rect 159085 56964 159097 56967
rect 151320 56936 159097 56964
rect 151320 56924 151326 56936
rect 159085 56933 159097 56936
rect 159131 56933 159143 56967
rect 159085 56927 159143 56933
rect 130068 56868 137324 56896
rect 130068 56856 130074 56868
rect 137922 56856 137928 56908
rect 137980 56896 137986 56908
rect 143077 56899 143135 56905
rect 137980 56868 142476 56896
rect 137980 56856 137986 56868
rect 68511 56800 69980 56828
rect 68511 56797 68523 56800
rect 68465 56791 68523 56797
rect 70394 56788 70400 56840
rect 70452 56828 70458 56840
rect 74534 56828 74540 56840
rect 70452 56800 74540 56828
rect 70452 56788 70458 56800
rect 74534 56788 74540 56800
rect 74592 56788 74598 56840
rect 80882 56788 80888 56840
rect 80940 56828 80946 56840
rect 83182 56828 83188 56840
rect 80940 56800 83188 56828
rect 80940 56788 80946 56800
rect 83182 56788 83188 56800
rect 83240 56788 83246 56840
rect 84746 56788 84752 56840
rect 84804 56828 84810 56840
rect 87598 56828 87604 56840
rect 84804 56800 87604 56828
rect 84804 56788 84810 56800
rect 87598 56788 87604 56800
rect 87656 56788 87662 56840
rect 122006 56788 122012 56840
rect 122064 56828 122070 56840
rect 122742 56828 122748 56840
rect 122064 56800 122748 56828
rect 122064 56788 122070 56800
rect 122742 56788 122748 56800
rect 122800 56788 122806 56840
rect 123297 56831 123355 56837
rect 123297 56797 123309 56831
rect 123343 56828 123355 56831
rect 124677 56831 124735 56837
rect 124677 56828 124689 56831
rect 123343 56800 124689 56828
rect 123343 56797 123355 56800
rect 123297 56791 123355 56797
rect 124677 56797 124689 56800
rect 124723 56797 124735 56831
rect 124677 56791 124735 56797
rect 124769 56831 124827 56837
rect 124769 56797 124781 56831
rect 124815 56828 124827 56831
rect 129734 56828 129740 56840
rect 124815 56800 129740 56828
rect 124815 56797 124827 56800
rect 124769 56791 124827 56797
rect 129734 56788 129740 56800
rect 129792 56788 129798 56840
rect 132466 56800 133368 56828
rect 68370 56720 68376 56772
rect 68428 56760 68434 56772
rect 74902 56760 74908 56772
rect 68428 56732 74908 56760
rect 68428 56720 68434 56732
rect 74902 56720 74908 56732
rect 74960 56720 74966 56772
rect 82078 56720 82084 56772
rect 82136 56760 82142 56772
rect 83458 56760 83464 56772
rect 82136 56732 83464 56760
rect 82136 56720 82142 56732
rect 83458 56720 83464 56732
rect 83516 56720 83522 56772
rect 84194 56720 84200 56772
rect 84252 56760 84258 56772
rect 86218 56760 86224 56772
rect 84252 56732 86224 56760
rect 84252 56720 84258 56732
rect 86218 56720 86224 56732
rect 86276 56720 86282 56772
rect 114002 56720 114008 56772
rect 114060 56760 114066 56772
rect 122653 56763 122711 56769
rect 122653 56760 122665 56763
rect 114060 56732 122665 56760
rect 114060 56720 114066 56732
rect 122653 56729 122665 56732
rect 122699 56729 122711 56763
rect 122653 56723 122711 56729
rect 122926 56720 122932 56772
rect 122984 56760 122990 56772
rect 124030 56760 124036 56772
rect 122984 56732 124036 56760
rect 122984 56720 122990 56732
rect 124030 56720 124036 56732
rect 124088 56720 124094 56772
rect 124398 56720 124404 56772
rect 124456 56760 124462 56772
rect 125318 56760 125324 56772
rect 124456 56732 125324 56760
rect 124456 56720 124462 56732
rect 125318 56720 125324 56732
rect 125376 56720 125382 56772
rect 129182 56720 129188 56772
rect 129240 56760 129246 56772
rect 129642 56760 129648 56772
rect 129240 56732 129648 56760
rect 129240 56720 129246 56732
rect 129642 56720 129648 56732
rect 129700 56720 129706 56772
rect 71498 56692 71504 56704
rect 64380 56664 68140 56692
rect 68296 56664 71504 56692
rect 64380 56652 64386 56664
rect 62850 56584 62856 56636
rect 62908 56624 62914 56636
rect 64785 56627 64843 56633
rect 62908 56596 64736 56624
rect 62908 56584 62914 56596
rect 29638 56516 29644 56568
rect 29696 56556 29702 56568
rect 63034 56556 63040 56568
rect 29696 56528 63040 56556
rect 29696 56516 29702 56528
rect 63034 56516 63040 56528
rect 63092 56516 63098 56568
rect 64233 56559 64291 56565
rect 64233 56525 64245 56559
rect 64279 56556 64291 56559
rect 64598 56556 64604 56568
rect 64279 56528 64604 56556
rect 64279 56525 64291 56528
rect 64233 56519 64291 56525
rect 64598 56516 64604 56528
rect 64656 56516 64662 56568
rect 64708 56556 64736 56596
rect 64785 56593 64797 56627
rect 64831 56624 64843 56627
rect 65702 56624 65708 56636
rect 64831 56596 65708 56624
rect 64831 56593 64843 56596
rect 64785 56587 64843 56593
rect 65702 56584 65708 56596
rect 65760 56584 65766 56636
rect 65978 56584 65984 56636
rect 66036 56624 66042 56636
rect 67450 56624 67456 56636
rect 66036 56596 67456 56624
rect 66036 56584 66042 56596
rect 67450 56584 67456 56596
rect 67508 56584 67514 56636
rect 68112 56624 68140 56664
rect 71498 56652 71504 56664
rect 71556 56652 71562 56704
rect 81802 56652 81808 56704
rect 81860 56692 81866 56704
rect 82722 56692 82728 56704
rect 81860 56664 82728 56692
rect 81860 56652 81866 56664
rect 82722 56652 82728 56664
rect 82780 56652 82786 56704
rect 82998 56652 83004 56704
rect 83056 56692 83062 56704
rect 84010 56692 84016 56704
rect 83056 56664 84016 56692
rect 83056 56652 83062 56664
rect 84010 56652 84016 56664
rect 84068 56652 84074 56704
rect 85942 56652 85948 56704
rect 86000 56692 86006 56704
rect 86862 56692 86868 56704
rect 86000 56664 86868 56692
rect 86000 56652 86006 56664
rect 86862 56652 86868 56664
rect 86920 56652 86926 56704
rect 88334 56652 88340 56704
rect 88392 56692 88398 56704
rect 89438 56692 89444 56704
rect 88392 56664 89444 56692
rect 88392 56652 88398 56664
rect 89438 56652 89444 56664
rect 89496 56652 89502 56704
rect 123018 56652 123024 56704
rect 123076 56692 123082 56704
rect 124122 56692 124128 56704
rect 123076 56664 124128 56692
rect 123076 56652 123082 56664
rect 124122 56652 124128 56664
rect 124180 56652 124186 56704
rect 124214 56652 124220 56704
rect 124272 56692 124278 56704
rect 125042 56692 125048 56704
rect 124272 56664 125048 56692
rect 124272 56652 124278 56664
rect 125042 56652 125048 56664
rect 125100 56652 125106 56704
rect 70946 56624 70952 56636
rect 68112 56596 70952 56624
rect 70946 56584 70952 56596
rect 71004 56584 71010 56636
rect 71038 56584 71044 56636
rect 71096 56624 71102 56636
rect 75546 56624 75552 56636
rect 71096 56596 75552 56624
rect 71096 56584 71102 56596
rect 75546 56584 75552 56596
rect 75604 56584 75610 56636
rect 80606 56584 80612 56636
rect 80664 56624 80670 56636
rect 81250 56624 81256 56636
rect 80664 56596 81256 56624
rect 80664 56584 80670 56596
rect 81250 56584 81256 56596
rect 81308 56584 81314 56636
rect 81526 56584 81532 56636
rect 81584 56624 81590 56636
rect 82538 56624 82544 56636
rect 81584 56596 82544 56624
rect 81584 56584 81590 56596
rect 82538 56584 82544 56596
rect 82596 56584 82602 56636
rect 83274 56584 83280 56636
rect 83332 56624 83338 56636
rect 83918 56624 83924 56636
rect 83332 56596 83924 56624
rect 83332 56584 83338 56596
rect 83918 56584 83924 56596
rect 83976 56584 83982 56636
rect 85666 56584 85672 56636
rect 85724 56624 85730 56636
rect 86770 56624 86776 56636
rect 85724 56596 86776 56624
rect 85724 56584 85730 56596
rect 86770 56584 86776 56596
rect 86828 56584 86834 56636
rect 87506 56584 87512 56636
rect 87564 56624 87570 56636
rect 88242 56624 88248 56636
rect 87564 56596 88248 56624
rect 87564 56584 87570 56596
rect 88242 56584 88248 56596
rect 88300 56584 88306 56636
rect 88978 56584 88984 56636
rect 89036 56624 89042 56636
rect 89530 56624 89536 56636
rect 89036 56596 89536 56624
rect 89036 56584 89042 56596
rect 89530 56584 89536 56596
rect 89588 56584 89594 56636
rect 122837 56627 122895 56633
rect 122837 56593 122849 56627
rect 122883 56624 122895 56627
rect 132466 56624 132494 56800
rect 133340 56692 133368 56800
rect 133966 56788 133972 56840
rect 134024 56828 134030 56840
rect 135070 56828 135076 56840
rect 134024 56800 135076 56828
rect 134024 56788 134030 56800
rect 135070 56788 135076 56800
rect 135128 56788 135134 56840
rect 135165 56831 135223 56837
rect 135165 56797 135177 56831
rect 135211 56828 135223 56831
rect 140038 56828 140044 56840
rect 135211 56800 140044 56828
rect 135211 56797 135223 56800
rect 135165 56791 135223 56797
rect 140038 56788 140044 56800
rect 140096 56788 140102 56840
rect 142448 56828 142476 56868
rect 143077 56865 143089 56899
rect 143123 56896 143135 56899
rect 151906 56896 151912 56908
rect 143123 56868 151912 56896
rect 143123 56865 143135 56868
rect 143077 56859 143135 56865
rect 151906 56856 151912 56868
rect 151964 56856 151970 56908
rect 153930 56856 153936 56908
rect 153988 56896 153994 56908
rect 153988 56868 156552 56896
rect 153988 56856 153994 56868
rect 146938 56828 146944 56840
rect 142448 56800 146944 56828
rect 146938 56788 146944 56800
rect 146996 56788 147002 56840
rect 150526 56828 150532 56840
rect 147784 56800 150532 56828
rect 133877 56763 133935 56769
rect 133877 56729 133889 56763
rect 133923 56760 133935 56763
rect 138017 56763 138075 56769
rect 138017 56760 138029 56763
rect 133923 56732 138029 56760
rect 133923 56729 133935 56732
rect 133877 56723 133935 56729
rect 138017 56729 138029 56732
rect 138063 56729 138075 56763
rect 138017 56723 138075 56729
rect 138201 56763 138259 56769
rect 138201 56729 138213 56763
rect 138247 56760 138259 56763
rect 139670 56760 139676 56772
rect 138247 56732 139676 56760
rect 138247 56729 138259 56732
rect 138201 56723 138259 56729
rect 139670 56720 139676 56732
rect 139728 56720 139734 56772
rect 140133 56763 140191 56769
rect 140133 56729 140145 56763
rect 140179 56760 140191 56763
rect 146297 56763 146355 56769
rect 146297 56760 146309 56763
rect 140179 56732 146309 56760
rect 140179 56729 140191 56732
rect 140133 56723 140191 56729
rect 146297 56729 146309 56732
rect 146343 56729 146355 56763
rect 146297 56723 146355 56729
rect 146389 56763 146447 56769
rect 146389 56729 146401 56763
rect 146435 56760 146447 56763
rect 147674 56760 147680 56772
rect 146435 56732 147680 56760
rect 146435 56729 146447 56732
rect 146389 56723 146447 56729
rect 147674 56720 147680 56732
rect 147732 56720 147738 56772
rect 134242 56692 134248 56704
rect 133340 56664 134248 56692
rect 134242 56652 134248 56664
rect 134300 56652 134306 56704
rect 134426 56652 134432 56704
rect 134484 56692 134490 56704
rect 138109 56695 138167 56701
rect 138109 56692 138121 56695
rect 134484 56664 138121 56692
rect 134484 56652 134490 56664
rect 138109 56661 138121 56664
rect 138155 56661 138167 56695
rect 147784 56692 147812 56800
rect 150526 56788 150532 56800
rect 150584 56788 150590 56840
rect 153010 56788 153016 56840
rect 153068 56828 153074 56840
rect 155218 56828 155224 56840
rect 153068 56800 155224 56828
rect 153068 56788 153074 56800
rect 155218 56788 155224 56800
rect 155276 56788 155282 56840
rect 147858 56720 147864 56772
rect 147916 56760 147922 56772
rect 147916 56732 153240 56760
rect 147916 56720 147922 56732
rect 148318 56692 148324 56704
rect 138109 56655 138167 56661
rect 138308 56664 147812 56692
rect 147876 56664 148324 56692
rect 122883 56596 132494 56624
rect 122883 56593 122895 56596
rect 122837 56587 122895 56593
rect 133322 56584 133328 56636
rect 133380 56624 133386 56636
rect 133380 56596 136680 56624
rect 133380 56584 133386 56596
rect 64969 56559 65027 56565
rect 64969 56556 64981 56559
rect 64708 56528 64981 56556
rect 64969 56525 64981 56528
rect 65015 56525 65027 56559
rect 64969 56519 65027 56525
rect 66717 56559 66775 56565
rect 66717 56525 66729 56559
rect 66763 56556 66775 56559
rect 68465 56559 68523 56565
rect 68465 56556 68477 56559
rect 66763 56528 68477 56556
rect 66763 56525 66775 56528
rect 66717 56519 66775 56525
rect 68465 56525 68477 56528
rect 68511 56525 68523 56559
rect 136652 56556 136680 56596
rect 136726 56584 136732 56636
rect 136784 56624 136790 56636
rect 137922 56624 137928 56636
rect 136784 56596 137928 56624
rect 136784 56584 136790 56596
rect 137922 56584 137928 56596
rect 137980 56584 137986 56636
rect 138308 56624 138336 56664
rect 138032 56596 138336 56624
rect 138032 56556 138060 56596
rect 138382 56584 138388 56636
rect 138440 56624 138446 56636
rect 139118 56624 139124 56636
rect 138440 56596 139124 56624
rect 138440 56584 138446 56596
rect 139118 56584 139124 56596
rect 139176 56584 139182 56636
rect 139578 56584 139584 56636
rect 139636 56624 139642 56636
rect 140866 56624 140872 56636
rect 139636 56596 140872 56624
rect 139636 56584 139642 56596
rect 140866 56584 140872 56596
rect 140924 56584 140930 56636
rect 141142 56584 141148 56636
rect 141200 56624 141206 56636
rect 141970 56624 141976 56636
rect 141200 56596 141976 56624
rect 141200 56584 141206 56596
rect 141970 56584 141976 56596
rect 142028 56584 142034 56636
rect 143810 56584 143816 56636
rect 143868 56624 143874 56636
rect 144454 56624 144460 56636
rect 143868 56596 144460 56624
rect 143868 56584 143874 56596
rect 144454 56584 144460 56596
rect 144512 56584 144518 56636
rect 145282 56584 145288 56636
rect 145340 56624 145346 56636
rect 146202 56624 146208 56636
rect 145340 56596 146208 56624
rect 145340 56584 145346 56596
rect 146202 56584 146208 56596
rect 146260 56584 146266 56636
rect 146297 56627 146355 56633
rect 146297 56593 146309 56627
rect 146343 56624 146355 56627
rect 147876 56624 147904 56664
rect 148318 56652 148324 56664
rect 148376 56652 148382 56704
rect 151814 56652 151820 56704
rect 151872 56692 151878 56704
rect 153010 56692 153016 56704
rect 151872 56664 153016 56692
rect 151872 56652 151878 56664
rect 153010 56652 153016 56664
rect 153068 56652 153074 56704
rect 146343 56596 147904 56624
rect 146343 56593 146355 56596
rect 146297 56587 146355 56593
rect 147950 56584 147956 56636
rect 148008 56624 148014 56636
rect 148962 56624 148968 56636
rect 148008 56596 148968 56624
rect 148008 56584 148014 56596
rect 148962 56584 148968 56596
rect 149020 56584 149026 56636
rect 150618 56584 150624 56636
rect 150676 56624 150682 56636
rect 151722 56624 151728 56636
rect 150676 56596 151728 56624
rect 150676 56584 150682 56596
rect 151722 56584 151728 56596
rect 151780 56584 151786 56636
rect 152458 56584 152464 56636
rect 152516 56624 152522 56636
rect 153102 56624 153108 56636
rect 152516 56596 153108 56624
rect 152516 56584 152522 56596
rect 153102 56584 153108 56596
rect 153160 56584 153166 56636
rect 153212 56624 153240 56732
rect 153286 56720 153292 56772
rect 153344 56760 153350 56772
rect 156524 56760 156552 56868
rect 156598 56856 156604 56908
rect 156656 56896 156662 56908
rect 157702 56896 157708 56908
rect 156656 56868 157708 56896
rect 156656 56856 156662 56868
rect 157702 56856 157708 56868
rect 157760 56856 157766 56908
rect 159192 56896 159220 57004
rect 159284 56964 159312 57140
rect 166966 57140 173164 57168
rect 159361 57103 159419 57109
rect 159361 57069 159373 57103
rect 159407 57100 159419 57103
rect 166966 57100 166994 57140
rect 173158 57128 173164 57140
rect 173216 57128 173222 57180
rect 173618 57128 173624 57180
rect 173676 57168 173682 57180
rect 175918 57168 175924 57180
rect 173676 57140 175924 57168
rect 173676 57128 173682 57140
rect 175918 57128 175924 57140
rect 175976 57128 175982 57180
rect 176286 57128 176292 57180
rect 176344 57168 176350 57180
rect 176344 57140 177068 57168
rect 176344 57128 176350 57140
rect 159407 57072 166994 57100
rect 159407 57069 159419 57072
rect 159361 57063 159419 57069
rect 169110 57060 169116 57112
rect 169168 57100 169174 57112
rect 176565 57103 176623 57109
rect 176565 57100 176577 57103
rect 169168 57072 176577 57100
rect 169168 57060 169174 57072
rect 176565 57069 176577 57072
rect 176611 57069 176623 57103
rect 177040 57100 177068 57140
rect 177114 57128 177120 57180
rect 177172 57168 177178 57180
rect 177942 57168 177948 57180
rect 177172 57140 177948 57168
rect 177172 57128 177178 57140
rect 177942 57128 177948 57140
rect 178000 57128 178006 57180
rect 178037 57171 178095 57177
rect 178037 57137 178049 57171
rect 178083 57168 178095 57171
rect 216030 57168 216036 57180
rect 178083 57140 216036 57168
rect 178083 57137 178095 57140
rect 178037 57131 178095 57137
rect 216030 57128 216036 57140
rect 216088 57128 216094 57180
rect 223390 57128 223396 57180
rect 223448 57168 223454 57180
rect 233602 57168 233608 57180
rect 223448 57140 233608 57168
rect 223448 57128 223454 57140
rect 233602 57128 233608 57140
rect 233660 57128 233666 57180
rect 183925 57103 183983 57109
rect 183925 57100 183937 57103
rect 177040 57072 183937 57100
rect 176565 57063 176623 57069
rect 183925 57069 183937 57072
rect 183971 57069 183983 57103
rect 217318 57100 217324 57112
rect 183925 57063 183983 57069
rect 185596 57072 217324 57100
rect 162121 57035 162179 57041
rect 162121 57001 162133 57035
rect 162167 57032 162179 57035
rect 172514 57032 172520 57044
rect 162167 57004 172520 57032
rect 162167 57001 162179 57004
rect 162121 56995 162179 57001
rect 172514 56992 172520 57004
rect 172572 56992 172578 57044
rect 172698 56992 172704 57044
rect 172756 57032 172762 57044
rect 177945 57035 178003 57041
rect 177945 57032 177957 57035
rect 172756 57004 177957 57032
rect 172756 56992 172762 57004
rect 177945 57001 177957 57004
rect 177991 57001 178003 57035
rect 177945 56995 178003 57001
rect 178034 56992 178040 57044
rect 178092 57032 178098 57044
rect 185489 57035 185547 57041
rect 185489 57032 185501 57035
rect 178092 57004 185501 57032
rect 178092 56992 178098 57004
rect 185489 57001 185501 57004
rect 185535 57001 185547 57035
rect 185489 56995 185547 57001
rect 166905 56967 166963 56973
rect 166905 56964 166917 56967
rect 159284 56936 166917 56964
rect 166905 56933 166917 56936
rect 166951 56933 166963 56967
rect 166905 56927 166963 56933
rect 170030 56924 170036 56976
rect 170088 56964 170094 56976
rect 174538 56964 174544 56976
rect 170088 56936 174544 56964
rect 170088 56924 170094 56936
rect 174538 56924 174544 56936
rect 174596 56924 174602 56976
rect 174630 56924 174636 56976
rect 174688 56964 174694 56976
rect 185596 56964 185624 57072
rect 217318 57060 217324 57072
rect 217376 57060 217382 57112
rect 223117 57103 223175 57109
rect 223117 57069 223129 57103
rect 223163 57100 223175 57103
rect 230474 57100 230480 57112
rect 223163 57072 230480 57100
rect 223163 57069 223175 57072
rect 223117 57063 223175 57069
rect 230474 57060 230480 57072
rect 230532 57060 230538 57112
rect 185673 57035 185731 57041
rect 185673 57001 185685 57035
rect 185719 57032 185731 57035
rect 220170 57032 220176 57044
rect 185719 57004 220176 57032
rect 185719 57001 185731 57004
rect 185673 56995 185731 57001
rect 220170 56992 220176 57004
rect 220228 56992 220234 57044
rect 174688 56936 185624 56964
rect 174688 56924 174694 56936
rect 185762 56924 185768 56976
rect 185820 56964 185826 56976
rect 186130 56964 186136 56976
rect 185820 56936 186136 56964
rect 185820 56924 185826 56936
rect 186130 56924 186136 56936
rect 186188 56924 186194 56976
rect 186314 56924 186320 56976
rect 186372 56964 186378 56976
rect 186682 56964 186688 56976
rect 186372 56936 186688 56964
rect 186372 56924 186378 56936
rect 186682 56924 186688 56936
rect 186740 56924 186746 56976
rect 187878 56924 187884 56976
rect 187936 56964 187942 56976
rect 188890 56964 188896 56976
rect 187936 56936 188896 56964
rect 187936 56924 187942 56936
rect 188890 56924 188896 56936
rect 188948 56924 188954 56976
rect 210418 56964 210424 56976
rect 190426 56936 210424 56964
rect 162213 56899 162271 56905
rect 159192 56868 162072 56896
rect 158809 56763 158867 56769
rect 158809 56760 158821 56763
rect 153344 56732 154620 56760
rect 156524 56732 158821 56760
rect 153344 56720 153350 56732
rect 154206 56652 154212 56704
rect 154264 56692 154270 56704
rect 154482 56692 154488 56704
rect 154264 56664 154488 56692
rect 154264 56652 154270 56664
rect 154482 56652 154488 56664
rect 154540 56652 154546 56704
rect 154592 56624 154620 56732
rect 158809 56729 158821 56732
rect 158855 56729 158867 56763
rect 158809 56723 158867 56729
rect 158990 56720 158996 56772
rect 159048 56760 159054 56772
rect 159818 56760 159824 56772
rect 159048 56732 159824 56760
rect 159048 56720 159054 56732
rect 159818 56720 159824 56732
rect 159876 56720 159882 56772
rect 162044 56760 162072 56868
rect 162213 56865 162225 56899
rect 162259 56896 162271 56899
rect 162259 56868 181852 56896
rect 162259 56865 162271 56868
rect 162213 56859 162271 56865
rect 162121 56831 162179 56837
rect 162121 56797 162133 56831
rect 162167 56828 162179 56831
rect 169018 56828 169024 56840
rect 162167 56800 169024 56828
rect 162167 56797 162179 56800
rect 162121 56791 162179 56797
rect 169018 56788 169024 56800
rect 169076 56788 169082 56840
rect 171137 56831 171195 56837
rect 171137 56797 171149 56831
rect 171183 56828 171195 56831
rect 173250 56828 173256 56840
rect 171183 56800 173256 56828
rect 171183 56797 171195 56800
rect 171137 56791 171195 56797
rect 173250 56788 173256 56800
rect 173308 56788 173314 56840
rect 174814 56788 174820 56840
rect 174872 56828 174878 56840
rect 175182 56828 175188 56840
rect 174872 56800 175188 56828
rect 174872 56788 174878 56800
rect 175182 56788 175188 56800
rect 175240 56788 175246 56840
rect 180150 56788 180156 56840
rect 180208 56828 180214 56840
rect 180702 56828 180708 56840
rect 180208 56800 180708 56828
rect 180208 56788 180214 56800
rect 180702 56788 180708 56800
rect 180760 56788 180766 56840
rect 181824 56828 181852 56868
rect 182266 56856 182272 56908
rect 182324 56896 182330 56908
rect 183370 56896 183376 56908
rect 182324 56868 183376 56896
rect 182324 56856 182330 56868
rect 183370 56856 183376 56868
rect 183428 56856 183434 56908
rect 183925 56899 183983 56905
rect 183925 56865 183937 56899
rect 183971 56896 183983 56899
rect 190426 56896 190454 56936
rect 210418 56924 210424 56936
rect 210476 56924 210482 56976
rect 215018 56924 215024 56976
rect 215076 56964 215082 56976
rect 228726 56964 228732 56976
rect 215076 56936 228732 56964
rect 215076 56924 215082 56936
rect 228726 56924 228732 56936
rect 228784 56924 228790 56976
rect 183971 56868 190454 56896
rect 183971 56865 183983 56868
rect 183925 56859 183983 56865
rect 192110 56856 192116 56908
rect 192168 56896 192174 56908
rect 192938 56896 192944 56908
rect 192168 56868 192944 56896
rect 192168 56856 192174 56868
rect 192938 56856 192944 56868
rect 192996 56856 193002 56908
rect 193490 56856 193496 56908
rect 193548 56896 193554 56908
rect 194134 56896 194140 56908
rect 193548 56868 194140 56896
rect 193548 56856 193554 56868
rect 194134 56856 194140 56868
rect 194192 56856 194198 56908
rect 194778 56856 194784 56908
rect 194836 56896 194842 56908
rect 195698 56896 195704 56908
rect 194836 56868 195704 56896
rect 194836 56856 194842 56868
rect 195698 56856 195704 56868
rect 195756 56856 195762 56908
rect 196250 56856 196256 56908
rect 196308 56896 196314 56908
rect 196894 56896 196900 56908
rect 196308 56868 196900 56896
rect 196308 56856 196314 56868
rect 196894 56856 196900 56868
rect 196952 56856 196958 56908
rect 197630 56856 197636 56908
rect 197688 56896 197694 56908
rect 198642 56896 198648 56908
rect 197688 56868 198648 56896
rect 197688 56856 197694 56868
rect 198642 56856 198648 56868
rect 198700 56856 198706 56908
rect 198918 56856 198924 56908
rect 198976 56896 198982 56908
rect 199930 56896 199936 56908
rect 198976 56868 199936 56896
rect 198976 56856 198982 56868
rect 199930 56856 199936 56868
rect 199988 56856 199994 56908
rect 207014 56856 207020 56908
rect 207072 56896 207078 56908
rect 242158 56896 242164 56908
rect 207072 56868 242164 56896
rect 207072 56856 207078 56868
rect 242158 56856 242164 56868
rect 242216 56856 242222 56908
rect 184198 56828 184204 56840
rect 181824 56800 184204 56828
rect 184198 56788 184204 56800
rect 184256 56788 184262 56840
rect 189534 56788 189540 56840
rect 189592 56828 189598 56840
rect 190362 56828 190368 56840
rect 189592 56800 190368 56828
rect 189592 56788 189598 56800
rect 190362 56788 190368 56800
rect 190420 56788 190426 56840
rect 190822 56788 190828 56840
rect 190880 56828 190886 56840
rect 191374 56828 191380 56840
rect 190880 56800 191380 56828
rect 190880 56788 190886 56800
rect 191374 56788 191380 56800
rect 191432 56788 191438 56840
rect 193306 56788 193312 56840
rect 193364 56828 193370 56840
rect 194410 56828 194416 56840
rect 193364 56800 194416 56828
rect 193364 56788 193370 56800
rect 194410 56788 194416 56800
rect 194468 56788 194474 56840
rect 200945 56831 201003 56837
rect 200945 56797 200957 56831
rect 200991 56828 201003 56831
rect 209130 56828 209136 56840
rect 200991 56800 209136 56828
rect 200991 56797 201003 56800
rect 200945 56791 201003 56797
rect 209130 56788 209136 56800
rect 209188 56788 209194 56840
rect 210878 56788 210884 56840
rect 210936 56828 210942 56840
rect 233234 56828 233240 56840
rect 210936 56800 233240 56828
rect 210936 56788 210942 56800
rect 233234 56788 233240 56800
rect 233292 56788 233298 56840
rect 170490 56760 170496 56772
rect 162044 56732 170496 56760
rect 170490 56720 170496 56732
rect 170548 56720 170554 56772
rect 175642 56720 175648 56772
rect 175700 56760 175706 56772
rect 176470 56760 176476 56772
rect 175700 56732 176476 56760
rect 175700 56720 175706 56732
rect 176470 56720 176476 56732
rect 176528 56720 176534 56772
rect 176565 56763 176623 56769
rect 176565 56729 176577 56763
rect 176611 56760 176623 56763
rect 188338 56760 188344 56772
rect 176611 56732 188344 56760
rect 176611 56729 176623 56732
rect 176565 56723 176623 56729
rect 188338 56720 188344 56732
rect 188396 56720 188402 56772
rect 207566 56720 207572 56772
rect 207624 56760 207630 56772
rect 229554 56760 229560 56772
rect 207624 56732 229560 56760
rect 207624 56720 207630 56732
rect 229554 56720 229560 56732
rect 229612 56720 229618 56772
rect 157794 56652 157800 56704
rect 157852 56692 157858 56704
rect 158622 56692 158628 56704
rect 157852 56664 158628 56692
rect 157852 56652 157858 56664
rect 158622 56652 158628 56664
rect 158680 56652 158686 56704
rect 158898 56652 158904 56704
rect 158956 56692 158962 56704
rect 159634 56692 159640 56704
rect 158956 56664 159640 56692
rect 158956 56652 158962 56664
rect 159634 56652 159640 56664
rect 159692 56652 159698 56704
rect 160462 56652 160468 56704
rect 160520 56692 160526 56704
rect 161382 56692 161388 56704
rect 160520 56664 161388 56692
rect 160520 56652 160526 56664
rect 161382 56652 161388 56664
rect 161440 56652 161446 56704
rect 166350 56692 166356 56704
rect 164206 56664 166356 56692
rect 153212 56596 154436 56624
rect 136652 56528 138060 56556
rect 68465 56519 68523 56525
rect 34422 56448 34428 56500
rect 34480 56488 34486 56500
rect 68186 56488 68192 56500
rect 34480 56460 68192 56488
rect 34480 56448 34486 56460
rect 68186 56448 68192 56460
rect 68244 56448 68250 56500
rect 154408 56488 154436 56596
rect 154500 56596 154620 56624
rect 154500 56568 154528 56596
rect 156322 56584 156328 56636
rect 156380 56624 156386 56636
rect 156966 56624 156972 56636
rect 156380 56596 156972 56624
rect 156380 56584 156386 56596
rect 156966 56584 156972 56596
rect 157024 56584 157030 56636
rect 157061 56627 157119 56633
rect 157061 56593 157073 56627
rect 157107 56624 157119 56627
rect 157981 56627 158039 56633
rect 157981 56624 157993 56627
rect 157107 56596 157993 56624
rect 157107 56593 157119 56596
rect 157061 56587 157119 56593
rect 157981 56593 157993 56596
rect 158027 56593 158039 56627
rect 157981 56587 158039 56593
rect 158070 56584 158076 56636
rect 158128 56624 158134 56636
rect 158530 56624 158536 56636
rect 158128 56596 158536 56624
rect 158128 56584 158134 56596
rect 158530 56584 158536 56596
rect 158588 56584 158594 56636
rect 159542 56584 159548 56636
rect 159600 56624 159606 56636
rect 159910 56624 159916 56636
rect 159600 56596 159916 56624
rect 159600 56584 159606 56596
rect 159910 56584 159916 56596
rect 159968 56584 159974 56636
rect 160738 56584 160744 56636
rect 160796 56624 160802 56636
rect 161290 56624 161296 56636
rect 160796 56596 161296 56624
rect 160796 56584 160802 56596
rect 161290 56584 161296 56596
rect 161348 56584 161354 56636
rect 161658 56584 161664 56636
rect 161716 56624 161722 56636
rect 162578 56624 162584 56636
rect 161716 56596 162584 56624
rect 161716 56584 161722 56596
rect 162578 56584 162584 56596
rect 162636 56584 162642 56636
rect 162854 56584 162860 56636
rect 162912 56624 162918 56636
rect 164050 56624 164056 56636
rect 162912 56596 164056 56624
rect 162912 56584 162918 56596
rect 164050 56584 164056 56596
rect 164108 56584 164114 56636
rect 154482 56516 154488 56568
rect 154540 56516 154546 56568
rect 156877 56559 156935 56565
rect 156877 56525 156889 56559
rect 156923 56556 156935 56559
rect 164206 56556 164234 56664
rect 166350 56652 166356 56664
rect 166408 56652 166414 56704
rect 170398 56692 170404 56704
rect 167012 56664 170404 56692
rect 164326 56584 164332 56636
rect 164384 56624 164390 56636
rect 165154 56624 165160 56636
rect 164384 56596 165160 56624
rect 164384 56584 164390 56596
rect 165154 56584 165160 56596
rect 165212 56584 165218 56636
rect 165246 56584 165252 56636
rect 165304 56624 165310 56636
rect 165430 56624 165436 56636
rect 165304 56596 165436 56624
rect 165304 56584 165310 56596
rect 165430 56584 165436 56596
rect 165488 56584 165494 56636
rect 166166 56584 166172 56636
rect 166224 56624 166230 56636
rect 166902 56624 166908 56636
rect 166224 56596 166908 56624
rect 166224 56584 166230 56596
rect 166902 56584 166908 56596
rect 166960 56584 166966 56636
rect 156923 56528 164234 56556
rect 166721 56559 166779 56565
rect 156923 56525 156935 56528
rect 156877 56519 156935 56525
rect 166721 56525 166733 56559
rect 166767 56556 166779 56559
rect 167012 56556 167040 56664
rect 170398 56652 170404 56664
rect 170456 56652 170462 56704
rect 170585 56695 170643 56701
rect 170585 56661 170597 56695
rect 170631 56692 170643 56695
rect 170631 56664 172928 56692
rect 170631 56661 170643 56664
rect 170585 56655 170643 56661
rect 167089 56627 167147 56633
rect 167089 56593 167101 56627
rect 167135 56624 167147 56627
rect 169110 56624 169116 56636
rect 167135 56596 169116 56624
rect 167135 56593 167147 56596
rect 167089 56587 167147 56593
rect 169110 56584 169116 56596
rect 169168 56584 169174 56636
rect 172900 56624 172928 56664
rect 172974 56652 172980 56704
rect 173032 56692 173038 56704
rect 173802 56692 173808 56704
rect 173032 56664 173808 56692
rect 173032 56652 173038 56664
rect 173802 56652 173808 56664
rect 173860 56652 173866 56704
rect 179782 56652 179788 56704
rect 179840 56692 179846 56704
rect 180610 56692 180616 56704
rect 179840 56664 180616 56692
rect 179840 56652 179846 56664
rect 180610 56652 180616 56664
rect 180668 56652 180674 56704
rect 182453 56695 182511 56701
rect 182453 56661 182465 56695
rect 182499 56692 182511 56695
rect 186958 56692 186964 56704
rect 182499 56664 186964 56692
rect 182499 56661 182511 56664
rect 182453 56655 182511 56661
rect 186958 56652 186964 56664
rect 187016 56652 187022 56704
rect 201773 56695 201831 56701
rect 201773 56661 201785 56695
rect 201819 56692 201831 56695
rect 209038 56692 209044 56704
rect 201819 56664 209044 56692
rect 201819 56661 201831 56664
rect 201773 56655 201831 56661
rect 209038 56652 209044 56664
rect 209096 56652 209102 56704
rect 209958 56652 209964 56704
rect 210016 56692 210022 56704
rect 230566 56692 230572 56704
rect 210016 56664 230572 56692
rect 210016 56652 210022 56664
rect 230566 56652 230572 56664
rect 230624 56652 230630 56704
rect 179506 56624 179512 56636
rect 172900 56596 179512 56624
rect 179506 56584 179512 56596
rect 179564 56584 179570 56636
rect 185210 56584 185216 56636
rect 185268 56624 185274 56636
rect 185946 56624 185952 56636
rect 185268 56596 185952 56624
rect 185268 56584 185274 56596
rect 185946 56584 185952 56596
rect 186004 56584 186010 56636
rect 212902 56584 212908 56636
rect 212960 56624 212966 56636
rect 225046 56624 225052 56636
rect 212960 56596 225052 56624
rect 212960 56584 212966 56596
rect 225046 56584 225052 56596
rect 225104 56584 225110 56636
rect 166767 56528 167040 56556
rect 166767 56525 166779 56528
rect 166721 56519 166779 56525
rect 171502 56516 171508 56568
rect 171560 56556 171566 56568
rect 436738 56556 436744 56568
rect 171560 56528 436744 56556
rect 171560 56516 171566 56528
rect 436738 56516 436744 56528
rect 436796 56516 436802 56568
rect 162121 56491 162179 56497
rect 162121 56488 162133 56491
rect 154408 56460 162133 56488
rect 162121 56457 162133 56460
rect 162167 56457 162179 56491
rect 162121 56451 162179 56457
rect 181070 56448 181076 56500
rect 181128 56488 181134 56500
rect 454678 56488 454684 56500
rect 181128 56460 454684 56488
rect 181128 56448 181134 56460
rect 454678 56448 454684 56460
rect 454736 56448 454742 56500
rect 30282 56380 30288 56432
rect 30340 56420 30346 56432
rect 30340 56392 64874 56420
rect 30340 56380 30346 56392
rect 21358 56312 21364 56364
rect 21416 56352 21422 56364
rect 60366 56352 60372 56364
rect 21416 56324 60372 56352
rect 21416 56312 21422 56324
rect 60366 56312 60372 56324
rect 60424 56312 60430 56364
rect 64846 56352 64874 56392
rect 183738 56380 183744 56432
rect 183796 56420 183802 56432
rect 468478 56420 468484 56432
rect 183796 56392 468484 56420
rect 183796 56380 183802 56392
rect 468478 56380 468484 56392
rect 468536 56380 468542 56432
rect 65978 56352 65984 56364
rect 64846 56324 65984 56352
rect 65978 56312 65984 56324
rect 66036 56312 66042 56364
rect 182818 56312 182824 56364
rect 182876 56352 182882 56364
rect 461578 56352 461584 56364
rect 182876 56324 461584 56352
rect 182876 56312 182882 56324
rect 461578 56312 461584 56324
rect 461636 56312 461642 56364
rect 27522 56244 27528 56296
rect 27580 56284 27586 56296
rect 66070 56284 66076 56296
rect 27580 56256 66076 56284
rect 27580 56244 27586 56256
rect 66070 56244 66076 56256
rect 66128 56244 66134 56296
rect 184842 56244 184848 56296
rect 184900 56284 184906 56296
rect 472618 56284 472624 56296
rect 184900 56256 472624 56284
rect 184900 56244 184906 56256
rect 472618 56244 472624 56256
rect 472676 56244 472682 56296
rect 22830 56176 22836 56228
rect 22888 56216 22894 56228
rect 65426 56216 65432 56228
rect 22888 56188 65432 56216
rect 22888 56176 22894 56188
rect 65426 56176 65432 56188
rect 65484 56176 65490 56228
rect 185486 56176 185492 56228
rect 185544 56216 185550 56228
rect 475378 56216 475384 56228
rect 185544 56188 475384 56216
rect 185544 56176 185550 56188
rect 475378 56176 475384 56188
rect 475436 56176 475442 56228
rect 17862 56108 17868 56160
rect 17920 56148 17926 56160
rect 64046 56148 64052 56160
rect 17920 56120 64052 56148
rect 17920 56108 17926 56120
rect 64046 56108 64052 56120
rect 64104 56108 64110 56160
rect 187326 56108 187332 56160
rect 187384 56148 187390 56160
rect 479518 56148 479524 56160
rect 187384 56120 479524 56148
rect 187384 56108 187390 56120
rect 479518 56108 479524 56120
rect 479576 56108 479582 56160
rect 8202 56040 8208 56092
rect 8260 56080 8266 56092
rect 61838 56080 61844 56092
rect 8260 56052 61844 56080
rect 8260 56040 8266 56052
rect 61838 56040 61844 56052
rect 61896 56040 61902 56092
rect 182082 56040 182088 56092
rect 182140 56080 182146 56092
rect 483014 56080 483020 56092
rect 182140 56052 483020 56080
rect 182140 56040 182146 56052
rect 483014 56040 483020 56052
rect 483072 56040 483078 56092
rect 4798 55972 4804 56024
rect 4856 56012 4862 56024
rect 60642 56012 60648 56024
rect 4856 55984 60648 56012
rect 4856 55972 4862 55984
rect 60642 55972 60648 55984
rect 60700 55972 60706 56024
rect 93118 55972 93124 56024
rect 93176 56012 93182 56024
rect 112438 56012 112444 56024
rect 93176 55984 112444 56012
rect 93176 55972 93182 55984
rect 112438 55972 112444 55984
rect 112496 55972 112502 56024
rect 186590 55972 186596 56024
rect 186648 56012 186654 56024
rect 500954 56012 500960 56024
rect 186648 55984 500960 56012
rect 186648 55972 186654 55984
rect 500954 55972 500960 55984
rect 501012 55972 501018 56024
rect 56134 55904 56140 55956
rect 56192 55944 56198 55956
rect 580258 55944 580264 55956
rect 56192 55916 580264 55944
rect 56192 55904 56198 55916
rect 580258 55904 580264 55916
rect 580316 55904 580322 55956
rect 11698 55836 11704 55888
rect 11756 55876 11762 55888
rect 60090 55876 60096 55888
rect 11756 55848 60096 55876
rect 11756 55836 11762 55848
rect 60090 55836 60096 55848
rect 60148 55836 60154 55888
rect 99374 55836 99380 55888
rect 99432 55876 99438 55888
rect 152458 55876 152464 55888
rect 99432 55848 152464 55876
rect 99432 55836 99438 55848
rect 152458 55836 152464 55848
rect 152516 55836 152522 55888
rect 189350 55836 189356 55888
rect 189408 55876 189414 55888
rect 512638 55876 512644 55888
rect 189408 55848 512644 55876
rect 189408 55836 189414 55848
rect 512638 55836 512644 55848
rect 512696 55836 512702 55888
rect 41322 55768 41328 55820
rect 41380 55808 41386 55820
rect 69934 55808 69940 55820
rect 41380 55780 69940 55808
rect 41380 55768 41386 55780
rect 69934 55768 69940 55780
rect 69992 55768 69998 55820
rect 167638 55768 167644 55820
rect 167696 55808 167702 55820
rect 425698 55808 425704 55820
rect 167696 55780 425704 55808
rect 167696 55768 167702 55780
rect 425698 55768 425704 55780
rect 425756 55768 425762 55820
rect 48222 55700 48228 55752
rect 48280 55740 48286 55752
rect 71958 55740 71964 55752
rect 48280 55712 71964 55740
rect 48280 55700 48286 55712
rect 71958 55700 71964 55712
rect 72016 55700 72022 55752
rect 163130 55700 163136 55752
rect 163188 55740 163194 55752
rect 407758 55740 407764 55752
rect 163188 55712 407764 55740
rect 163188 55700 163194 55712
rect 407758 55700 407764 55712
rect 407816 55700 407822 55752
rect 52362 55632 52368 55684
rect 52420 55672 52426 55684
rect 72878 55672 72884 55684
rect 52420 55644 72884 55672
rect 52420 55632 52426 55644
rect 72878 55632 72884 55644
rect 72936 55632 72942 55684
rect 116670 55632 116676 55684
rect 116728 55672 116734 55684
rect 224954 55672 224960 55684
rect 116728 55644 224960 55672
rect 116728 55632 116734 55644
rect 224954 55632 224960 55644
rect 225012 55632 225018 55684
rect 55122 55564 55128 55616
rect 55180 55604 55186 55616
rect 73798 55604 73804 55616
rect 55180 55576 73804 55604
rect 55180 55564 55186 55576
rect 73798 55564 73804 55576
rect 73856 55564 73862 55616
rect 114922 55564 114928 55616
rect 114980 55604 114986 55616
rect 218054 55604 218060 55616
rect 114980 55576 218060 55604
rect 114980 55564 114986 55576
rect 218054 55564 218060 55576
rect 218112 55564 218118 55616
rect 59262 55496 59268 55548
rect 59320 55536 59326 55548
rect 70394 55536 70400 55548
rect 59320 55508 70400 55536
rect 59320 55496 59326 55508
rect 70394 55496 70400 55508
rect 70452 55496 70458 55548
rect 113082 55496 113088 55548
rect 113140 55536 113146 55548
rect 209774 55536 209780 55548
rect 113140 55508 209780 55536
rect 113140 55496 113146 55508
rect 209774 55496 209780 55508
rect 209832 55496 209838 55548
rect 133506 55428 133512 55480
rect 133564 55468 133570 55480
rect 227714 55468 227720 55480
rect 133564 55440 227720 55468
rect 133564 55428 133570 55440
rect 227714 55428 227720 55440
rect 227772 55428 227778 55480
rect 112162 55360 112168 55412
rect 112220 55400 112226 55412
rect 207014 55400 207020 55412
rect 112220 55372 207020 55400
rect 112220 55360 112226 55372
rect 207014 55360 207020 55372
rect 207072 55360 207078 55412
rect 129734 55292 129740 55344
rect 129792 55332 129798 55344
rect 213914 55332 213920 55344
rect 129792 55304 213920 55332
rect 129792 55292 129798 55304
rect 213914 55292 213920 55304
rect 213972 55292 213978 55344
rect 139946 55156 139952 55208
rect 140004 55196 140010 55208
rect 316034 55196 316040 55208
rect 140004 55168 316040 55196
rect 140004 55156 140010 55168
rect 316034 55156 316040 55168
rect 316092 55156 316098 55208
rect 140774 55088 140780 55140
rect 140832 55128 140838 55140
rect 320174 55128 320180 55140
rect 140832 55100 320180 55128
rect 140832 55088 140838 55100
rect 320174 55088 320180 55100
rect 320232 55088 320238 55140
rect 141694 55020 141700 55072
rect 141752 55060 141758 55072
rect 324314 55060 324320 55072
rect 141752 55032 324320 55060
rect 141752 55020 141758 55032
rect 324314 55020 324320 55032
rect 324372 55020 324378 55072
rect 142522 54952 142528 55004
rect 142580 54992 142586 55004
rect 327074 54992 327080 55004
rect 142580 54964 327080 54992
rect 142580 54952 142586 54964
rect 327074 54952 327080 54964
rect 327132 54952 327138 55004
rect 162302 54884 162308 54936
rect 162360 54924 162366 54936
rect 405734 54924 405740 54936
rect 162360 54896 405740 54924
rect 162360 54884 162366 54896
rect 405734 54884 405740 54896
rect 405792 54884 405798 54936
rect 164142 54816 164148 54868
rect 164200 54856 164206 54868
rect 412634 54856 412640 54868
rect 164200 54828 412640 54856
rect 164200 54816 164206 54828
rect 412634 54816 412640 54828
rect 412692 54816 412698 54868
rect 164970 54748 164976 54800
rect 165028 54788 165034 54800
rect 414658 54788 414664 54800
rect 165028 54760 414664 54788
rect 165028 54748 165034 54760
rect 414658 54748 414664 54760
rect 414716 54748 414722 54800
rect 167730 54680 167736 54732
rect 167788 54720 167794 54732
rect 427814 54720 427820 54732
rect 167788 54692 427820 54720
rect 167788 54680 167794 54692
rect 427814 54680 427820 54692
rect 427872 54680 427878 54732
rect 189534 54612 189540 54664
rect 189592 54652 189598 54664
rect 485038 54652 485044 54664
rect 189592 54624 485044 54652
rect 189592 54612 189598 54624
rect 485038 54612 485044 54624
rect 485096 54612 485102 54664
rect 187970 54544 187976 54596
rect 188028 54584 188034 54596
rect 507854 54584 507860 54596
rect 188028 54556 507860 54584
rect 188028 54544 188034 54556
rect 507854 54544 507860 54556
rect 507912 54544 507918 54596
rect 37182 54476 37188 54528
rect 37240 54516 37246 54528
rect 69198 54516 69204 54528
rect 37240 54488 69204 54516
rect 37240 54476 37246 54488
rect 69198 54476 69204 54488
rect 69256 54476 69262 54528
rect 193398 54476 193404 54528
rect 193456 54516 193462 54528
rect 530578 54516 530584 54528
rect 193456 54488 530584 54516
rect 193456 54476 193462 54488
rect 530578 54476 530584 54488
rect 530636 54476 530642 54528
rect 139026 54408 139032 54460
rect 139084 54448 139090 54460
rect 313274 54448 313280 54460
rect 139084 54420 313280 54448
rect 139084 54408 139090 54420
rect 313274 54408 313280 54420
rect 313332 54408 313338 54460
rect 140314 54340 140320 54392
rect 140372 54380 140378 54392
rect 309134 54380 309140 54392
rect 140372 54352 309140 54380
rect 140372 54340 140378 54352
rect 309134 54340 309140 54352
rect 309192 54340 309198 54392
rect 137186 54272 137192 54324
rect 137244 54312 137250 54324
rect 306374 54312 306380 54324
rect 137244 54284 306380 54312
rect 137244 54272 137250 54284
rect 306374 54272 306380 54284
rect 306432 54272 306438 54324
rect 136634 54204 136640 54256
rect 136692 54244 136698 54256
rect 302234 54244 302240 54256
rect 136692 54216 302240 54244
rect 136692 54204 136698 54216
rect 302234 54204 302240 54216
rect 302292 54204 302298 54256
rect 134058 54136 134064 54188
rect 134116 54176 134122 54188
rect 231854 54176 231860 54188
rect 134116 54148 231860 54176
rect 134116 54136 134122 54148
rect 231854 54136 231860 54148
rect 231912 54136 231918 54188
rect 155862 54068 155868 54120
rect 155920 54108 155926 54120
rect 222838 54108 222844 54120
rect 155920 54080 222844 54108
rect 155920 54068 155926 54080
rect 222838 54068 222844 54080
rect 222896 54068 222902 54120
rect 155494 53932 155500 53984
rect 155552 53972 155558 53984
rect 155862 53972 155868 53984
rect 155552 53944 155868 53972
rect 155552 53932 155558 53944
rect 155862 53932 155868 53944
rect 155920 53932 155926 53984
rect 149146 53728 149152 53780
rect 149204 53768 149210 53780
rect 353294 53768 353300 53780
rect 149204 53740 353300 53768
rect 149204 53728 149210 53740
rect 353294 53728 353300 53740
rect 353352 53728 353358 53780
rect 165798 53660 165804 53712
rect 165856 53700 165862 53712
rect 418798 53700 418804 53712
rect 165856 53672 418804 53700
rect 165856 53660 165862 53672
rect 418798 53660 418804 53672
rect 418856 53660 418862 53712
rect 166718 53592 166724 53644
rect 166776 53632 166782 53644
rect 421558 53632 421564 53644
rect 166776 53604 421564 53632
rect 166776 53592 166782 53604
rect 421558 53592 421564 53604
rect 421616 53592 421622 53644
rect 187786 53524 187792 53576
rect 187844 53564 187850 53576
rect 447778 53564 447784 53576
rect 187844 53536 447784 53564
rect 187844 53524 187850 53536
rect 447778 53524 447784 53536
rect 447836 53524 447842 53576
rect 168374 53456 168380 53508
rect 168432 53496 168438 53508
rect 430574 53496 430580 53508
rect 168432 53468 430580 53496
rect 168432 53456 168438 53468
rect 430574 53456 430580 53468
rect 430632 53456 430638 53508
rect 186498 53388 186504 53440
rect 186556 53428 186562 53440
rect 450538 53428 450544 53440
rect 186556 53400 450544 53428
rect 186556 53388 186562 53400
rect 450538 53388 450544 53400
rect 450596 53388 450602 53440
rect 171318 53320 171324 53372
rect 171376 53360 171382 53372
rect 445754 53360 445760 53372
rect 171376 53332 445760 53360
rect 171376 53320 171382 53332
rect 445754 53320 445760 53332
rect 445812 53320 445818 53372
rect 186314 53252 186320 53304
rect 186372 53292 186378 53304
rect 502334 53292 502340 53304
rect 186372 53264 502340 53292
rect 186372 53252 186378 53264
rect 502334 53252 502340 53264
rect 502392 53252 502398 53304
rect 191926 53184 191932 53236
rect 191984 53224 191990 53236
rect 519538 53224 519544 53236
rect 191984 53196 519544 53224
rect 191984 53184 191990 53196
rect 519538 53184 519544 53196
rect 519596 53184 519602 53236
rect 190914 53116 190920 53168
rect 190972 53156 190978 53168
rect 520274 53156 520280 53168
rect 190972 53128 520280 53156
rect 190972 53116 190978 53128
rect 520274 53116 520280 53128
rect 520332 53116 520338 53168
rect 192110 53048 192116 53100
rect 192168 53088 192174 53100
rect 526438 53088 526444 53100
rect 192168 53060 526444 53088
rect 192168 53048 192174 53060
rect 526438 53048 526444 53060
rect 526496 53048 526502 53100
rect 143442 52980 143448 53032
rect 143500 53020 143506 53032
rect 331214 53020 331220 53032
rect 143500 52992 331220 53020
rect 143500 52980 143506 52992
rect 331214 52980 331220 52992
rect 331272 52980 331278 53032
rect 124214 52912 124220 52964
rect 124272 52952 124278 52964
rect 258074 52952 258080 52964
rect 124272 52924 258080 52952
rect 124272 52912 124278 52924
rect 258074 52912 258080 52924
rect 258132 52912 258138 52964
rect 123202 52844 123208 52896
rect 123260 52884 123266 52896
rect 251174 52884 251180 52896
rect 123260 52856 251180 52884
rect 123260 52844 123266 52856
rect 251174 52844 251180 52856
rect 251232 52844 251238 52896
rect 118878 52776 118884 52828
rect 118936 52816 118942 52828
rect 233234 52816 233240 52828
rect 118936 52788 233240 52816
rect 118936 52776 118942 52788
rect 233234 52776 233240 52788
rect 233292 52776 233298 52828
rect 117682 52708 117688 52760
rect 117740 52748 117746 52760
rect 229094 52748 229100 52760
rect 117740 52720 229100 52748
rect 117740 52708 117746 52720
rect 229094 52708 229100 52720
rect 229152 52708 229158 52760
rect 144638 52368 144644 52420
rect 144696 52408 144702 52420
rect 335354 52408 335360 52420
rect 144696 52380 335360 52408
rect 144696 52368 144702 52380
rect 335354 52368 335360 52380
rect 335412 52368 335418 52420
rect 145558 52300 145564 52352
rect 145616 52340 145622 52352
rect 339494 52340 339500 52352
rect 145616 52312 339500 52340
rect 145616 52300 145622 52312
rect 339494 52300 339500 52312
rect 339552 52300 339558 52352
rect 146478 52232 146484 52284
rect 146536 52272 146542 52284
rect 342254 52272 342260 52284
rect 146536 52244 342260 52272
rect 146536 52232 146542 52244
rect 342254 52232 342260 52244
rect 342312 52232 342318 52284
rect 147398 52164 147404 52216
rect 147456 52204 147462 52216
rect 346394 52204 346400 52216
rect 147456 52176 346400 52204
rect 147456 52164 147462 52176
rect 346394 52164 346400 52176
rect 346452 52164 346458 52216
rect 148226 52096 148232 52148
rect 148284 52136 148290 52148
rect 349154 52136 349160 52148
rect 148284 52108 349160 52136
rect 148284 52096 148290 52108
rect 349154 52096 349160 52108
rect 349212 52096 349218 52148
rect 150066 52028 150072 52080
rect 150124 52068 150130 52080
rect 357434 52068 357440 52080
rect 150124 52040 357440 52068
rect 150124 52028 150130 52040
rect 357434 52028 357440 52040
rect 357492 52028 357498 52080
rect 168742 51960 168748 52012
rect 168800 52000 168806 52012
rect 431954 52000 431960 52012
rect 168800 51972 431960 52000
rect 168800 51960 168806 51972
rect 431954 51960 431960 51972
rect 432012 51960 432018 52012
rect 169938 51892 169944 51944
rect 169996 51932 170002 51944
rect 434714 51932 434720 51944
rect 169996 51904 434720 51932
rect 169996 51892 170002 51904
rect 434714 51892 434720 51904
rect 434772 51892 434778 51944
rect 174078 51824 174084 51876
rect 174136 51864 174142 51876
rect 452654 51864 452660 51876
rect 174136 51836 452660 51864
rect 174136 51824 174142 51836
rect 452654 51824 452660 51836
rect 452712 51824 452718 51876
rect 193674 51756 193680 51808
rect 193732 51796 193738 51808
rect 528554 51796 528560 51808
rect 193732 51768 528560 51796
rect 193732 51756 193738 51768
rect 528554 51756 528560 51768
rect 528612 51756 528618 51808
rect 97534 51688 97540 51740
rect 97592 51728 97598 51740
rect 142154 51728 142160 51740
rect 97592 51700 142160 51728
rect 97592 51688 97598 51700
rect 142154 51688 142160 51700
rect 142212 51688 142218 51740
rect 200390 51688 200396 51740
rect 200448 51728 200454 51740
rect 544378 51728 544384 51740
rect 200448 51700 544384 51728
rect 200448 51688 200454 51700
rect 544378 51688 544384 51700
rect 544436 51688 544442 51740
rect 144362 51620 144368 51672
rect 144420 51660 144426 51672
rect 328454 51660 328460 51672
rect 144420 51632 328460 51660
rect 144420 51620 144426 51632
rect 328454 51620 328460 51632
rect 328512 51620 328518 51672
rect 123018 51552 123024 51604
rect 123076 51592 123082 51604
rect 253934 51592 253940 51604
rect 123076 51564 253940 51592
rect 123076 51552 123082 51564
rect 253934 51552 253940 51564
rect 253992 51552 253998 51604
rect 119246 51484 119252 51536
rect 119304 51524 119310 51536
rect 235994 51524 236000 51536
rect 119304 51496 236000 51524
rect 119304 51484 119310 51496
rect 235994 51484 236000 51496
rect 236052 51484 236058 51536
rect 142246 51416 142252 51468
rect 142304 51456 142310 51468
rect 240134 51456 240140 51468
rect 142304 51428 240140 51456
rect 142304 51416 142310 51428
rect 240134 51416 240140 51428
rect 240192 51416 240198 51468
rect 159082 51008 159088 51060
rect 159140 51048 159146 51060
rect 393314 51048 393320 51060
rect 159140 51020 393320 51048
rect 159140 51008 159146 51020
rect 393314 51008 393320 51020
rect 393372 51008 393378 51060
rect 170306 50940 170312 50992
rect 170364 50980 170370 50992
rect 438854 50980 438860 50992
rect 170364 50952 438860 50980
rect 170364 50940 170370 50952
rect 438854 50940 438860 50952
rect 438912 50940 438918 50992
rect 173066 50872 173072 50924
rect 173124 50912 173130 50924
rect 443638 50912 443644 50924
rect 173124 50884 443644 50912
rect 173124 50872 173130 50884
rect 443638 50872 443644 50884
rect 443696 50872 443702 50924
rect 173986 50804 173992 50856
rect 174044 50844 174050 50856
rect 456886 50844 456892 50856
rect 174044 50816 456892 50844
rect 174044 50804 174050 50816
rect 456886 50804 456892 50816
rect 456944 50804 456950 50856
rect 193490 50736 193496 50788
rect 193548 50776 193554 50788
rect 489178 50776 489184 50788
rect 193548 50748 489184 50776
rect 193548 50736 193554 50748
rect 489178 50736 489184 50748
rect 489236 50736 489242 50788
rect 197630 50668 197636 50720
rect 197688 50708 197694 50720
rect 533338 50708 533344 50720
rect 197688 50680 533344 50708
rect 197688 50668 197694 50680
rect 533338 50668 533344 50680
rect 533396 50668 533402 50720
rect 199286 50600 199292 50652
rect 199344 50640 199350 50652
rect 537478 50640 537484 50652
rect 199344 50612 537484 50640
rect 199344 50600 199350 50612
rect 537478 50600 537484 50612
rect 537536 50600 537542 50652
rect 194870 50532 194876 50584
rect 194928 50572 194934 50584
rect 535454 50572 535460 50584
rect 194928 50544 535460 50572
rect 194928 50532 194934 50544
rect 535454 50532 535460 50544
rect 535512 50532 535518 50584
rect 196158 50464 196164 50516
rect 196216 50504 196222 50516
rect 539594 50504 539600 50516
rect 196216 50476 539600 50504
rect 196216 50464 196222 50476
rect 539594 50464 539600 50476
rect 539652 50464 539658 50516
rect 196618 50396 196624 50448
rect 196676 50436 196682 50448
rect 542354 50436 542360 50448
rect 196676 50408 542360 50436
rect 196676 50396 196682 50408
rect 542354 50396 542360 50408
rect 542412 50396 542418 50448
rect 197722 50328 197728 50380
rect 197780 50368 197786 50380
rect 546494 50368 546500 50380
rect 197780 50340 546500 50368
rect 197780 50328 197786 50340
rect 546494 50328 546500 50340
rect 546552 50328 546558 50380
rect 150894 50260 150900 50312
rect 150952 50300 150958 50312
rect 322934 50300 322940 50312
rect 150952 50272 322940 50300
rect 150952 50260 150958 50272
rect 322934 50260 322940 50272
rect 322992 50260 322998 50312
rect 137922 50192 137928 50244
rect 137980 50232 137986 50244
rect 284294 50232 284300 50244
rect 137980 50204 284300 50232
rect 137980 50192 137986 50204
rect 284294 50192 284300 50204
rect 284352 50192 284358 50244
rect 150618 49648 150624 49700
rect 150676 49688 150682 49700
rect 291194 49688 291200 49700
rect 150676 49660 291200 49688
rect 150676 49648 150682 49660
rect 291194 49648 291200 49660
rect 291252 49648 291258 49700
rect 151814 49580 151820 49632
rect 151872 49620 151878 49632
rect 298094 49620 298100 49632
rect 151872 49592 298100 49620
rect 151872 49580 151878 49592
rect 298094 49580 298100 49592
rect 298152 49580 298158 49632
rect 139670 49512 139676 49564
rect 139728 49552 139734 49564
rect 293954 49552 293960 49564
rect 139728 49524 293960 49552
rect 139728 49512 139734 49524
rect 293954 49512 293960 49524
rect 294012 49512 294018 49564
rect 155862 49444 155868 49496
rect 155920 49484 155926 49496
rect 311894 49484 311900 49496
rect 155920 49456 311900 49484
rect 155920 49444 155926 49456
rect 311894 49444 311900 49456
rect 311952 49444 311958 49496
rect 147950 49376 147956 49428
rect 148008 49416 148014 49428
rect 304994 49416 305000 49428
rect 148008 49388 305000 49416
rect 148008 49376 148014 49388
rect 304994 49376 305000 49388
rect 305052 49376 305058 49428
rect 172514 49308 172520 49360
rect 172572 49348 172578 49360
rect 340874 49348 340880 49360
rect 172572 49320 340880 49348
rect 172572 49308 172578 49320
rect 340874 49308 340880 49320
rect 340932 49308 340938 49360
rect 161566 49240 161572 49292
rect 161624 49280 161630 49292
rect 329834 49280 329840 49292
rect 161624 49252 329840 49280
rect 161624 49240 161630 49252
rect 329834 49240 329840 49252
rect 329892 49240 329898 49292
rect 140866 49172 140872 49224
rect 140924 49212 140930 49224
rect 316126 49212 316132 49224
rect 140924 49184 316132 49212
rect 140924 49172 140930 49184
rect 316126 49172 316132 49184
rect 316184 49172 316190 49224
rect 154850 49104 154856 49156
rect 154908 49144 154914 49156
rect 375374 49144 375380 49156
rect 154908 49116 375380 49144
rect 154908 49104 154914 49116
rect 375374 49104 375380 49116
rect 375432 49104 375438 49156
rect 157794 49036 157800 49088
rect 157852 49076 157858 49088
rect 382274 49076 382280 49088
rect 157852 49048 382280 49076
rect 157852 49036 157858 49048
rect 382274 49036 382280 49048
rect 382332 49036 382338 49088
rect 160370 48968 160376 49020
rect 160428 49008 160434 49020
rect 396718 49008 396724 49020
rect 160428 48980 396724 49008
rect 160428 48968 160434 48980
rect 396718 48968 396724 48980
rect 396776 48968 396782 49020
rect 147398 48900 147404 48952
rect 147456 48940 147462 48952
rect 276014 48940 276020 48952
rect 147456 48912 276020 48940
rect 147456 48900 147462 48912
rect 276014 48900 276020 48912
rect 276072 48900 276078 48952
rect 158438 47948 158444 48000
rect 158496 47988 158502 48000
rect 388438 47988 388444 48000
rect 158496 47960 388444 47988
rect 158496 47948 158502 47960
rect 388438 47948 388444 47960
rect 388496 47948 388502 48000
rect 179506 47880 179512 47932
rect 179564 47920 179570 47932
rect 411254 47920 411260 47932
rect 179564 47892 411260 47920
rect 179564 47880 179570 47892
rect 411254 47880 411260 47892
rect 411312 47880 411318 47932
rect 161106 47812 161112 47864
rect 161164 47852 161170 47864
rect 400214 47852 400220 47864
rect 161164 47824 400220 47852
rect 161164 47812 161170 47824
rect 400214 47812 400220 47824
rect 400272 47812 400278 47864
rect 164050 47744 164056 47796
rect 164108 47784 164114 47796
rect 407114 47784 407120 47796
rect 164108 47756 407120 47784
rect 164108 47744 164114 47756
rect 407114 47744 407120 47756
rect 407172 47744 407178 47796
rect 188338 47676 188344 47728
rect 188396 47716 188402 47728
rect 432046 47716 432052 47728
rect 188396 47688 432052 47716
rect 188396 47676 188402 47688
rect 432046 47676 432052 47688
rect 432104 47676 432110 47728
rect 210418 47608 210424 47660
rect 210476 47648 210482 47660
rect 460934 47648 460940 47660
rect 210476 47620 460940 47648
rect 210476 47608 210482 47620
rect 460934 47608 460940 47620
rect 460992 47608 460998 47660
rect 165338 47540 165344 47592
rect 165396 47580 165402 47592
rect 418154 47580 418160 47592
rect 165396 47552 418160 47580
rect 165396 47540 165402 47552
rect 418154 47540 418160 47552
rect 418212 47540 418218 47592
rect 287698 46860 287704 46912
rect 287756 46900 287762 46912
rect 580166 46900 580172 46912
rect 287756 46872 580172 46900
rect 287756 46860 287762 46872
rect 580166 46860 580172 46872
rect 580224 46860 580230 46912
rect 3510 45500 3516 45552
rect 3568 45540 3574 45552
rect 40678 45540 40684 45552
rect 3568 45512 40684 45540
rect 3568 45500 3574 45512
rect 40678 45500 40684 45512
rect 40736 45500 40742 45552
rect 3510 33056 3516 33108
rect 3568 33096 3574 33108
rect 22738 33096 22744 33108
rect 3568 33068 22744 33096
rect 3568 33056 3574 33068
rect 22738 33056 22744 33068
rect 22796 33056 22802 33108
rect 55766 33056 55772 33108
rect 55824 33096 55830 33108
rect 580166 33096 580172 33108
rect 55824 33068 580172 33096
rect 55824 33056 55830 33068
rect 580166 33056 580172 33068
rect 580224 33056 580230 33108
rect 216030 24148 216036 24200
rect 216088 24188 216094 24200
rect 447134 24188 447140 24200
rect 216088 24160 447140 24188
rect 216088 24148 216094 24160
rect 447134 24148 447140 24160
rect 447192 24148 447198 24200
rect 220170 24080 220176 24132
rect 220228 24120 220234 24132
rect 467834 24120 467840 24132
rect 220228 24092 467840 24120
rect 220228 24080 220234 24092
rect 467834 24080 467840 24092
rect 467892 24080 467898 24132
rect 86586 22720 86592 22772
rect 86644 22760 86650 22772
rect 103514 22760 103520 22772
rect 86644 22732 103520 22760
rect 86644 22720 86650 22732
rect 103514 22720 103520 22732
rect 103572 22720 103578 22772
rect 217318 22720 217324 22772
rect 217376 22760 217382 22772
rect 454034 22760 454040 22772
rect 217376 22732 454040 22760
rect 217376 22720 217382 22732
rect 454034 22720 454040 22732
rect 454092 22720 454098 22772
rect 214558 21360 214564 21412
rect 214616 21400 214622 21412
rect 440234 21400 440240 21412
rect 214616 21372 440240 21400
rect 214616 21360 214622 21372
rect 440234 21360 440240 21372
rect 440292 21360 440298 21412
rect 3510 20612 3516 20664
rect 3568 20652 3574 20664
rect 33778 20652 33784 20664
rect 3568 20624 33784 20652
rect 3568 20612 3574 20624
rect 33778 20612 33784 20624
rect 33836 20612 33842 20664
rect 55674 20612 55680 20664
rect 55732 20652 55738 20664
rect 580166 20652 580172 20664
rect 55732 20624 580172 20652
rect 55732 20612 55738 20624
rect 580166 20612 580172 20624
rect 580224 20612 580230 20664
rect 186958 20204 186964 20256
rect 187016 20244 187022 20256
rect 357526 20244 357532 20256
rect 187016 20216 357532 20244
rect 187016 20204 187022 20216
rect 357526 20204 357532 20216
rect 357584 20204 357590 20256
rect 213270 20136 213276 20188
rect 213328 20176 213334 20188
rect 404354 20176 404360 20188
rect 213328 20148 404360 20176
rect 213328 20136 213334 20148
rect 404354 20136 404360 20148
rect 404412 20136 404418 20188
rect 184198 20068 184204 20120
rect 184256 20108 184262 20120
rect 386414 20108 386420 20120
rect 184256 20080 386420 20108
rect 184256 20068 184262 20080
rect 386414 20068 386420 20080
rect 386472 20068 386478 20120
rect 220078 20000 220084 20052
rect 220136 20040 220142 20052
rect 425054 20040 425060 20052
rect 220136 20012 425060 20040
rect 220136 20000 220142 20012
rect 425054 20000 425060 20012
rect 425112 20000 425118 20052
rect 213178 19932 213184 19984
rect 213236 19972 213242 19984
rect 422294 19972 422300 19984
rect 213236 19944 422300 19972
rect 213236 19932 213242 19944
rect 422294 19932 422300 19944
rect 422352 19932 422358 19984
rect 147030 19252 147036 19304
rect 147088 19292 147094 19304
rect 287054 19292 287060 19304
rect 147088 19264 287060 19292
rect 147088 19252 147094 19264
rect 287054 19252 287060 19264
rect 287112 19252 287118 19304
rect 209130 19184 209136 19236
rect 209188 19224 209194 19236
rect 365714 19224 365720 19236
rect 209188 19196 365720 19224
rect 209188 19184 209194 19196
rect 365714 19184 365720 19196
rect 365772 19184 365778 19236
rect 173250 19116 173256 19168
rect 173308 19156 173314 19168
rect 336734 19156 336740 19168
rect 173308 19128 336740 19156
rect 173308 19116 173314 19128
rect 336734 19116 336740 19128
rect 336792 19116 336798 19168
rect 162118 19048 162124 19100
rect 162176 19088 162182 19100
rect 332594 19088 332600 19100
rect 162176 19060 332600 19088
rect 162176 19048 162182 19060
rect 332594 19048 332600 19060
rect 332652 19048 332658 19100
rect 169110 18980 169116 19032
rect 169168 19020 169174 19032
rect 343634 19020 343640 19032
rect 169168 18992 343640 19020
rect 169168 18980 169174 18992
rect 343634 18980 343640 18992
rect 343692 18980 343698 19032
rect 169018 18912 169024 18964
rect 169076 18952 169082 18964
rect 347774 18952 347780 18964
rect 169076 18924 347780 18952
rect 169076 18912 169082 18924
rect 347774 18912 347780 18924
rect 347832 18912 347838 18964
rect 170490 18844 170496 18896
rect 170548 18884 170554 18896
rect 350534 18884 350540 18896
rect 170548 18856 350540 18884
rect 170548 18844 170554 18856
rect 350534 18844 350540 18856
rect 350592 18844 350598 18896
rect 166350 18776 166356 18828
rect 166408 18816 166414 18828
rect 354674 18816 354680 18828
rect 166408 18788 354680 18816
rect 166408 18776 166414 18788
rect 354674 18776 354680 18788
rect 354732 18776 354738 18828
rect 173158 18708 173164 18760
rect 173216 18748 173222 18760
rect 361574 18748 361580 18760
rect 173216 18720 361580 18748
rect 173216 18708 173222 18720
rect 361574 18708 361580 18720
rect 361632 18708 361638 18760
rect 155218 18640 155224 18692
rect 155276 18680 155282 18692
rect 368474 18680 368480 18692
rect 155276 18652 368480 18680
rect 155276 18640 155282 18652
rect 368474 18640 368480 18652
rect 368532 18640 368538 18692
rect 88978 18572 88984 18624
rect 89036 18612 89042 18624
rect 96614 18612 96620 18624
rect 89036 18584 96620 18612
rect 89036 18572 89042 18584
rect 96614 18572 96620 18584
rect 96672 18572 96678 18624
rect 97626 18572 97632 18624
rect 97684 18612 97690 18624
rect 147122 18612 147128 18624
rect 97684 18584 147128 18612
rect 97684 18572 97690 18584
rect 147122 18572 147128 18584
rect 147180 18572 147186 18624
rect 161198 18572 161204 18624
rect 161256 18612 161262 18624
rect 401594 18612 401600 18624
rect 161256 18584 401600 18612
rect 161256 18572 161262 18584
rect 401594 18572 401600 18584
rect 401652 18572 401658 18624
rect 122466 18504 122472 18556
rect 122524 18544 122530 18556
rect 247034 18544 247040 18556
rect 122524 18516 247040 18544
rect 122524 18504 122530 18516
rect 247034 18504 247040 18516
rect 247092 18504 247098 18556
rect 115566 18436 115572 18488
rect 115624 18476 115630 18488
rect 220814 18476 220820 18488
rect 115624 18448 220820 18476
rect 115624 18436 115630 18448
rect 220814 18436 220820 18448
rect 220872 18436 220878 18488
rect 126514 17892 126520 17944
rect 126572 17932 126578 17944
rect 262214 17932 262220 17944
rect 126572 17904 262220 17932
rect 126572 17892 126578 17904
rect 262214 17892 262220 17904
rect 262272 17892 262278 17944
rect 127894 17824 127900 17876
rect 127952 17864 127958 17876
rect 266354 17864 266360 17876
rect 127952 17836 266360 17864
rect 127952 17824 127958 17836
rect 266354 17824 266360 17836
rect 266412 17824 266418 17876
rect 127986 17756 127992 17808
rect 128044 17796 128050 17808
rect 269114 17796 269120 17808
rect 128044 17768 269120 17796
rect 128044 17756 128050 17768
rect 269114 17756 269120 17768
rect 269172 17756 269178 17808
rect 129366 17688 129372 17740
rect 129424 17728 129430 17740
rect 273254 17728 273260 17740
rect 129424 17700 273260 17728
rect 129424 17688 129430 17700
rect 273254 17688 273260 17700
rect 273312 17688 273318 17740
rect 130746 17620 130752 17672
rect 130804 17660 130810 17672
rect 280154 17660 280160 17672
rect 130804 17632 280160 17660
rect 130804 17620 130810 17632
rect 280154 17620 280160 17632
rect 280212 17620 280218 17672
rect 166258 17552 166264 17604
rect 166316 17592 166322 17604
rect 318794 17592 318800 17604
rect 166316 17564 318800 17592
rect 166316 17552 166322 17564
rect 318794 17552 318800 17564
rect 318852 17552 318858 17604
rect 170398 17484 170404 17536
rect 170456 17524 170462 17536
rect 325694 17524 325700 17536
rect 170456 17496 325700 17524
rect 170456 17484 170462 17496
rect 325694 17484 325700 17496
rect 325752 17484 325758 17536
rect 142982 17416 142988 17468
rect 143040 17456 143046 17468
rect 300854 17456 300860 17468
rect 143040 17428 300860 17456
rect 143040 17416 143046 17428
rect 300854 17416 300860 17428
rect 300912 17416 300918 17468
rect 146938 17348 146944 17400
rect 146996 17388 147002 17400
rect 307754 17388 307760 17400
rect 146996 17360 307760 17388
rect 146996 17348 147002 17360
rect 307754 17348 307760 17360
rect 307812 17348 307818 17400
rect 97718 17280 97724 17332
rect 97776 17320 97782 17332
rect 119338 17320 119344 17332
rect 97776 17292 119344 17320
rect 97776 17280 97782 17292
rect 119338 17280 119344 17292
rect 119396 17280 119402 17332
rect 144730 17280 144736 17332
rect 144788 17320 144794 17332
rect 332686 17320 332692 17332
rect 144788 17292 332692 17320
rect 144788 17280 144794 17292
rect 332686 17280 332692 17292
rect 332744 17280 332750 17332
rect 94866 17212 94872 17264
rect 94924 17252 94930 17264
rect 122098 17252 122104 17264
rect 94924 17224 122104 17252
rect 94924 17212 94930 17224
rect 122098 17212 122104 17224
rect 122156 17212 122162 17264
rect 209038 17212 209044 17264
rect 209096 17252 209102 17264
rect 415486 17252 415492 17264
rect 209096 17224 415492 17252
rect 209096 17212 209102 17224
rect 415486 17212 415492 17224
rect 415544 17212 415550 17264
rect 125410 17144 125416 17196
rect 125468 17184 125474 17196
rect 259454 17184 259460 17196
rect 125468 17156 259460 17184
rect 125468 17144 125474 17156
rect 259454 17144 259460 17156
rect 259512 17144 259518 17196
rect 125318 17076 125324 17128
rect 125376 17116 125382 17128
rect 255314 17116 255320 17128
rect 125376 17088 255320 17116
rect 125376 17076 125382 17088
rect 255314 17076 255320 17088
rect 255372 17076 255378 17128
rect 142890 17008 142896 17060
rect 142948 17048 142954 17060
rect 242894 17048 242900 17060
rect 142948 17020 242900 17048
rect 142948 17008 142954 17020
rect 242894 17008 242900 17020
rect 242952 17008 242958 17060
rect 119798 16532 119804 16584
rect 119856 16572 119862 16584
rect 238110 16572 238116 16584
rect 119856 16544 238116 16572
rect 119856 16532 119862 16544
rect 238110 16532 238116 16544
rect 238168 16532 238174 16584
rect 121178 16464 121184 16516
rect 121236 16504 121242 16516
rect 241698 16504 241704 16516
rect 121236 16476 241704 16504
rect 121236 16464 121242 16476
rect 241698 16464 241704 16476
rect 241756 16464 241762 16516
rect 122558 16396 122564 16448
rect 122616 16436 122622 16448
rect 245194 16436 245200 16448
rect 122616 16408 245200 16436
rect 122616 16396 122622 16408
rect 245194 16396 245200 16408
rect 245252 16396 245258 16448
rect 122650 16328 122656 16380
rect 122708 16368 122714 16380
rect 248782 16368 248788 16380
rect 122708 16340 248788 16368
rect 122708 16328 122714 16340
rect 248782 16328 248788 16340
rect 248840 16328 248846 16380
rect 123938 16260 123944 16312
rect 123996 16300 124002 16312
rect 252370 16300 252376 16312
rect 123996 16272 252376 16300
rect 123996 16260 124002 16272
rect 252370 16260 252376 16272
rect 252428 16260 252434 16312
rect 201126 16192 201132 16244
rect 201184 16232 201190 16244
rect 560846 16232 560852 16244
rect 201184 16204 560852 16232
rect 201184 16192 201190 16204
rect 560846 16192 560852 16204
rect 560904 16192 560910 16244
rect 202414 16124 202420 16176
rect 202472 16164 202478 16176
rect 564434 16164 564440 16176
rect 202472 16136 564440 16164
rect 202472 16124 202478 16136
rect 564434 16124 564440 16136
rect 564492 16124 564498 16176
rect 203886 16056 203892 16108
rect 203944 16096 203950 16108
rect 568022 16096 568028 16108
rect 203944 16068 568028 16096
rect 203944 16056 203950 16068
rect 568022 16056 568028 16068
rect 568080 16056 568086 16108
rect 99006 15988 99012 16040
rect 99064 16028 99070 16040
rect 116578 16028 116584 16040
rect 99064 16000 116584 16028
rect 99064 15988 99070 16000
rect 116578 15988 116584 16000
rect 116636 15988 116642 16040
rect 203978 15988 203984 16040
rect 204036 16028 204042 16040
rect 571518 16028 571524 16040
rect 204036 16000 571524 16028
rect 204036 15988 204042 16000
rect 571518 15988 571524 16000
rect 571576 15988 571582 16040
rect 94958 15920 94964 15972
rect 95016 15960 95022 15972
rect 115198 15960 115204 15972
rect 95016 15932 115204 15960
rect 95016 15920 95022 15932
rect 115198 15920 115204 15932
rect 115256 15920 115262 15972
rect 205174 15920 205180 15972
rect 205232 15960 205238 15972
rect 575106 15960 575112 15972
rect 205232 15932 575112 15960
rect 205232 15920 205238 15932
rect 575106 15920 575112 15932
rect 575164 15920 575170 15972
rect 112990 15852 112996 15904
rect 113048 15892 113054 15904
rect 206186 15892 206192 15904
rect 113048 15864 206192 15892
rect 113048 15852 113054 15864
rect 206186 15852 206192 15864
rect 206244 15852 206250 15904
rect 206738 15852 206744 15904
rect 206796 15892 206802 15904
rect 578602 15892 578608 15904
rect 206796 15864 578608 15892
rect 206796 15852 206802 15864
rect 578602 15852 578608 15864
rect 578660 15852 578666 15904
rect 119890 15784 119896 15836
rect 119948 15824 119954 15836
rect 234614 15824 234620 15836
rect 119948 15796 234620 15824
rect 119948 15784 119954 15796
rect 234614 15784 234620 15796
rect 234672 15784 234678 15836
rect 118602 15716 118608 15768
rect 118660 15756 118666 15768
rect 231026 15756 231032 15768
rect 118660 15728 231032 15756
rect 118660 15716 118666 15728
rect 231026 15716 231032 15728
rect 231084 15716 231090 15768
rect 117038 15648 117044 15700
rect 117096 15688 117102 15700
rect 226334 15688 226340 15700
rect 117096 15660 226340 15688
rect 117096 15648 117102 15660
rect 226334 15648 226340 15660
rect 226392 15648 226398 15700
rect 116946 15580 116952 15632
rect 117004 15620 117010 15632
rect 223942 15620 223948 15632
rect 117004 15592 223948 15620
rect 117004 15580 117010 15592
rect 223942 15580 223948 15592
rect 224000 15580 224006 15632
rect 115750 15512 115756 15564
rect 115808 15552 115814 15564
rect 220446 15552 220452 15564
rect 115808 15524 220452 15552
rect 115808 15512 115814 15524
rect 220446 15512 220452 15524
rect 220504 15512 220510 15564
rect 115658 15444 115664 15496
rect 115716 15484 115722 15496
rect 216858 15484 216864 15496
rect 115716 15456 216864 15484
rect 115716 15444 115722 15456
rect 216858 15444 216864 15456
rect 216916 15444 216922 15496
rect 114278 15376 114284 15428
rect 114336 15416 114342 15428
rect 213362 15416 213368 15428
rect 114336 15388 213368 15416
rect 114336 15376 114342 15388
rect 213362 15376 213368 15388
rect 213420 15376 213426 15428
rect 112898 15308 112904 15360
rect 112956 15348 112962 15360
rect 209866 15348 209872 15360
rect 112956 15320 209872 15348
rect 112956 15308 112962 15320
rect 209866 15308 209872 15320
rect 209924 15308 209930 15360
rect 183186 15104 183192 15156
rect 183244 15144 183250 15156
rect 489914 15144 489920 15156
rect 183244 15116 489920 15144
rect 183244 15104 183250 15116
rect 489914 15104 489920 15116
rect 489972 15104 489978 15156
rect 184750 15036 184756 15088
rect 184808 15076 184814 15088
rect 493502 15076 493508 15088
rect 184808 15048 493508 15076
rect 184808 15036 184814 15048
rect 493502 15036 493508 15048
rect 493560 15036 493566 15088
rect 185946 14968 185952 15020
rect 186004 15008 186010 15020
rect 497090 15008 497096 15020
rect 186004 14980 497096 15008
rect 186004 14968 186010 14980
rect 497090 14968 497096 14980
rect 497148 14968 497154 15020
rect 186038 14900 186044 14952
rect 186096 14940 186102 14952
rect 500586 14940 500592 14952
rect 186096 14912 500592 14940
rect 186096 14900 186102 14912
rect 500586 14900 500592 14912
rect 500644 14900 500650 14952
rect 187326 14832 187332 14884
rect 187384 14872 187390 14884
rect 504174 14872 504180 14884
rect 187384 14844 504180 14872
rect 187384 14832 187390 14844
rect 504174 14832 504180 14844
rect 504232 14832 504238 14884
rect 188890 14764 188896 14816
rect 188948 14804 188954 14816
rect 507670 14804 507676 14816
rect 188948 14776 507676 14804
rect 188948 14764 188954 14776
rect 507670 14764 507676 14776
rect 507728 14764 507734 14816
rect 188706 14696 188712 14748
rect 188764 14736 188770 14748
rect 511258 14736 511264 14748
rect 188764 14708 511264 14736
rect 188764 14696 188770 14708
rect 511258 14696 511264 14708
rect 511316 14696 511322 14748
rect 190178 14628 190184 14680
rect 190236 14668 190242 14680
rect 514754 14668 514760 14680
rect 190236 14640 514760 14668
rect 190236 14628 190242 14640
rect 514754 14628 514760 14640
rect 514812 14628 514818 14680
rect 191558 14560 191564 14612
rect 191616 14600 191622 14612
rect 518342 14600 518348 14612
rect 191616 14572 518348 14600
rect 191616 14560 191622 14572
rect 518342 14560 518348 14572
rect 518400 14560 518406 14612
rect 191466 14492 191472 14544
rect 191524 14532 191530 14544
rect 521838 14532 521844 14544
rect 191524 14504 521844 14532
rect 191524 14492 191530 14504
rect 521838 14492 521844 14504
rect 521896 14492 521902 14544
rect 105998 14424 106004 14476
rect 106056 14464 106062 14476
rect 182542 14464 182548 14476
rect 106056 14436 182548 14464
rect 106056 14424 106062 14436
rect 182542 14424 182548 14436
rect 182600 14424 182606 14476
rect 193030 14424 193036 14476
rect 193088 14464 193094 14476
rect 525426 14464 525432 14476
rect 193088 14436 525432 14464
rect 193088 14424 193094 14436
rect 525426 14424 525432 14436
rect 525484 14424 525490 14476
rect 183278 14356 183284 14408
rect 183336 14396 183342 14408
rect 486418 14396 486424 14408
rect 183336 14368 486424 14396
rect 183336 14356 183342 14368
rect 486418 14356 486424 14368
rect 486476 14356 486482 14408
rect 181990 14288 181996 14340
rect 182048 14328 182054 14340
rect 481634 14328 481640 14340
rect 182048 14300 481640 14328
rect 182048 14288 182054 14300
rect 481634 14288 481640 14300
rect 481692 14288 481698 14340
rect 180518 14220 180524 14272
rect 180576 14260 180582 14272
rect 478138 14260 478144 14272
rect 180576 14232 478144 14260
rect 180576 14220 180582 14232
rect 478138 14220 478144 14232
rect 478196 14220 478202 14272
rect 180610 14152 180616 14204
rect 180668 14192 180674 14204
rect 473354 14192 473360 14204
rect 180668 14164 473360 14192
rect 180668 14152 180674 14164
rect 473354 14152 473360 14164
rect 473412 14152 473418 14204
rect 179046 14084 179052 14136
rect 179104 14124 179110 14136
rect 471054 14124 471060 14136
rect 179104 14096 471060 14124
rect 179104 14084 179110 14096
rect 471054 14084 471060 14096
rect 471112 14084 471118 14136
rect 177758 14016 177764 14068
rect 177816 14056 177822 14068
rect 467466 14056 467472 14068
rect 177816 14028 467472 14056
rect 177816 14016 177822 14028
rect 467466 14016 467472 14028
rect 467524 14016 467530 14068
rect 177666 13948 177672 14000
rect 177724 13988 177730 14000
rect 463970 13988 463976 14000
rect 177724 13960 463976 13988
rect 177724 13948 177730 13960
rect 463970 13948 463976 13960
rect 464028 13948 464034 14000
rect 176286 13880 176292 13932
rect 176344 13920 176350 13932
rect 460382 13920 460388 13932
rect 176344 13892 460388 13920
rect 176344 13880 176350 13892
rect 460382 13880 460388 13892
rect 460440 13880 460446 13932
rect 158530 13744 158536 13796
rect 158588 13784 158594 13796
rect 389450 13784 389456 13796
rect 158588 13756 389456 13784
rect 158588 13744 158594 13756
rect 389450 13744 389456 13756
rect 389508 13744 389514 13796
rect 159818 13676 159824 13728
rect 159876 13716 159882 13728
rect 393038 13716 393044 13728
rect 159876 13688 393044 13716
rect 159876 13676 159882 13688
rect 393038 13676 393044 13688
rect 393096 13676 393102 13728
rect 159726 13608 159732 13660
rect 159784 13648 159790 13660
rect 396534 13648 396540 13660
rect 159784 13620 396540 13648
rect 159784 13608 159790 13620
rect 396534 13608 396540 13620
rect 396592 13608 396598 13660
rect 161290 13540 161296 13592
rect 161348 13580 161354 13592
rect 398834 13580 398840 13592
rect 161348 13552 398840 13580
rect 161348 13540 161354 13552
rect 398834 13540 398840 13552
rect 398892 13540 398898 13592
rect 162578 13472 162584 13524
rect 162636 13512 162642 13524
rect 403618 13512 403624 13524
rect 162636 13484 403624 13512
rect 162636 13472 162642 13484
rect 403618 13472 403624 13484
rect 403676 13472 403682 13524
rect 162670 13404 162676 13456
rect 162728 13444 162734 13456
rect 407206 13444 407212 13456
rect 162728 13416 407212 13444
rect 162728 13404 162734 13416
rect 407206 13404 407212 13416
rect 407264 13404 407270 13456
rect 163958 13336 163964 13388
rect 164016 13376 164022 13388
rect 410794 13376 410800 13388
rect 164016 13348 410800 13376
rect 164016 13336 164022 13348
rect 410794 13336 410800 13348
rect 410852 13336 410858 13388
rect 165246 13268 165252 13320
rect 165304 13308 165310 13320
rect 414290 13308 414296 13320
rect 165304 13280 414296 13308
rect 165304 13268 165310 13280
rect 414290 13268 414296 13280
rect 414348 13268 414354 13320
rect 165430 13200 165436 13252
rect 165488 13240 165494 13252
rect 417878 13240 417884 13252
rect 165488 13212 417884 13240
rect 165488 13200 165494 13212
rect 417878 13200 417884 13212
rect 417936 13200 417942 13252
rect 166902 13132 166908 13184
rect 166960 13172 166966 13184
rect 421374 13172 421380 13184
rect 166960 13144 421380 13172
rect 166960 13132 166966 13144
rect 421374 13132 421380 13144
rect 421432 13132 421438 13184
rect 168190 13064 168196 13116
rect 168248 13104 168254 13116
rect 423766 13104 423772 13116
rect 168248 13076 423772 13104
rect 168248 13064 168254 13076
rect 423766 13064 423772 13076
rect 423824 13064 423830 13116
rect 157058 12996 157064 13048
rect 157116 13036 157122 13048
rect 385954 13036 385960 13048
rect 157116 13008 385960 13036
rect 157116 12996 157122 13008
rect 385954 12996 385960 13008
rect 386012 12996 386018 13048
rect 156966 12928 156972 12980
rect 157024 12968 157030 12980
rect 382366 12968 382372 12980
rect 157024 12940 382372 12968
rect 157024 12928 157030 12940
rect 382366 12928 382372 12940
rect 382424 12928 382430 12980
rect 155770 12860 155776 12912
rect 155828 12900 155834 12912
rect 378870 12900 378876 12912
rect 155828 12872 378876 12900
rect 155828 12860 155834 12872
rect 378870 12860 378876 12872
rect 378928 12860 378934 12912
rect 154206 12792 154212 12844
rect 154264 12832 154270 12844
rect 373994 12832 374000 12844
rect 154264 12804 374000 12832
rect 154264 12792 154270 12804
rect 373994 12792 374000 12804
rect 374052 12792 374058 12844
rect 154298 12724 154304 12776
rect 154356 12764 154362 12776
rect 371694 12764 371700 12776
rect 154356 12736 371700 12764
rect 154356 12724 154362 12736
rect 371694 12724 371700 12736
rect 371752 12724 371758 12776
rect 152918 12656 152924 12708
rect 152976 12696 152982 12708
rect 368198 12696 368204 12708
rect 152976 12668 368204 12696
rect 152976 12656 152982 12668
rect 368198 12656 368204 12668
rect 368256 12656 368262 12708
rect 153010 12588 153016 12640
rect 153068 12628 153074 12640
rect 364610 12628 364616 12640
rect 153068 12600 364616 12628
rect 153068 12588 153074 12600
rect 364610 12588 364616 12600
rect 364668 12588 364674 12640
rect 151538 12520 151544 12572
rect 151596 12560 151602 12572
rect 361114 12560 361120 12572
rect 151596 12532 361120 12560
rect 151596 12520 151602 12532
rect 361114 12520 361120 12532
rect 361172 12520 361178 12572
rect 133598 12384 133604 12436
rect 133656 12424 133662 12436
rect 290182 12424 290188 12436
rect 133656 12396 290188 12424
rect 133656 12384 133662 12396
rect 290182 12384 290188 12396
rect 290240 12384 290246 12436
rect 135070 12316 135076 12368
rect 135128 12356 135134 12368
rect 293678 12356 293684 12368
rect 135128 12328 293684 12356
rect 135128 12316 135134 12328
rect 293678 12316 293684 12328
rect 293736 12316 293742 12368
rect 134978 12248 134984 12300
rect 135036 12288 135042 12300
rect 297266 12288 297272 12300
rect 135036 12260 297272 12288
rect 135036 12248 135042 12260
rect 297266 12248 297272 12260
rect 297324 12248 297330 12300
rect 136450 12180 136456 12232
rect 136508 12220 136514 12232
rect 299474 12220 299480 12232
rect 136508 12192 299480 12220
rect 136508 12180 136514 12192
rect 299474 12180 299480 12192
rect 299532 12180 299538 12232
rect 137830 12112 137836 12164
rect 137888 12152 137894 12164
rect 304350 12152 304356 12164
rect 137888 12124 304356 12152
rect 137888 12112 137894 12124
rect 304350 12112 304356 12124
rect 304408 12112 304414 12164
rect 137738 12044 137744 12096
rect 137796 12084 137802 12096
rect 307938 12084 307944 12096
rect 137796 12056 307944 12084
rect 137796 12044 137802 12056
rect 307938 12044 307944 12056
rect 307996 12044 308002 12096
rect 139118 11976 139124 12028
rect 139176 12016 139182 12028
rect 311434 12016 311440 12028
rect 139176 11988 311440 12016
rect 139176 11976 139182 11988
rect 311434 11976 311440 11988
rect 311492 11976 311498 12028
rect 139210 11908 139216 11960
rect 139268 11948 139274 11960
rect 315022 11948 315028 11960
rect 139268 11920 315028 11948
rect 139268 11908 139274 11920
rect 315022 11908 315028 11920
rect 315080 11908 315086 11960
rect 140682 11840 140688 11892
rect 140740 11880 140746 11892
rect 318518 11880 318524 11892
rect 140740 11852 318524 11880
rect 140740 11840 140746 11852
rect 318518 11840 318524 11852
rect 318576 11840 318582 11892
rect 141970 11772 141976 11824
rect 142028 11812 142034 11824
rect 322106 11812 322112 11824
rect 142028 11784 322112 11812
rect 142028 11772 142034 11784
rect 322106 11772 322112 11784
rect 322164 11772 322170 11824
rect 141786 11704 141792 11756
rect 141844 11744 141850 11756
rect 325602 11744 325608 11756
rect 141844 11716 325608 11744
rect 141844 11704 141850 11716
rect 325602 11704 325608 11716
rect 325660 11704 325666 11756
rect 357526 11704 357532 11756
rect 357584 11744 357590 11756
rect 358722 11744 358728 11756
rect 357584 11716 358728 11744
rect 357584 11704 357590 11716
rect 358722 11704 358728 11716
rect 358780 11704 358786 11756
rect 432046 11704 432052 11756
rect 432104 11744 432110 11756
rect 433242 11744 433248 11756
rect 432104 11716 433248 11744
rect 432104 11704 432110 11716
rect 433242 11704 433248 11716
rect 433300 11704 433306 11756
rect 132310 11636 132316 11688
rect 132368 11676 132374 11688
rect 286594 11676 286600 11688
rect 132368 11648 286600 11676
rect 132368 11636 132374 11648
rect 286594 11636 286600 11648
rect 286652 11636 286658 11688
rect 132218 11568 132224 11620
rect 132276 11608 132282 11620
rect 283098 11608 283104 11620
rect 132276 11580 283104 11608
rect 132276 11568 132282 11580
rect 283098 11568 283104 11580
rect 283156 11568 283162 11620
rect 130838 11500 130844 11552
rect 130896 11540 130902 11552
rect 279510 11540 279516 11552
rect 130896 11512 279516 11540
rect 130896 11500 130902 11512
rect 279510 11500 279516 11512
rect 279568 11500 279574 11552
rect 129458 11432 129464 11484
rect 129516 11472 129522 11484
rect 276106 11472 276112 11484
rect 129516 11444 276112 11472
rect 129516 11432 129522 11444
rect 276106 11432 276112 11444
rect 276164 11432 276170 11484
rect 129550 11364 129556 11416
rect 129608 11404 129614 11416
rect 272426 11404 272432 11416
rect 129608 11376 272432 11404
rect 129608 11364 129614 11376
rect 272426 11364 272432 11376
rect 272484 11364 272490 11416
rect 128078 11296 128084 11348
rect 128136 11336 128142 11348
rect 268838 11336 268844 11348
rect 128136 11308 268844 11336
rect 128136 11296 128142 11308
rect 268838 11296 268844 11308
rect 268896 11296 268902 11348
rect 126606 11228 126612 11280
rect 126664 11268 126670 11280
rect 265342 11268 265348 11280
rect 126664 11240 265348 11268
rect 126664 11228 126670 11240
rect 265342 11228 265348 11240
rect 265400 11228 265406 11280
rect 126698 11160 126704 11212
rect 126756 11200 126762 11212
rect 261754 11200 261760 11212
rect 126756 11172 261760 11200
rect 126756 11160 126762 11172
rect 261754 11160 261760 11172
rect 261812 11160 261818 11212
rect 107286 10956 107292 11008
rect 107344 10996 107350 11008
rect 187326 10996 187332 11008
rect 107344 10968 187332 10996
rect 107344 10956 107350 10968
rect 187326 10956 187332 10968
rect 187384 10956 187390 11008
rect 197078 10956 197084 11008
rect 197136 10996 197142 11008
rect 541986 10996 541992 11008
rect 197136 10968 541992 10996
rect 197136 10956 197142 10968
rect 541986 10956 541992 10968
rect 542044 10956 542050 11008
rect 107378 10888 107384 10940
rect 107436 10928 107442 10940
rect 188522 10928 188528 10940
rect 107436 10900 188528 10928
rect 107436 10888 107442 10900
rect 188522 10888 188528 10900
rect 188580 10888 188586 10940
rect 198458 10888 198464 10940
rect 198516 10928 198522 10940
rect 545482 10928 545488 10940
rect 198516 10900 545488 10928
rect 198516 10888 198522 10900
rect 545482 10888 545488 10900
rect 545540 10888 545546 10940
rect 108666 10820 108672 10872
rect 108724 10860 108730 10872
rect 190822 10860 190828 10872
rect 108724 10832 190828 10860
rect 108724 10820 108730 10832
rect 190822 10820 190828 10832
rect 190880 10820 190886 10872
rect 198550 10820 198556 10872
rect 198608 10860 198614 10872
rect 547874 10860 547880 10872
rect 198608 10832 547880 10860
rect 198608 10820 198614 10832
rect 547874 10820 547880 10832
rect 547932 10820 547938 10872
rect 108758 10752 108764 10804
rect 108816 10792 108822 10804
rect 192018 10792 192024 10804
rect 108816 10764 192024 10792
rect 108816 10752 108822 10764
rect 192018 10752 192024 10764
rect 192076 10752 192082 10804
rect 199838 10752 199844 10804
rect 199896 10792 199902 10804
rect 552658 10792 552664 10804
rect 199896 10764 552664 10792
rect 199896 10752 199902 10764
rect 552658 10752 552664 10764
rect 552716 10752 552722 10804
rect 110230 10684 110236 10736
rect 110288 10724 110294 10736
rect 195606 10724 195612 10736
rect 110288 10696 195612 10724
rect 110288 10684 110294 10696
rect 195606 10684 195612 10696
rect 195664 10684 195670 10736
rect 201218 10684 201224 10736
rect 201276 10724 201282 10736
rect 556154 10724 556160 10736
rect 201276 10696 556160 10724
rect 201276 10684 201282 10696
rect 556154 10684 556160 10696
rect 556212 10684 556218 10736
rect 108574 10616 108580 10668
rect 108632 10656 108638 10668
rect 193214 10656 193220 10668
rect 108632 10628 193220 10656
rect 108632 10616 108638 10628
rect 193214 10616 193220 10628
rect 193272 10616 193278 10668
rect 201310 10616 201316 10668
rect 201368 10656 201374 10668
rect 559742 10656 559748 10668
rect 201368 10628 559748 10656
rect 201368 10616 201374 10628
rect 559742 10616 559748 10628
rect 559800 10616 559806 10668
rect 110138 10548 110144 10600
rect 110196 10588 110202 10600
rect 197906 10588 197912 10600
rect 110196 10560 197912 10588
rect 110196 10548 110202 10560
rect 197906 10548 197912 10560
rect 197964 10548 197970 10600
rect 202506 10548 202512 10600
rect 202564 10548 202570 10600
rect 202598 10548 202604 10600
rect 202656 10588 202662 10600
rect 563238 10588 563244 10600
rect 202656 10560 563244 10588
rect 202656 10548 202662 10560
rect 563238 10548 563244 10560
rect 563296 10548 563302 10600
rect 110046 10480 110052 10532
rect 110104 10520 110110 10532
rect 199102 10520 199108 10532
rect 110104 10492 199108 10520
rect 110104 10480 110110 10492
rect 199102 10480 199108 10492
rect 199160 10480 199166 10532
rect 202524 10520 202552 10548
rect 566826 10520 566832 10532
rect 202524 10492 566832 10520
rect 566826 10480 566832 10492
rect 566884 10480 566890 10532
rect 111518 10412 111524 10464
rect 111576 10452 111582 10464
rect 202506 10452 202512 10464
rect 111576 10424 202512 10452
rect 111576 10412 111582 10424
rect 202506 10412 202512 10424
rect 202564 10412 202570 10464
rect 204070 10412 204076 10464
rect 204128 10452 204134 10464
rect 570322 10452 570328 10464
rect 204128 10424 570328 10452
rect 204128 10412 204134 10424
rect 570322 10412 570328 10424
rect 570380 10412 570386 10464
rect 111426 10344 111432 10396
rect 111484 10384 111490 10396
rect 201494 10384 201500 10396
rect 111484 10356 201500 10384
rect 111484 10344 111490 10356
rect 201494 10344 201500 10356
rect 201552 10344 201558 10396
rect 205358 10344 205364 10396
rect 205416 10384 205422 10396
rect 572714 10384 572720 10396
rect 205416 10356 572720 10384
rect 205416 10344 205422 10356
rect 572714 10344 572720 10356
rect 572772 10344 572778 10396
rect 88150 10276 88156 10328
rect 88208 10316 88214 10328
rect 106918 10316 106924 10328
rect 88208 10288 106924 10316
rect 88208 10276 88214 10288
rect 106918 10276 106924 10288
rect 106976 10276 106982 10328
rect 111334 10276 111340 10328
rect 111392 10316 111398 10328
rect 205082 10316 205088 10328
rect 111392 10288 205088 10316
rect 111392 10276 111398 10288
rect 205082 10276 205088 10288
rect 205140 10276 205146 10328
rect 205266 10276 205272 10328
rect 205324 10316 205330 10328
rect 577406 10316 577412 10328
rect 205324 10288 577412 10316
rect 205324 10276 205330 10288
rect 577406 10276 577412 10288
rect 577464 10276 577470 10328
rect 195790 10208 195796 10260
rect 195848 10248 195854 10260
rect 538398 10248 538404 10260
rect 195848 10220 538404 10248
rect 195848 10208 195854 10220
rect 538398 10208 538404 10220
rect 538456 10208 538462 10260
rect 195698 10140 195704 10192
rect 195756 10180 195762 10192
rect 534902 10180 534908 10192
rect 195756 10152 534908 10180
rect 195756 10140 195762 10152
rect 534902 10140 534908 10152
rect 534960 10140 534966 10192
rect 114370 10072 114376 10124
rect 114428 10112 114434 10124
rect 215662 10112 215668 10124
rect 114428 10084 215668 10112
rect 114428 10072 114434 10084
rect 215662 10072 215668 10084
rect 215720 10072 215726 10124
rect 215938 10072 215944 10124
rect 215996 10112 216002 10124
rect 372890 10112 372896 10124
rect 215996 10084 372896 10112
rect 215996 10072 216002 10084
rect 372890 10072 372896 10084
rect 372948 10072 372954 10124
rect 117130 10004 117136 10056
rect 117188 10044 117194 10056
rect 226426 10044 226432 10056
rect 117188 10016 226432 10044
rect 117188 10004 117194 10016
rect 226426 10004 226432 10016
rect 226484 10004 226490 10056
rect 116854 9936 116860 9988
rect 116912 9976 116918 9988
rect 222746 9976 222752 9988
rect 116912 9948 222752 9976
rect 116912 9936 116918 9948
rect 222746 9936 222752 9948
rect 222804 9936 222810 9988
rect 115474 9868 115480 9920
rect 115532 9908 115538 9920
rect 219250 9908 219256 9920
rect 115532 9880 219256 9908
rect 115532 9868 115538 9880
rect 219250 9868 219256 9880
rect 219308 9868 219314 9920
rect 114462 9800 114468 9852
rect 114520 9840 114526 9852
rect 212166 9840 212172 9852
rect 114520 9812 212172 9840
rect 114520 9800 114526 9812
rect 212166 9800 212172 9812
rect 212224 9800 212230 9852
rect 112806 9732 112812 9784
rect 112864 9772 112870 9784
rect 208578 9772 208584 9784
rect 112864 9744 208584 9772
rect 112864 9732 112870 9744
rect 208578 9732 208584 9744
rect 208636 9732 208642 9784
rect 176378 9596 176384 9648
rect 176436 9636 176442 9648
rect 462774 9636 462780 9648
rect 176436 9608 462780 9636
rect 176436 9596 176442 9608
rect 462774 9596 462780 9608
rect 462832 9596 462838 9648
rect 101858 9528 101864 9580
rect 101916 9568 101922 9580
rect 163682 9568 163688 9580
rect 101916 9540 163688 9568
rect 101916 9528 101922 9540
rect 163682 9528 163688 9540
rect 163740 9528 163746 9580
rect 177850 9528 177856 9580
rect 177908 9568 177914 9580
rect 466270 9568 466276 9580
rect 177908 9540 466276 9568
rect 177908 9528 177914 9540
rect 466270 9528 466276 9540
rect 466328 9528 466334 9580
rect 101766 9460 101772 9512
rect 101824 9500 101830 9512
rect 167178 9500 167184 9512
rect 101824 9472 167184 9500
rect 101824 9460 101830 9472
rect 167178 9460 167184 9472
rect 167236 9460 167242 9512
rect 179230 9460 179236 9512
rect 179288 9500 179294 9512
rect 469858 9500 469864 9512
rect 179288 9472 469864 9500
rect 179288 9460 179294 9472
rect 469858 9460 469864 9472
rect 469916 9460 469922 9512
rect 103330 9392 103336 9444
rect 103388 9432 103394 9444
rect 170766 9432 170772 9444
rect 103388 9404 170772 9432
rect 103388 9392 103394 9404
rect 170766 9392 170772 9404
rect 170824 9392 170830 9444
rect 179138 9392 179144 9444
rect 179196 9432 179202 9444
rect 473446 9432 473452 9444
rect 179196 9404 473452 9432
rect 179196 9392 179202 9404
rect 473446 9392 473452 9404
rect 473504 9392 473510 9444
rect 104710 9324 104716 9376
rect 104768 9364 104774 9376
rect 174262 9364 174268 9376
rect 104768 9336 174268 9364
rect 104768 9324 104774 9336
rect 174262 9324 174268 9336
rect 174320 9324 174326 9376
rect 180702 9324 180708 9376
rect 180760 9364 180766 9376
rect 476942 9364 476948 9376
rect 180760 9336 476948 9364
rect 180760 9324 180766 9336
rect 476942 9324 476948 9336
rect 477000 9324 477006 9376
rect 104618 9256 104624 9308
rect 104676 9296 104682 9308
rect 177850 9296 177856 9308
rect 104676 9268 177856 9296
rect 104676 9256 104682 9268
rect 177850 9256 177856 9268
rect 177908 9256 177914 9308
rect 181898 9256 181904 9308
rect 181956 9296 181962 9308
rect 481726 9296 481732 9308
rect 181956 9268 481732 9296
rect 181956 9256 181962 9268
rect 481726 9256 481732 9268
rect 481784 9256 481790 9308
rect 104526 9188 104532 9240
rect 104584 9228 104590 9240
rect 176654 9228 176660 9240
rect 104584 9200 176660 9228
rect 104584 9188 104590 9200
rect 176654 9188 176660 9200
rect 176712 9188 176718 9240
rect 183370 9188 183376 9240
rect 183428 9228 183434 9240
rect 485222 9228 485228 9240
rect 183428 9200 485228 9228
rect 183428 9188 183434 9200
rect 485222 9188 485228 9200
rect 485280 9188 485286 9240
rect 106182 9120 106188 9172
rect 106240 9160 106246 9172
rect 180242 9160 180248 9172
rect 106240 9132 180248 9160
rect 106240 9120 106246 9132
rect 180242 9120 180248 9132
rect 180300 9120 180306 9172
rect 183094 9120 183100 9172
rect 183152 9160 183158 9172
rect 488810 9160 488816 9172
rect 183152 9132 488816 9160
rect 183152 9120 183158 9132
rect 488810 9120 488816 9132
rect 488868 9120 488874 9172
rect 106090 9052 106096 9104
rect 106148 9092 106154 9104
rect 181438 9092 181444 9104
rect 106148 9064 181444 9092
rect 106148 9052 106154 9064
rect 181438 9052 181444 9064
rect 181496 9052 181502 9104
rect 184658 9052 184664 9104
rect 184716 9092 184722 9104
rect 492306 9092 492312 9104
rect 184716 9064 492312 9092
rect 184716 9052 184722 9064
rect 492306 9052 492312 9064
rect 492364 9052 492370 9104
rect 107562 8984 107568 9036
rect 107620 9024 107626 9036
rect 183738 9024 183744 9036
rect 107620 8996 183744 9024
rect 107620 8984 107626 8996
rect 183738 8984 183744 8996
rect 183796 8984 183802 9036
rect 185854 8984 185860 9036
rect 185912 9024 185918 9036
rect 495894 9024 495900 9036
rect 185912 8996 495900 9024
rect 185912 8984 185918 8996
rect 495894 8984 495900 8996
rect 495952 8984 495958 9036
rect 107470 8916 107476 8968
rect 107528 8956 107534 8968
rect 184934 8956 184940 8968
rect 107528 8928 184940 8956
rect 107528 8916 107534 8928
rect 184934 8916 184940 8928
rect 184992 8916 184998 8968
rect 186130 8916 186136 8968
rect 186188 8956 186194 8968
rect 499390 8956 499396 8968
rect 186188 8928 499396 8956
rect 186188 8916 186194 8928
rect 499390 8916 499396 8928
rect 499448 8916 499454 8968
rect 176470 8848 176476 8900
rect 176528 8888 176534 8900
rect 459186 8888 459192 8900
rect 176528 8860 459192 8888
rect 176528 8848 176534 8860
rect 459186 8848 459192 8860
rect 459244 8848 459250 8900
rect 175182 8780 175188 8832
rect 175240 8820 175246 8832
rect 455690 8820 455696 8832
rect 175240 8792 455696 8820
rect 175240 8780 175246 8792
rect 455690 8780 455696 8792
rect 455748 8780 455754 8832
rect 175090 8712 175096 8764
rect 175148 8752 175154 8764
rect 452102 8752 452108 8764
rect 175148 8724 452108 8752
rect 175148 8712 175154 8724
rect 452102 8712 452108 8724
rect 452160 8712 452166 8764
rect 173802 8644 173808 8696
rect 173860 8684 173866 8696
rect 448606 8684 448612 8696
rect 173860 8656 448612 8684
rect 173860 8644 173866 8656
rect 448606 8644 448612 8656
rect 448664 8644 448670 8696
rect 172330 8576 172336 8628
rect 172388 8616 172394 8628
rect 445018 8616 445024 8628
rect 172388 8588 445024 8616
rect 172388 8576 172394 8588
rect 445018 8576 445024 8588
rect 445076 8576 445082 8628
rect 172238 8508 172244 8560
rect 172296 8548 172302 8560
rect 441522 8548 441528 8560
rect 172296 8520 441528 8548
rect 172296 8508 172302 8520
rect 441522 8508 441528 8520
rect 441580 8508 441586 8560
rect 171042 8440 171048 8492
rect 171100 8480 171106 8492
rect 437934 8480 437940 8492
rect 171100 8452 437940 8480
rect 171100 8440 171106 8452
rect 437934 8440 437940 8452
rect 437992 8440 437998 8492
rect 169662 8372 169668 8424
rect 169720 8412 169726 8424
rect 434438 8412 434444 8424
rect 169720 8384 434444 8412
rect 169720 8372 169726 8384
rect 434438 8372 434444 8384
rect 434496 8372 434502 8424
rect 151630 8236 151636 8288
rect 151688 8276 151694 8288
rect 363506 8276 363512 8288
rect 151688 8248 363512 8276
rect 151688 8236 151694 8248
rect 363506 8236 363512 8248
rect 363564 8236 363570 8288
rect 153102 8168 153108 8220
rect 153160 8208 153166 8220
rect 367002 8208 367008 8220
rect 153160 8180 367008 8208
rect 153160 8168 153166 8180
rect 367002 8168 367008 8180
rect 367060 8168 367066 8220
rect 154482 8100 154488 8152
rect 154540 8140 154546 8152
rect 370590 8140 370596 8152
rect 154540 8112 370596 8140
rect 154540 8100 154546 8112
rect 370590 8100 370596 8112
rect 370648 8100 370654 8152
rect 154390 8032 154396 8084
rect 154448 8072 154454 8084
rect 374086 8072 374092 8084
rect 154448 8044 374092 8072
rect 154448 8032 154454 8044
rect 374086 8032 374092 8044
rect 374144 8032 374150 8084
rect 155586 7964 155592 8016
rect 155644 8004 155650 8016
rect 377674 8004 377680 8016
rect 155644 7976 377680 8004
rect 155644 7964 155650 7976
rect 377674 7964 377680 7976
rect 377732 7964 377738 8016
rect 157150 7896 157156 7948
rect 157208 7936 157214 7948
rect 381170 7936 381176 7948
rect 157208 7908 381176 7936
rect 157208 7896 157214 7908
rect 381170 7896 381176 7908
rect 381228 7896 381234 7948
rect 95050 7828 95056 7880
rect 95108 7868 95114 7880
rect 137646 7868 137652 7880
rect 95108 7840 137652 7868
rect 95108 7828 95114 7840
rect 137646 7828 137652 7840
rect 137704 7828 137710 7880
rect 157242 7828 157248 7880
rect 157300 7868 157306 7880
rect 384758 7868 384764 7880
rect 157300 7840 384764 7868
rect 157300 7828 157306 7840
rect 384758 7828 384764 7840
rect 384816 7828 384822 7880
rect 96338 7760 96344 7812
rect 96396 7800 96402 7812
rect 141234 7800 141240 7812
rect 96396 7772 141240 7800
rect 96396 7760 96402 7772
rect 141234 7760 141240 7772
rect 141292 7760 141298 7812
rect 158622 7760 158628 7812
rect 158680 7800 158686 7812
rect 388254 7800 388260 7812
rect 158680 7772 388260 7800
rect 158680 7760 158686 7772
rect 388254 7760 388260 7772
rect 388312 7760 388318 7812
rect 99098 7692 99104 7744
rect 99156 7732 99162 7744
rect 151814 7732 151820 7744
rect 99156 7704 151820 7732
rect 99156 7692 99162 7704
rect 151814 7692 151820 7704
rect 151872 7692 151878 7744
rect 159634 7692 159640 7744
rect 159692 7732 159698 7744
rect 391842 7732 391848 7744
rect 159692 7704 391848 7732
rect 159692 7692 159698 7704
rect 391842 7692 391848 7704
rect 391900 7692 391906 7744
rect 99190 7624 99196 7676
rect 99248 7664 99254 7676
rect 155402 7664 155408 7676
rect 99248 7636 155408 7664
rect 99248 7624 99254 7636
rect 155402 7624 155408 7636
rect 155460 7624 155466 7676
rect 159910 7624 159916 7676
rect 159968 7664 159974 7676
rect 395338 7664 395344 7676
rect 159968 7636 395344 7664
rect 159968 7624 159974 7636
rect 395338 7624 395344 7636
rect 395396 7624 395402 7676
rect 100478 7556 100484 7608
rect 100536 7596 100542 7608
rect 158898 7596 158904 7608
rect 100536 7568 158904 7596
rect 100536 7556 100542 7568
rect 158898 7556 158904 7568
rect 158956 7556 158962 7608
rect 161382 7556 161388 7608
rect 161440 7596 161446 7608
rect 398926 7596 398932 7608
rect 161440 7568 398932 7596
rect 161440 7556 161446 7568
rect 398926 7556 398932 7568
rect 398984 7556 398990 7608
rect 151722 7488 151728 7540
rect 151780 7528 151786 7540
rect 359918 7528 359924 7540
rect 151780 7500 359924 7528
rect 151780 7488 151786 7500
rect 359918 7488 359924 7500
rect 359976 7488 359982 7540
rect 150342 7420 150348 7472
rect 150400 7460 150406 7472
rect 356330 7460 356336 7472
rect 150400 7432 356336 7460
rect 150400 7420 150406 7432
rect 356330 7420 356336 7432
rect 356388 7420 356394 7472
rect 148870 7352 148876 7404
rect 148928 7392 148934 7404
rect 352834 7392 352840 7404
rect 148928 7364 352840 7392
rect 148928 7352 148934 7364
rect 352834 7352 352840 7364
rect 352892 7352 352898 7404
rect 148962 7284 148968 7336
rect 149020 7324 149026 7336
rect 349246 7324 349252 7336
rect 149020 7296 349252 7324
rect 149020 7284 149026 7296
rect 349246 7284 349252 7296
rect 349304 7284 349310 7336
rect 147582 7216 147588 7268
rect 147640 7256 147646 7268
rect 345750 7256 345756 7268
rect 147640 7228 345756 7256
rect 147640 7216 147646 7228
rect 345750 7216 345756 7228
rect 345808 7216 345814 7268
rect 146110 7148 146116 7200
rect 146168 7188 146174 7200
rect 342162 7188 342168 7200
rect 146168 7160 342168 7188
rect 146168 7148 146174 7160
rect 342162 7148 342168 7160
rect 342220 7148 342226 7200
rect 146202 7080 146208 7132
rect 146260 7120 146266 7132
rect 338666 7120 338672 7132
rect 146260 7092 338672 7120
rect 146260 7080 146266 7092
rect 338666 7080 338672 7092
rect 338724 7080 338730 7132
rect 144822 7012 144828 7064
rect 144880 7052 144886 7064
rect 335078 7052 335084 7064
rect 144880 7024 335084 7052
rect 144880 7012 144886 7024
rect 335078 7012 335084 7024
rect 335136 7012 335142 7064
rect 126790 6808 126796 6860
rect 126848 6848 126854 6860
rect 264146 6848 264152 6860
rect 126848 6820 264152 6848
rect 126848 6808 126854 6820
rect 264146 6808 264152 6820
rect 264204 6808 264210 6860
rect 128170 6740 128176 6792
rect 128228 6780 128234 6792
rect 267734 6780 267740 6792
rect 128228 6752 267740 6780
rect 128228 6740 128234 6752
rect 267734 6740 267740 6752
rect 267792 6740 267798 6792
rect 128262 6672 128268 6724
rect 128320 6712 128326 6724
rect 271230 6712 271236 6724
rect 128320 6684 271236 6712
rect 128320 6672 128326 6684
rect 271230 6672 271236 6684
rect 271288 6672 271294 6724
rect 129642 6604 129648 6656
rect 129700 6644 129706 6656
rect 274818 6644 274824 6656
rect 129700 6616 274824 6644
rect 129700 6604 129706 6616
rect 274818 6604 274824 6616
rect 274876 6604 274882 6656
rect 130930 6536 130936 6588
rect 130988 6576 130994 6588
rect 278314 6576 278320 6588
rect 130988 6548 278320 6576
rect 130988 6536 130994 6548
rect 278314 6536 278320 6548
rect 278372 6536 278378 6588
rect 131022 6468 131028 6520
rect 131080 6508 131086 6520
rect 281902 6508 281908 6520
rect 131080 6480 281908 6508
rect 131080 6468 131086 6480
rect 281902 6468 281908 6480
rect 281960 6468 281966 6520
rect 132402 6400 132408 6452
rect 132460 6440 132466 6452
rect 285398 6440 285404 6452
rect 132460 6412 285404 6440
rect 132460 6400 132466 6412
rect 285398 6400 285404 6412
rect 285456 6400 285462 6452
rect 133690 6332 133696 6384
rect 133748 6372 133754 6384
rect 288986 6372 288992 6384
rect 133748 6344 288992 6372
rect 133748 6332 133754 6344
rect 288986 6332 288992 6344
rect 289044 6332 289050 6384
rect 105630 6264 105636 6316
rect 105688 6304 105694 6316
rect 128170 6304 128176 6316
rect 105688 6276 128176 6304
rect 105688 6264 105694 6276
rect 128170 6264 128176 6276
rect 128228 6264 128234 6316
rect 133782 6264 133788 6316
rect 133840 6304 133846 6316
rect 292574 6304 292580 6316
rect 133840 6276 292580 6304
rect 133840 6264 133846 6276
rect 292574 6264 292580 6276
rect 292632 6264 292638 6316
rect 93578 6196 93584 6248
rect 93636 6236 93642 6248
rect 130562 6236 130568 6248
rect 93636 6208 130568 6236
rect 93636 6196 93642 6208
rect 130562 6196 130568 6208
rect 130620 6196 130626 6248
rect 135162 6196 135168 6248
rect 135220 6236 135226 6248
rect 296070 6236 296076 6248
rect 135220 6208 296076 6236
rect 135220 6196 135226 6208
rect 296070 6196 296076 6208
rect 296128 6196 296134 6248
rect 93486 6128 93492 6180
rect 93544 6168 93550 6180
rect 134150 6168 134156 6180
rect 93544 6140 134156 6168
rect 93544 6128 93550 6140
rect 134150 6128 134156 6140
rect 134208 6128 134214 6180
rect 136542 6128 136548 6180
rect 136600 6168 136606 6180
rect 299658 6168 299664 6180
rect 136600 6140 299664 6168
rect 136600 6128 136606 6140
rect 299658 6128 299664 6140
rect 299716 6128 299722 6180
rect 126882 6060 126888 6112
rect 126940 6100 126946 6112
rect 260650 6100 260656 6112
rect 126940 6072 260656 6100
rect 126940 6060 126946 6072
rect 260650 6060 260656 6072
rect 260708 6060 260714 6112
rect 125226 5992 125232 6044
rect 125284 6032 125290 6044
rect 257062 6032 257068 6044
rect 125284 6004 257068 6032
rect 125284 5992 125290 6004
rect 257062 5992 257068 6004
rect 257120 5992 257126 6044
rect 123754 5924 123760 5976
rect 123812 5964 123818 5976
rect 253474 5964 253480 5976
rect 123812 5936 253480 5964
rect 123812 5924 123818 5936
rect 253474 5924 253480 5936
rect 253532 5924 253538 5976
rect 124030 5856 124036 5908
rect 124088 5896 124094 5908
rect 249978 5896 249984 5908
rect 124088 5868 249984 5896
rect 124088 5856 124094 5868
rect 249978 5856 249984 5868
rect 250036 5856 250042 5908
rect 122742 5788 122748 5840
rect 122800 5828 122806 5840
rect 246390 5828 246396 5840
rect 122800 5800 246396 5828
rect 122800 5788 122806 5800
rect 246390 5788 246396 5800
rect 246448 5788 246454 5840
rect 121362 5720 121368 5772
rect 121420 5760 121426 5772
rect 242986 5760 242992 5772
rect 121420 5732 242992 5760
rect 121420 5720 121426 5732
rect 242986 5720 242992 5732
rect 243044 5720 243050 5772
rect 121270 5652 121276 5704
rect 121328 5692 121334 5704
rect 239306 5692 239312 5704
rect 121328 5664 239312 5692
rect 121328 5652 121334 5664
rect 239306 5652 239312 5664
rect 239364 5652 239370 5704
rect 119614 5584 119620 5636
rect 119672 5624 119678 5636
rect 235810 5624 235816 5636
rect 119672 5596 235816 5624
rect 119672 5584 119678 5596
rect 235810 5584 235816 5596
rect 235868 5584 235874 5636
rect 99282 5448 99288 5500
rect 99340 5488 99346 5500
rect 154206 5488 154212 5500
rect 99340 5460 154212 5488
rect 99340 5448 99346 5460
rect 154206 5448 154212 5460
rect 154264 5448 154270 5500
rect 196894 5448 196900 5500
rect 196952 5488 196958 5500
rect 540790 5488 540796 5500
rect 196952 5460 540796 5488
rect 196952 5448 196958 5460
rect 540790 5448 540796 5460
rect 540848 5448 540854 5500
rect 100570 5380 100576 5432
rect 100628 5420 100634 5432
rect 157794 5420 157800 5432
rect 100628 5392 157800 5420
rect 100628 5380 100634 5392
rect 157794 5380 157800 5392
rect 157852 5380 157858 5432
rect 197170 5380 197176 5432
rect 197228 5420 197234 5432
rect 544286 5420 544292 5432
rect 197228 5392 544292 5420
rect 197228 5380 197234 5392
rect 544286 5380 544292 5392
rect 544344 5380 544350 5432
rect 102042 5312 102048 5364
rect 102100 5352 102106 5364
rect 162486 5352 162492 5364
rect 102100 5324 162492 5352
rect 102100 5312 102106 5324
rect 162486 5312 162492 5324
rect 162544 5312 162550 5364
rect 198274 5312 198280 5364
rect 198332 5352 198338 5364
rect 547966 5352 547972 5364
rect 198332 5324 547972 5352
rect 198332 5312 198338 5324
rect 547966 5312 547972 5324
rect 548024 5312 548030 5364
rect 101950 5244 101956 5296
rect 102008 5284 102014 5296
rect 166074 5284 166080 5296
rect 102008 5256 166080 5284
rect 102008 5244 102014 5256
rect 166074 5244 166080 5256
rect 166132 5244 166138 5296
rect 199930 5244 199936 5296
rect 199988 5284 199994 5296
rect 551462 5284 551468 5296
rect 199988 5256 551468 5284
rect 199988 5244 199994 5256
rect 551462 5244 551468 5256
rect 551520 5244 551526 5296
rect 103422 5176 103428 5228
rect 103480 5216 103486 5228
rect 169570 5216 169576 5228
rect 103480 5188 169576 5216
rect 103480 5176 103486 5188
rect 169570 5176 169576 5188
rect 169628 5176 169634 5228
rect 200022 5176 200028 5228
rect 200080 5216 200086 5228
rect 554958 5216 554964 5228
rect 200080 5188 554964 5216
rect 200080 5176 200086 5188
rect 554958 5176 554964 5188
rect 555016 5176 555022 5228
rect 104802 5108 104808 5160
rect 104860 5148 104866 5160
rect 173158 5148 173164 5160
rect 104860 5120 173164 5148
rect 104860 5108 104866 5120
rect 173158 5108 173164 5120
rect 173216 5108 173222 5160
rect 202598 5108 202604 5160
rect 202656 5148 202662 5160
rect 205085 5151 205143 5157
rect 205085 5148 205097 5151
rect 202656 5120 205097 5148
rect 202656 5108 202662 5120
rect 205085 5117 205097 5120
rect 205131 5117 205143 5151
rect 205085 5111 205143 5117
rect 205177 5151 205235 5157
rect 205177 5117 205189 5151
rect 205223 5148 205235 5151
rect 558546 5148 558552 5160
rect 205223 5120 558552 5148
rect 205223 5117 205235 5120
rect 205177 5111 205235 5117
rect 558546 5108 558552 5120
rect 558604 5108 558610 5160
rect 108942 5040 108948 5092
rect 109000 5080 109006 5092
rect 189718 5080 189724 5092
rect 109000 5052 189724 5080
rect 109000 5040 109006 5052
rect 189718 5040 189724 5052
rect 189776 5040 189782 5092
rect 202782 5040 202788 5092
rect 202840 5080 202846 5092
rect 562042 5080 562048 5092
rect 202840 5052 562048 5080
rect 202840 5040 202846 5052
rect 562042 5040 562048 5052
rect 562100 5040 562106 5092
rect 108850 4972 108856 5024
rect 108908 5012 108914 5024
rect 193306 5012 193312 5024
rect 108908 4984 193312 5012
rect 108908 4972 108914 4984
rect 193306 4972 193312 4984
rect 193364 4972 193370 5024
rect 194134 4972 194140 5024
rect 194192 5012 194198 5024
rect 204993 5015 205051 5021
rect 204993 5012 205005 5015
rect 194192 4984 205005 5012
rect 194192 4972 194198 4984
rect 204993 4981 205005 4984
rect 205039 4981 205051 5015
rect 204993 4975 205051 4981
rect 205085 5015 205143 5021
rect 205085 4981 205097 5015
rect 205131 5012 205143 5015
rect 565630 5012 565636 5024
rect 205131 4984 565636 5012
rect 205131 4981 205143 4984
rect 205085 4975 205143 4981
rect 565630 4972 565636 4984
rect 565688 4972 565694 5024
rect 110322 4904 110328 4956
rect 110380 4944 110386 4956
rect 196802 4944 196808 4956
rect 110380 4916 196808 4944
rect 110380 4904 110386 4916
rect 196802 4904 196808 4916
rect 196860 4904 196866 4956
rect 204162 4904 204168 4956
rect 204220 4944 204226 4956
rect 569126 4944 569132 4956
rect 204220 4916 569132 4944
rect 204220 4904 204226 4916
rect 569126 4904 569132 4916
rect 569184 4904 569190 4956
rect 111702 4836 111708 4888
rect 111760 4876 111766 4888
rect 195241 4879 195299 4885
rect 195241 4876 195253 4879
rect 111760 4848 195253 4876
rect 111760 4836 111766 4848
rect 195241 4845 195253 4848
rect 195287 4845 195299 4879
rect 195241 4839 195299 4845
rect 201034 4836 201040 4888
rect 201092 4876 201098 4888
rect 205177 4879 205235 4885
rect 205177 4876 205189 4879
rect 201092 4848 205189 4876
rect 201092 4836 201098 4848
rect 205177 4845 205189 4848
rect 205223 4845 205235 4879
rect 205177 4839 205235 4845
rect 205542 4836 205548 4888
rect 205600 4876 205606 4888
rect 572806 4876 572812 4888
rect 205600 4848 572812 4876
rect 205600 4836 205606 4848
rect 572806 4836 572812 4848
rect 572864 4836 572870 4888
rect 62022 4768 62028 4820
rect 62080 4808 62086 4820
rect 71038 4808 71044 4820
rect 62080 4780 71044 4808
rect 62080 4768 62086 4780
rect 71038 4768 71044 4780
rect 71096 4768 71102 4820
rect 111610 4768 111616 4820
rect 111668 4808 111674 4820
rect 203886 4808 203892 4820
rect 111668 4780 203892 4808
rect 111668 4768 111674 4780
rect 203886 4768 203892 4780
rect 203944 4768 203950 4820
rect 205450 4768 205456 4820
rect 205508 4808 205514 4820
rect 576302 4808 576308 4820
rect 205508 4780 576308 4808
rect 205508 4768 205514 4780
rect 576302 4768 576308 4780
rect 576360 4768 576366 4820
rect 97810 4700 97816 4752
rect 97868 4740 97874 4752
rect 150618 4740 150624 4752
rect 97868 4712 150624 4740
rect 97868 4700 97874 4712
rect 150618 4700 150624 4712
rect 150676 4700 150682 4752
rect 195241 4743 195299 4749
rect 195241 4709 195253 4743
rect 195287 4740 195299 4743
rect 200298 4740 200304 4752
rect 195287 4712 200304 4740
rect 195287 4709 195299 4712
rect 195241 4703 195299 4709
rect 200298 4700 200304 4712
rect 200356 4700 200362 4752
rect 537202 4740 537208 4752
rect 204916 4712 537208 4740
rect 93394 4632 93400 4684
rect 93452 4672 93458 4684
rect 132954 4672 132960 4684
rect 93452 4644 132960 4672
rect 93452 4632 93458 4644
rect 132954 4632 132960 4644
rect 133012 4632 133018 4684
rect 133138 4632 133144 4684
rect 133196 4672 133202 4684
rect 186130 4672 186136 4684
rect 133196 4644 186136 4672
rect 133196 4632 133202 4644
rect 186130 4632 186136 4644
rect 186188 4632 186194 4684
rect 195882 4632 195888 4684
rect 195940 4672 195946 4684
rect 204916 4672 204944 4712
rect 537202 4700 537208 4712
rect 537260 4700 537266 4752
rect 195940 4644 204944 4672
rect 204993 4675 205051 4681
rect 195940 4632 195946 4644
rect 204993 4641 205005 4675
rect 205039 4672 205051 4675
rect 533706 4672 533712 4684
rect 205039 4644 533712 4672
rect 205039 4641 205051 4644
rect 204993 4635 205051 4641
rect 533706 4632 533712 4644
rect 533764 4632 533770 4684
rect 97902 4564 97908 4616
rect 97960 4604 97966 4616
rect 147030 4604 147036 4616
rect 97960 4576 147036 4604
rect 97960 4564 97966 4576
rect 147030 4564 147036 4576
rect 147088 4564 147094 4616
rect 148318 4564 148324 4616
rect 148376 4604 148382 4616
rect 175458 4604 175464 4616
rect 148376 4576 175464 4604
rect 148376 4564 148382 4576
rect 175458 4564 175464 4576
rect 175516 4564 175522 4616
rect 194502 4564 194508 4616
rect 194560 4604 194566 4616
rect 530118 4604 530124 4616
rect 194560 4576 530124 4604
rect 194560 4564 194566 4576
rect 530118 4564 530124 4576
rect 530176 4564 530182 4616
rect 96430 4496 96436 4548
rect 96488 4536 96494 4548
rect 143534 4536 143540 4548
rect 96488 4508 143540 4536
rect 96488 4496 96494 4508
rect 143534 4496 143540 4508
rect 143592 4496 143598 4548
rect 192846 4496 192852 4548
rect 192904 4536 192910 4548
rect 526622 4536 526628 4548
rect 192904 4508 526628 4536
rect 192904 4496 192910 4508
rect 526622 4496 526628 4508
rect 526680 4496 526686 4548
rect 96522 4428 96528 4480
rect 96580 4468 96586 4480
rect 140038 4468 140044 4480
rect 96580 4440 140044 4468
rect 96580 4428 96586 4440
rect 140038 4428 140044 4440
rect 140096 4428 140102 4480
rect 140130 4428 140136 4480
rect 140188 4468 140194 4480
rect 179046 4468 179052 4480
rect 140188 4440 179052 4468
rect 140188 4428 140194 4440
rect 179046 4428 179052 4440
rect 179104 4428 179110 4480
rect 191650 4428 191656 4480
rect 191708 4468 191714 4480
rect 523034 4468 523040 4480
rect 191708 4440 523040 4468
rect 191708 4428 191714 4440
rect 523034 4428 523040 4440
rect 523092 4428 523098 4480
rect 95142 4360 95148 4412
rect 95200 4400 95206 4412
rect 136450 4400 136456 4412
rect 95200 4372 136456 4400
rect 95200 4360 95206 4372
rect 136450 4360 136456 4372
rect 136508 4360 136514 4412
rect 191374 4360 191380 4412
rect 191432 4400 191438 4412
rect 519538 4400 519544 4412
rect 191432 4372 519544 4400
rect 191432 4360 191438 4372
rect 519538 4360 519544 4372
rect 519596 4360 519602 4412
rect 92290 4292 92296 4344
rect 92348 4332 92354 4344
rect 126974 4332 126980 4344
rect 92348 4304 126980 4332
rect 92348 4292 92354 4304
rect 126974 4292 126980 4304
rect 127032 4292 127038 4344
rect 190270 4292 190276 4344
rect 190328 4332 190334 4344
rect 515950 4332 515956 4344
rect 190328 4304 515956 4332
rect 190328 4292 190334 4304
rect 515950 4292 515956 4304
rect 516008 4292 516014 4344
rect 93670 4224 93676 4276
rect 93728 4264 93734 4276
rect 129366 4264 129372 4276
rect 93728 4236 129372 4264
rect 93728 4224 93734 4236
rect 129366 4224 129372 4236
rect 129424 4224 129430 4276
rect 190086 4224 190092 4276
rect 190144 4264 190150 4276
rect 512454 4264 512460 4276
rect 190144 4236 512460 4264
rect 190144 4224 190150 4236
rect 512454 4224 512460 4236
rect 512512 4224 512518 4276
rect 59924 4168 60136 4196
rect 43070 4088 43076 4140
rect 43128 4128 43134 4140
rect 59817 4131 59875 4137
rect 59817 4128 59829 4131
rect 43128 4100 59829 4128
rect 43128 4088 43134 4100
rect 59817 4097 59829 4100
rect 59863 4097 59875 4131
rect 59817 4091 59875 4097
rect 38378 4020 38384 4072
rect 38436 4060 38442 4072
rect 59924 4060 59952 4168
rect 60108 4128 60136 4168
rect 87690 4156 87696 4208
rect 87748 4196 87754 4208
rect 90358 4196 90364 4208
rect 87748 4168 90364 4196
rect 87748 4156 87754 4168
rect 90358 4156 90364 4168
rect 90416 4156 90422 4208
rect 98638 4156 98644 4208
rect 98696 4196 98702 4208
rect 101030 4196 101036 4208
rect 98696 4168 101036 4196
rect 98696 4156 98702 4168
rect 101030 4156 101036 4168
rect 101088 4156 101094 4208
rect 105538 4156 105544 4208
rect 105596 4196 105602 4208
rect 108114 4196 108120 4208
rect 105596 4168 108120 4196
rect 105596 4156 105602 4168
rect 108114 4156 108120 4168
rect 108172 4156 108178 4208
rect 64138 4128 64144 4140
rect 60108 4100 64144 4128
rect 64138 4088 64144 4100
rect 64196 4088 64202 4140
rect 64233 4131 64291 4137
rect 64233 4097 64245 4131
rect 64279 4128 64291 4131
rect 65518 4128 65524 4140
rect 64279 4100 65524 4128
rect 64279 4097 64291 4100
rect 64233 4091 64291 4097
rect 65518 4088 65524 4100
rect 65576 4088 65582 4140
rect 89438 4088 89444 4140
rect 89496 4128 89502 4140
rect 89496 4100 112392 4128
rect 89496 4088 89502 4100
rect 38436 4032 59952 4060
rect 60001 4063 60059 4069
rect 38436 4020 38442 4032
rect 60001 4029 60013 4063
rect 60047 4060 60059 4063
rect 67082 4060 67088 4072
rect 60047 4032 67088 4060
rect 60047 4029 60059 4032
rect 60001 4023 60059 4029
rect 67082 4020 67088 4032
rect 67140 4020 67146 4072
rect 89530 4020 89536 4072
rect 89588 4060 89594 4072
rect 111705 4063 111763 4069
rect 111705 4060 111717 4063
rect 89588 4032 111717 4060
rect 89588 4020 89594 4032
rect 111705 4029 111717 4032
rect 111751 4029 111763 4063
rect 112364 4060 112392 4100
rect 112438 4088 112444 4140
rect 112496 4128 112502 4140
rect 131758 4128 131764 4140
rect 112496 4100 131764 4128
rect 112496 4088 112502 4100
rect 131758 4088 131764 4100
rect 131816 4088 131822 4140
rect 141418 4088 141424 4140
rect 141476 4128 141482 4140
rect 144730 4128 144736 4140
rect 141476 4100 144736 4128
rect 141476 4088 141482 4100
rect 144730 4088 144736 4100
rect 144788 4088 144794 4140
rect 222838 4088 222844 4140
rect 222896 4128 222902 4140
rect 222896 4100 229094 4128
rect 222896 4088 222902 4100
rect 112806 4060 112812 4072
rect 112364 4032 112812 4060
rect 111705 4023 111763 4029
rect 112806 4020 112812 4032
rect 112864 4020 112870 4072
rect 115198 4020 115204 4072
rect 115256 4060 115262 4072
rect 138842 4060 138848 4072
rect 115256 4032 138848 4060
rect 115256 4020 115262 4032
rect 138842 4020 138848 4032
rect 138900 4020 138906 4072
rect 209774 4020 209780 4072
rect 209832 4060 209838 4072
rect 210970 4060 210976 4072
rect 209832 4032 210976 4060
rect 209832 4020 209838 4032
rect 210970 4020 210976 4032
rect 211028 4020 211034 4072
rect 226334 4020 226340 4072
rect 226392 4060 226398 4072
rect 227530 4060 227536 4072
rect 226392 4032 227536 4060
rect 226392 4020 226398 4032
rect 227530 4020 227536 4032
rect 227588 4020 227594 4072
rect 229066 4060 229094 4100
rect 276014 4088 276020 4140
rect 276072 4128 276078 4140
rect 277118 4128 277124 4140
rect 276072 4100 277124 4128
rect 276072 4088 276078 4100
rect 277118 4088 277124 4100
rect 277176 4088 277182 4140
rect 387058 4088 387064 4140
rect 387116 4128 387122 4140
rect 479334 4128 479340 4140
rect 387116 4100 479340 4128
rect 387116 4088 387122 4100
rect 479334 4088 479340 4100
rect 479392 4088 479398 4140
rect 379974 4060 379980 4072
rect 229066 4032 379980 4060
rect 379974 4020 379980 4032
rect 380032 4020 380038 4072
rect 391198 4020 391204 4072
rect 391256 4060 391262 4072
rect 582190 4060 582196 4072
rect 391256 4032 582196 4060
rect 391256 4020 391262 4032
rect 582190 4020 582196 4032
rect 582248 4020 582254 4072
rect 35986 3952 35992 4004
rect 36044 3992 36050 4004
rect 36044 3964 60136 3992
rect 36044 3952 36050 3964
rect 12342 3884 12348 3936
rect 12400 3924 12406 3936
rect 29638 3924 29644 3936
rect 12400 3896 29644 3924
rect 12400 3884 12406 3896
rect 29638 3884 29644 3896
rect 29696 3884 29702 3936
rect 31294 3884 31300 3936
rect 31352 3924 31358 3936
rect 58897 3927 58955 3933
rect 58897 3924 58909 3927
rect 31352 3896 58909 3924
rect 31352 3884 31358 3896
rect 58897 3893 58909 3896
rect 58943 3893 58955 3927
rect 58897 3887 58955 3893
rect 58989 3927 59047 3933
rect 58989 3893 59001 3927
rect 59035 3924 59047 3927
rect 60001 3927 60059 3933
rect 60001 3924 60013 3927
rect 59035 3896 60013 3924
rect 59035 3893 59047 3896
rect 58989 3887 59047 3893
rect 60001 3893 60013 3896
rect 60047 3893 60059 3927
rect 60001 3887 60059 3893
rect 28810 3816 28816 3868
rect 28868 3856 28874 3868
rect 59909 3859 59967 3865
rect 59909 3856 59921 3859
rect 28868 3828 59921 3856
rect 28868 3816 28874 3828
rect 59909 3825 59921 3828
rect 59955 3825 59967 3859
rect 59909 3819 59967 3825
rect 1670 3748 1676 3800
rect 1728 3788 1734 3800
rect 21358 3788 21364 3800
rect 1728 3760 21364 3788
rect 1728 3748 1734 3760
rect 21358 3748 21364 3760
rect 21416 3748 21422 3800
rect 23014 3748 23020 3800
rect 23072 3788 23078 3800
rect 60108 3788 60136 3964
rect 60826 3952 60832 4004
rect 60884 3992 60890 4004
rect 64233 3995 64291 4001
rect 64233 3992 64245 3995
rect 60884 3964 64245 3992
rect 60884 3952 60890 3964
rect 64233 3961 64245 3964
rect 64279 3961 64291 3995
rect 64233 3955 64291 3961
rect 64322 3952 64328 4004
rect 64380 3952 64386 4004
rect 90910 3952 90916 4004
rect 90968 3992 90974 4004
rect 119890 3992 119896 4004
rect 90968 3964 119896 3992
rect 90968 3952 90974 3964
rect 119890 3952 119896 3964
rect 119948 3952 119954 4004
rect 168098 3952 168104 4004
rect 168156 3992 168162 4004
rect 429654 3992 429660 4004
rect 168156 3964 429660 3992
rect 168156 3952 168162 3964
rect 429654 3952 429660 3964
rect 429712 3952 429718 4004
rect 436830 3952 436836 4004
rect 436888 3992 436894 4004
rect 442626 3992 442632 4004
rect 436888 3964 442632 3992
rect 436888 3952 436894 3964
rect 442626 3952 442632 3964
rect 442684 3952 442690 4004
rect 447778 3952 447784 4004
rect 447836 3992 447842 4004
rect 447836 3964 454632 3992
rect 447836 3952 447842 3964
rect 60185 3927 60243 3933
rect 60185 3893 60197 3927
rect 60231 3924 60243 3927
rect 63678 3924 63684 3936
rect 60231 3896 63684 3924
rect 60231 3893 60243 3896
rect 60185 3887 60243 3893
rect 63678 3884 63684 3896
rect 63736 3884 63742 3936
rect 63770 3884 63776 3936
rect 63828 3924 63834 3936
rect 64340 3924 64368 3952
rect 63828 3896 64368 3924
rect 63828 3884 63834 3896
rect 89622 3884 89628 3936
rect 89680 3924 89686 3936
rect 117590 3924 117596 3936
rect 89680 3896 117596 3924
rect 89680 3884 89686 3896
rect 117590 3884 117596 3896
rect 117648 3884 117654 3936
rect 144178 3884 144184 3936
rect 144236 3924 144242 3936
rect 161290 3924 161296 3936
rect 144236 3896 161296 3924
rect 144236 3884 144242 3896
rect 161290 3884 161296 3896
rect 161348 3884 161354 3936
rect 174538 3884 174544 3936
rect 174596 3924 174602 3936
rect 436738 3924 436744 3936
rect 174596 3896 436744 3924
rect 174596 3884 174602 3896
rect 436738 3884 436744 3896
rect 436796 3884 436802 3936
rect 64322 3816 64328 3868
rect 64380 3856 64386 3868
rect 66990 3856 66996 3868
rect 64380 3828 66996 3856
rect 64380 3816 64386 3828
rect 66990 3816 66996 3828
rect 67048 3816 67054 3868
rect 82538 3816 82544 3868
rect 82596 3856 82602 3868
rect 85666 3856 85672 3868
rect 82596 3828 85672 3856
rect 82596 3816 82602 3828
rect 85666 3816 85672 3828
rect 85724 3816 85730 3868
rect 90726 3816 90732 3868
rect 90784 3856 90790 3868
rect 118786 3856 118792 3868
rect 90784 3828 118792 3856
rect 90784 3816 90790 3828
rect 118786 3816 118792 3828
rect 118844 3816 118850 3868
rect 119338 3816 119344 3868
rect 119396 3856 119402 3868
rect 145926 3856 145932 3868
rect 119396 3828 145932 3856
rect 119396 3816 119402 3828
rect 145926 3816 145932 3828
rect 145984 3816 145990 3868
rect 172146 3816 172152 3868
rect 172204 3856 172210 3868
rect 443822 3856 443828 3868
rect 172204 3828 443828 3856
rect 172204 3816 172210 3828
rect 443822 3816 443828 3828
rect 443880 3816 443886 3868
rect 450538 3816 450544 3868
rect 450596 3856 450602 3868
rect 454604 3856 454632 3964
rect 479518 3952 479524 4004
rect 479576 3992 479582 4004
rect 505370 3992 505376 4004
rect 479576 3964 505376 3992
rect 479576 3952 479582 3964
rect 505370 3952 505376 3964
rect 505428 3952 505434 4004
rect 454678 3884 454684 3936
rect 454736 3924 454742 3936
rect 480530 3924 480536 3936
rect 454736 3896 480536 3924
rect 454736 3884 454742 3896
rect 480530 3884 480536 3896
rect 480588 3884 480594 3936
rect 510062 3856 510068 3868
rect 450596 3828 451274 3856
rect 454604 3828 510068 3856
rect 450596 3816 450602 3828
rect 66898 3788 66904 3800
rect 23072 3760 59124 3788
rect 60108 3760 66904 3788
rect 23072 3748 23078 3760
rect 19426 3680 19432 3732
rect 19484 3720 19490 3732
rect 58989 3723 59047 3729
rect 58989 3720 59001 3723
rect 19484 3692 59001 3720
rect 19484 3680 19490 3692
rect 58989 3689 59001 3692
rect 59035 3689 59047 3723
rect 59096 3720 59124 3760
rect 66898 3748 66904 3760
rect 66956 3748 66962 3800
rect 90818 3748 90824 3800
rect 90876 3788 90882 3800
rect 121086 3788 121092 3800
rect 90876 3760 121092 3788
rect 90876 3748 90882 3760
rect 121086 3748 121092 3760
rect 121144 3748 121150 3800
rect 122098 3748 122104 3800
rect 122156 3788 122162 3800
rect 122156 3760 122834 3788
rect 122156 3748 122162 3760
rect 62942 3720 62948 3732
rect 59096 3692 62948 3720
rect 58989 3683 59047 3689
rect 62942 3680 62948 3692
rect 63000 3680 63006 3732
rect 91002 3680 91008 3732
rect 91060 3720 91066 3732
rect 122282 3720 122288 3732
rect 91060 3692 122288 3720
rect 91060 3680 91066 3692
rect 122282 3680 122288 3692
rect 122340 3680 122346 3732
rect 122806 3720 122834 3760
rect 128998 3748 129004 3800
rect 129056 3788 129062 3800
rect 148318 3788 148324 3800
rect 129056 3760 148324 3788
rect 129056 3748 129062 3760
rect 148318 3748 148324 3760
rect 148376 3748 148382 3800
rect 175918 3748 175924 3800
rect 175976 3788 175982 3800
rect 450906 3788 450912 3800
rect 175976 3760 450912 3788
rect 175976 3748 175982 3760
rect 450906 3748 450912 3760
rect 450964 3748 450970 3800
rect 451246 3788 451274 3828
rect 510062 3816 510068 3828
rect 510120 3816 510126 3868
rect 506474 3788 506480 3800
rect 451246 3760 506480 3788
rect 506474 3748 506480 3760
rect 506532 3748 506538 3800
rect 135254 3720 135260 3732
rect 122806 3692 135260 3720
rect 135254 3680 135260 3692
rect 135312 3680 135318 3732
rect 142798 3680 142804 3732
rect 142856 3720 142862 3732
rect 171962 3720 171968 3732
rect 142856 3692 171968 3720
rect 142856 3680 142862 3692
rect 171962 3680 171968 3692
rect 172020 3680 172026 3732
rect 176562 3680 176568 3732
rect 176620 3720 176626 3732
rect 458082 3720 458088 3732
rect 176620 3692 458088 3720
rect 176620 3680 176626 3692
rect 458082 3680 458088 3692
rect 458140 3680 458146 3732
rect 461670 3680 461676 3732
rect 461728 3720 461734 3732
rect 487614 3720 487620 3732
rect 461728 3692 487620 3720
rect 461728 3680 461734 3692
rect 487614 3680 487620 3692
rect 487672 3680 487678 3732
rect 544378 3680 544384 3732
rect 544436 3720 544442 3732
rect 557350 3720 557356 3732
rect 544436 3692 557356 3720
rect 544436 3680 544442 3692
rect 557350 3680 557356 3692
rect 557408 3680 557414 3732
rect 8754 3612 8760 3664
rect 8812 3652 8818 3664
rect 8812 3624 11100 3652
rect 8812 3612 8818 3624
rect 9950 3544 9956 3596
rect 10008 3584 10014 3596
rect 10962 3584 10968 3596
rect 10008 3556 10968 3584
rect 10008 3544 10014 3556
rect 10962 3544 10968 3556
rect 11020 3544 11026 3596
rect 11072 3584 11100 3624
rect 11146 3612 11152 3664
rect 11204 3652 11210 3664
rect 62482 3652 62488 3664
rect 11204 3624 62488 3652
rect 11204 3612 11210 3624
rect 62482 3612 62488 3624
rect 62540 3612 62546 3664
rect 84010 3612 84016 3664
rect 84068 3652 84074 3664
rect 91554 3652 91560 3664
rect 84068 3624 91560 3652
rect 84068 3612 84074 3624
rect 91554 3612 91560 3624
rect 91612 3612 91618 3664
rect 92382 3612 92388 3664
rect 92440 3652 92446 3664
rect 124674 3652 124680 3664
rect 92440 3624 124680 3652
rect 92440 3612 92446 3624
rect 124674 3612 124680 3624
rect 124732 3612 124738 3664
rect 134518 3612 134524 3664
rect 134576 3652 134582 3664
rect 164878 3652 164884 3664
rect 134576 3624 164884 3652
rect 134576 3612 134582 3624
rect 164878 3612 164884 3624
rect 164936 3612 164942 3664
rect 177942 3612 177948 3664
rect 178000 3652 178006 3664
rect 465166 3652 465172 3664
rect 178000 3624 465172 3652
rect 178000 3612 178006 3624
rect 465166 3612 465172 3624
rect 465224 3612 465230 3664
rect 472618 3612 472624 3664
rect 472676 3652 472682 3664
rect 476485 3655 476543 3661
rect 476485 3652 476497 3655
rect 472676 3624 476497 3652
rect 472676 3612 472682 3624
rect 476485 3621 476497 3624
rect 476531 3621 476543 3655
rect 476485 3615 476543 3621
rect 485038 3612 485044 3664
rect 485096 3652 485102 3664
rect 517146 3652 517152 3664
rect 485096 3624 517152 3652
rect 485096 3612 485102 3624
rect 517146 3612 517152 3624
rect 517204 3612 517210 3664
rect 532510 3652 532516 3664
rect 528526 3624 532516 3652
rect 62114 3584 62120 3596
rect 11072 3556 62120 3584
rect 62114 3544 62120 3556
rect 62172 3544 62178 3596
rect 64138 3584 64144 3596
rect 62224 3556 64144 3584
rect 5258 3476 5264 3528
rect 5316 3516 5322 3528
rect 5316 3488 58112 3516
rect 5316 3476 5322 3488
rect 566 3408 572 3460
rect 624 3448 630 3460
rect 11698 3448 11704 3460
rect 624 3420 11704 3448
rect 624 3408 630 3420
rect 11698 3408 11704 3420
rect 11756 3408 11762 3460
rect 15930 3408 15936 3460
rect 15988 3448 15994 3460
rect 16482 3448 16488 3460
rect 15988 3420 16488 3448
rect 15988 3408 15994 3420
rect 16482 3408 16488 3420
rect 16540 3408 16546 3460
rect 17034 3408 17040 3460
rect 17092 3448 17098 3460
rect 17862 3448 17868 3460
rect 17092 3420 17868 3448
rect 17092 3408 17098 3420
rect 17862 3408 17868 3420
rect 17920 3408 17926 3460
rect 18230 3408 18236 3460
rect 18288 3448 18294 3460
rect 19242 3448 19248 3460
rect 18288 3420 19248 3448
rect 18288 3408 18294 3420
rect 19242 3408 19248 3420
rect 19300 3408 19306 3460
rect 21818 3408 21824 3460
rect 21876 3448 21882 3460
rect 22830 3448 22836 3460
rect 21876 3420 22836 3448
rect 21876 3408 21882 3420
rect 22830 3408 22836 3420
rect 22888 3408 22894 3460
rect 24210 3408 24216 3460
rect 24268 3448 24274 3460
rect 24762 3448 24768 3460
rect 24268 3420 24768 3448
rect 24268 3408 24274 3420
rect 24762 3408 24768 3420
rect 24820 3408 24826 3460
rect 25314 3408 25320 3460
rect 25372 3448 25378 3460
rect 26142 3448 26148 3460
rect 25372 3420 26148 3448
rect 25372 3408 25378 3420
rect 26142 3408 26148 3420
rect 26200 3408 26206 3460
rect 26510 3408 26516 3460
rect 26568 3448 26574 3460
rect 27522 3448 27528 3460
rect 26568 3420 27528 3448
rect 26568 3408 26574 3420
rect 27522 3408 27528 3420
rect 27580 3408 27586 3460
rect 27706 3408 27712 3460
rect 27764 3448 27770 3460
rect 28902 3448 28908 3460
rect 27764 3420 28908 3448
rect 27764 3408 27770 3420
rect 28902 3408 28908 3420
rect 28960 3408 28966 3460
rect 32398 3408 32404 3460
rect 32456 3448 32462 3460
rect 33042 3448 33048 3460
rect 32456 3420 33048 3448
rect 32456 3408 32462 3420
rect 33042 3408 33048 3420
rect 33100 3408 33106 3460
rect 33594 3408 33600 3460
rect 33652 3448 33658 3460
rect 34422 3448 34428 3460
rect 33652 3420 34428 3448
rect 33652 3408 33658 3420
rect 34422 3408 34428 3420
rect 34480 3408 34486 3460
rect 34790 3408 34796 3460
rect 34848 3448 34854 3460
rect 35802 3448 35808 3460
rect 34848 3420 35808 3448
rect 34848 3408 34854 3420
rect 35802 3408 35808 3420
rect 35860 3408 35866 3460
rect 40678 3408 40684 3460
rect 40736 3448 40742 3460
rect 41322 3448 41328 3460
rect 40736 3420 41328 3448
rect 40736 3408 40742 3420
rect 41322 3408 41328 3420
rect 41380 3408 41386 3460
rect 41874 3408 41880 3460
rect 41932 3448 41938 3460
rect 43438 3448 43444 3460
rect 41932 3420 43444 3448
rect 41932 3408 41938 3420
rect 43438 3408 43444 3420
rect 43496 3408 43502 3460
rect 46658 3408 46664 3460
rect 46716 3448 46722 3460
rect 50338 3448 50344 3460
rect 46716 3420 50344 3448
rect 46716 3408 46722 3420
rect 50338 3408 50344 3420
rect 50396 3408 50402 3460
rect 51350 3408 51356 3460
rect 51408 3448 51414 3460
rect 52362 3448 52368 3460
rect 51408 3420 52368 3448
rect 51408 3408 51414 3420
rect 52362 3408 52368 3420
rect 52420 3408 52426 3460
rect 45462 3340 45468 3392
rect 45520 3380 45526 3392
rect 57977 3383 58035 3389
rect 57977 3380 57989 3383
rect 45520 3352 57989 3380
rect 45520 3340 45526 3352
rect 57977 3349 57989 3352
rect 58023 3349 58035 3383
rect 58084 3380 58112 3488
rect 58434 3476 58440 3528
rect 58492 3516 58498 3528
rect 59262 3516 59268 3528
rect 58492 3488 59268 3516
rect 58492 3476 58498 3488
rect 59262 3476 59268 3488
rect 59320 3476 59326 3528
rect 62224 3516 62252 3556
rect 64138 3544 64144 3556
rect 64196 3544 64202 3596
rect 81342 3544 81348 3596
rect 81400 3584 81406 3596
rect 81400 3556 82216 3584
rect 81400 3544 81406 3556
rect 59372 3488 62252 3516
rect 58713 3451 58771 3457
rect 58713 3417 58725 3451
rect 58759 3448 58771 3451
rect 59372 3448 59400 3488
rect 63218 3476 63224 3528
rect 63276 3516 63282 3528
rect 74718 3516 74724 3528
rect 63276 3488 74724 3516
rect 63276 3476 63282 3488
rect 74718 3476 74724 3488
rect 74776 3476 74782 3528
rect 74994 3476 75000 3528
rect 75052 3516 75058 3528
rect 75822 3516 75828 3528
rect 75052 3488 75828 3516
rect 75052 3476 75058 3488
rect 75822 3476 75828 3488
rect 75880 3476 75886 3528
rect 76190 3476 76196 3528
rect 76248 3516 76254 3528
rect 77202 3516 77208 3528
rect 76248 3488 77208 3516
rect 76248 3476 76254 3488
rect 77202 3476 77208 3488
rect 77260 3476 77266 3528
rect 80330 3476 80336 3528
rect 80388 3516 80394 3528
rect 80882 3516 80888 3528
rect 80388 3488 80888 3516
rect 80388 3476 80394 3488
rect 80882 3476 80888 3488
rect 80940 3476 80946 3528
rect 81250 3476 81256 3528
rect 81308 3516 81314 3528
rect 82078 3516 82084 3528
rect 81308 3488 82084 3516
rect 81308 3476 81314 3488
rect 82078 3476 82084 3488
rect 82136 3476 82142 3528
rect 82188 3516 82216 3556
rect 83458 3544 83464 3596
rect 83516 3584 83522 3596
rect 87966 3584 87972 3596
rect 83516 3556 87972 3584
rect 83516 3544 83522 3556
rect 87966 3544 87972 3556
rect 88024 3544 88030 3596
rect 90634 3544 90640 3596
rect 90692 3584 90698 3596
rect 123478 3584 123484 3596
rect 90692 3556 123484 3584
rect 90692 3544 90698 3556
rect 123478 3544 123484 3556
rect 123536 3544 123542 3596
rect 124858 3544 124864 3596
rect 124916 3584 124922 3596
rect 125870 3584 125876 3596
rect 124916 3556 125876 3584
rect 124916 3544 124922 3556
rect 125870 3544 125876 3556
rect 125928 3544 125934 3596
rect 137278 3544 137284 3596
rect 137336 3584 137342 3596
rect 168374 3584 168380 3596
rect 137336 3556 168380 3584
rect 137336 3544 137342 3556
rect 168374 3544 168380 3556
rect 168432 3544 168438 3596
rect 179322 3544 179328 3596
rect 179380 3584 179386 3596
rect 472250 3584 472256 3596
rect 179380 3556 472256 3584
rect 179380 3544 179386 3556
rect 472250 3544 472256 3556
rect 472308 3544 472314 3596
rect 473354 3544 473360 3596
rect 473412 3584 473418 3596
rect 474550 3584 474556 3596
rect 473412 3556 474556 3584
rect 473412 3544 473418 3556
rect 474550 3544 474556 3556
rect 474608 3544 474614 3596
rect 481634 3544 481640 3596
rect 481692 3584 481698 3596
rect 482830 3584 482836 3596
rect 481692 3556 482836 3584
rect 481692 3544 481698 3556
rect 482830 3544 482836 3556
rect 482888 3544 482894 3596
rect 489178 3544 489184 3596
rect 489236 3584 489242 3596
rect 528526 3584 528554 3624
rect 532510 3612 532516 3624
rect 532568 3612 532574 3664
rect 537478 3612 537484 3664
rect 537536 3652 537542 3664
rect 553762 3652 553768 3664
rect 537536 3624 553768 3652
rect 537536 3612 537542 3624
rect 553762 3612 553768 3624
rect 553820 3612 553826 3664
rect 489236 3556 528554 3584
rect 489236 3544 489242 3556
rect 530578 3544 530584 3596
rect 530636 3584 530642 3596
rect 531314 3584 531320 3596
rect 530636 3556 531320 3584
rect 530636 3544 530642 3556
rect 531314 3544 531320 3556
rect 531372 3544 531378 3596
rect 533338 3544 533344 3596
rect 533396 3584 533402 3596
rect 550266 3584 550272 3596
rect 533396 3556 550272 3584
rect 533396 3544 533402 3556
rect 550266 3544 550272 3556
rect 550324 3544 550330 3596
rect 572714 3544 572720 3596
rect 572772 3584 572778 3596
rect 573910 3584 573916 3596
rect 572772 3556 573916 3584
rect 572772 3544 572778 3556
rect 573910 3544 573916 3556
rect 573968 3544 573974 3596
rect 84470 3516 84476 3528
rect 82188 3488 84476 3516
rect 84470 3476 84476 3488
rect 84528 3476 84534 3528
rect 85482 3476 85488 3528
rect 85540 3516 85546 3528
rect 85540 3488 89300 3516
rect 85540 3476 85546 3488
rect 58759 3420 59400 3448
rect 59909 3451 59967 3457
rect 58759 3417 58771 3420
rect 58713 3411 58771 3417
rect 59909 3417 59921 3451
rect 59955 3448 59967 3451
rect 66438 3448 66444 3460
rect 59955 3420 66444 3448
rect 59955 3417 59967 3420
rect 59909 3411 59967 3417
rect 66438 3408 66444 3420
rect 66496 3408 66502 3460
rect 66714 3408 66720 3460
rect 66772 3448 66778 3460
rect 67542 3448 67548 3460
rect 66772 3420 67548 3448
rect 66772 3408 66778 3420
rect 67542 3408 67548 3420
rect 67600 3408 67606 3460
rect 67910 3408 67916 3460
rect 67968 3448 67974 3460
rect 68922 3448 68928 3460
rect 67968 3420 68928 3448
rect 67968 3408 67974 3420
rect 68922 3408 68928 3420
rect 68980 3408 68986 3460
rect 69106 3408 69112 3460
rect 69164 3448 69170 3460
rect 70210 3448 70216 3460
rect 69164 3420 70216 3448
rect 69164 3408 69170 3420
rect 70210 3408 70216 3420
rect 70268 3408 70274 3460
rect 72602 3408 72608 3460
rect 72660 3448 72666 3460
rect 73062 3448 73068 3460
rect 72660 3420 73068 3448
rect 72660 3408 72666 3420
rect 73062 3408 73068 3420
rect 73120 3408 73126 3460
rect 73798 3408 73804 3460
rect 73856 3448 73862 3460
rect 75178 3448 75184 3460
rect 73856 3420 75184 3448
rect 73856 3408 73862 3420
rect 75178 3408 75184 3420
rect 75236 3408 75242 3460
rect 77386 3408 77392 3460
rect 77444 3448 77450 3460
rect 78950 3448 78956 3460
rect 77444 3420 78956 3448
rect 77444 3408 77450 3420
rect 78950 3408 78956 3420
rect 79008 3408 79014 3460
rect 79686 3408 79692 3460
rect 79744 3448 79750 3460
rect 80422 3448 80428 3460
rect 79744 3420 80428 3448
rect 79744 3408 79750 3420
rect 80422 3408 80428 3420
rect 80480 3408 80486 3460
rect 82630 3408 82636 3460
rect 82688 3448 82694 3460
rect 89162 3448 89168 3460
rect 82688 3420 89168 3448
rect 82688 3408 82694 3420
rect 89162 3408 89168 3420
rect 89220 3408 89226 3460
rect 89272 3448 89300 3488
rect 89346 3476 89352 3528
rect 89404 3516 89410 3528
rect 116394 3516 116400 3528
rect 89404 3488 116400 3516
rect 89404 3476 89410 3488
rect 116394 3476 116400 3488
rect 116452 3476 116458 3528
rect 116578 3476 116584 3528
rect 116636 3516 116642 3528
rect 153010 3516 153016 3528
rect 116636 3488 153016 3516
rect 116636 3476 116642 3488
rect 153010 3476 153016 3488
rect 153068 3476 153074 3528
rect 193214 3476 193220 3528
rect 193272 3516 193278 3528
rect 194410 3516 194416 3528
rect 193272 3488 194416 3516
rect 193272 3476 193278 3488
rect 194410 3476 194416 3488
rect 194468 3476 194474 3528
rect 206922 3476 206928 3528
rect 206980 3516 206986 3528
rect 580994 3516 581000 3528
rect 206980 3488 581000 3516
rect 206980 3476 206986 3488
rect 580994 3476 581000 3488
rect 581052 3476 581058 3528
rect 99834 3448 99840 3460
rect 89272 3420 99840 3448
rect 99834 3408 99840 3420
rect 99892 3408 99898 3460
rect 100386 3408 100392 3460
rect 100444 3448 100450 3460
rect 100444 3420 142154 3448
rect 100444 3408 100450 3420
rect 61010 3380 61016 3392
rect 58084 3352 61016 3380
rect 57977 3343 58035 3349
rect 61010 3340 61016 3352
rect 61068 3340 61074 3392
rect 65518 3340 65524 3392
rect 65576 3380 65582 3392
rect 76098 3380 76104 3392
rect 65576 3352 76104 3380
rect 65576 3340 65582 3352
rect 76098 3340 76104 3352
rect 76156 3340 76162 3392
rect 88242 3340 88248 3392
rect 88300 3380 88306 3392
rect 109310 3380 109316 3392
rect 88300 3352 109316 3380
rect 88300 3340 88306 3352
rect 109310 3340 109316 3352
rect 109368 3340 109374 3392
rect 142126 3380 142154 3420
rect 147122 3408 147128 3460
rect 147180 3448 147186 3460
rect 149514 3448 149520 3460
rect 147180 3420 149520 3448
rect 147180 3408 147186 3420
rect 149514 3408 149520 3420
rect 149572 3408 149578 3460
rect 152458 3408 152464 3460
rect 152516 3448 152522 3460
rect 156598 3448 156604 3460
rect 152516 3420 156604 3448
rect 152516 3408 152522 3420
rect 156598 3408 156604 3420
rect 156656 3408 156662 3460
rect 206830 3408 206836 3460
rect 206888 3448 206894 3460
rect 583386 3448 583392 3460
rect 206888 3420 583392 3448
rect 206888 3408 206894 3420
rect 583386 3408 583392 3420
rect 583444 3408 583450 3460
rect 160094 3380 160100 3392
rect 142126 3352 160100 3380
rect 160094 3340 160100 3352
rect 160152 3340 160158 3392
rect 242894 3340 242900 3392
rect 242952 3380 242958 3392
rect 244090 3380 244096 3392
rect 242952 3352 244096 3380
rect 242952 3340 242958 3352
rect 244090 3340 244096 3352
rect 244148 3340 244154 3392
rect 307754 3340 307760 3392
rect 307812 3380 307818 3392
rect 309042 3380 309048 3392
rect 307812 3352 309048 3380
rect 307812 3340 307818 3352
rect 309042 3340 309048 3352
rect 309100 3340 309106 3392
rect 316034 3340 316040 3392
rect 316092 3380 316098 3392
rect 317322 3380 317328 3392
rect 316092 3352 317328 3380
rect 316092 3340 316098 3352
rect 317322 3340 317328 3352
rect 317380 3340 317386 3392
rect 332594 3340 332600 3392
rect 332652 3380 332658 3392
rect 333882 3380 333888 3392
rect 332652 3352 333888 3380
rect 332652 3340 332658 3352
rect 333882 3340 333888 3352
rect 333940 3340 333946 3392
rect 349154 3340 349160 3392
rect 349212 3380 349218 3392
rect 350442 3380 350448 3392
rect 349212 3352 350448 3380
rect 349212 3340 349218 3352
rect 350442 3340 350448 3352
rect 350500 3340 350506 3392
rect 373994 3340 374000 3392
rect 374052 3380 374058 3392
rect 375282 3380 375288 3392
rect 374052 3352 375288 3380
rect 374052 3340 374058 3352
rect 375282 3340 375288 3352
rect 375340 3340 375346 3392
rect 382918 3340 382924 3392
rect 382976 3380 382982 3392
rect 475746 3380 475752 3392
rect 382976 3352 475752 3380
rect 382976 3340 382982 3352
rect 475746 3340 475752 3352
rect 475804 3340 475810 3392
rect 498194 3380 498200 3392
rect 475856 3352 498200 3380
rect 44266 3272 44272 3324
rect 44324 3312 44330 3324
rect 58897 3315 58955 3321
rect 44324 3284 58848 3312
rect 44324 3272 44330 3284
rect 50154 3204 50160 3256
rect 50212 3244 50218 3256
rect 58713 3247 58771 3253
rect 58713 3244 58725 3247
rect 50212 3216 58725 3244
rect 50212 3204 50218 3216
rect 58713 3213 58725 3216
rect 58759 3213 58771 3247
rect 58820 3244 58848 3284
rect 58897 3281 58909 3315
rect 58943 3312 58955 3315
rect 64414 3312 64420 3324
rect 58943 3284 64420 3312
rect 58943 3281 58955 3284
rect 58897 3275 58955 3281
rect 64414 3272 64420 3284
rect 64472 3272 64478 3324
rect 86678 3272 86684 3324
rect 86736 3312 86742 3324
rect 105722 3312 105728 3324
rect 86736 3284 105728 3312
rect 86736 3272 86742 3284
rect 105722 3272 105728 3284
rect 105780 3272 105786 3324
rect 106918 3272 106924 3324
rect 106976 3312 106982 3324
rect 111610 3312 111616 3324
rect 106976 3284 111616 3312
rect 106976 3272 106982 3284
rect 111610 3272 111616 3284
rect 111668 3272 111674 3324
rect 111705 3315 111763 3321
rect 111705 3281 111717 3315
rect 111751 3312 111763 3315
rect 115198 3312 115204 3324
rect 111751 3284 115204 3312
rect 111751 3281 111763 3284
rect 111705 3275 111763 3281
rect 115198 3272 115204 3284
rect 115256 3272 115262 3324
rect 382274 3272 382280 3324
rect 382332 3312 382338 3324
rect 383562 3312 383568 3324
rect 382332 3284 383568 3312
rect 382332 3272 382338 3284
rect 383562 3272 383568 3284
rect 383620 3272 383626 3324
rect 398834 3272 398840 3324
rect 398892 3312 398898 3324
rect 400122 3312 400128 3324
rect 398892 3284 400128 3312
rect 398892 3272 398898 3284
rect 400122 3272 400128 3284
rect 400180 3272 400186 3324
rect 407758 3272 407764 3324
rect 407816 3312 407822 3324
rect 409598 3312 409604 3324
rect 407816 3284 409604 3312
rect 407816 3272 407822 3284
rect 409598 3272 409604 3284
rect 409656 3272 409662 3324
rect 414658 3272 414664 3324
rect 414716 3312 414722 3324
rect 416682 3312 416688 3324
rect 414716 3284 416688 3312
rect 414716 3272 414722 3284
rect 416682 3272 416688 3284
rect 416740 3272 416746 3324
rect 423766 3272 423772 3324
rect 423824 3312 423830 3324
rect 424962 3312 424968 3324
rect 423824 3284 424968 3312
rect 423824 3272 423830 3284
rect 424962 3272 424968 3284
rect 425020 3272 425026 3324
rect 475378 3272 475384 3324
rect 475436 3312 475442 3324
rect 475856 3312 475884 3352
rect 498194 3340 498200 3352
rect 498252 3340 498258 3392
rect 512638 3340 512644 3392
rect 512696 3380 512702 3392
rect 513558 3380 513564 3392
rect 512696 3352 513564 3380
rect 512696 3340 512702 3352
rect 513558 3340 513564 3352
rect 513616 3340 513622 3392
rect 526438 3340 526444 3392
rect 526496 3380 526502 3392
rect 527818 3380 527824 3392
rect 526496 3352 527824 3380
rect 526496 3340 526502 3352
rect 527818 3340 527824 3352
rect 527876 3340 527882 3392
rect 547874 3340 547880 3392
rect 547932 3380 547938 3392
rect 549070 3380 549076 3392
rect 547932 3352 549076 3380
rect 547932 3340 547938 3352
rect 549070 3340 549076 3352
rect 549128 3340 549134 3392
rect 475436 3284 475884 3312
rect 476485 3315 476543 3321
rect 475436 3272 475442 3284
rect 476485 3281 476497 3315
rect 476531 3312 476543 3315
rect 494698 3312 494704 3324
rect 476531 3284 494704 3312
rect 476531 3281 476543 3284
rect 476485 3275 476543 3281
rect 494698 3272 494704 3284
rect 494756 3272 494762 3324
rect 62850 3244 62856 3256
rect 58820 3216 62856 3244
rect 58713 3207 58771 3213
rect 62850 3204 62856 3216
rect 62908 3204 62914 3256
rect 86770 3204 86776 3256
rect 86828 3244 86834 3256
rect 102226 3244 102232 3256
rect 86828 3216 102232 3244
rect 86828 3204 86834 3216
rect 102226 3204 102232 3216
rect 102284 3204 102290 3256
rect 102870 3204 102876 3256
rect 102928 3244 102934 3256
rect 114002 3244 114008 3256
rect 102928 3216 114008 3244
rect 102928 3204 102934 3216
rect 114002 3204 114008 3216
rect 114060 3204 114066 3256
rect 388438 3204 388444 3256
rect 388496 3244 388502 3256
rect 390646 3244 390652 3256
rect 388496 3216 390652 3244
rect 388496 3204 388502 3216
rect 390646 3204 390652 3216
rect 390704 3204 390710 3256
rect 407114 3204 407120 3256
rect 407172 3244 407178 3256
rect 408402 3244 408408 3256
rect 407172 3216 408408 3244
rect 407172 3204 407178 3216
rect 408402 3204 408408 3216
rect 408460 3204 408466 3256
rect 418798 3204 418804 3256
rect 418856 3244 418862 3256
rect 420178 3244 420184 3256
rect 418856 3216 420184 3244
rect 418856 3204 418862 3216
rect 420178 3204 420184 3216
rect 420236 3204 420242 3256
rect 468478 3204 468484 3256
rect 468536 3244 468542 3256
rect 491110 3244 491116 3256
rect 468536 3216 491116 3244
rect 468536 3204 468542 3216
rect 491110 3204 491116 3216
rect 491168 3204 491174 3256
rect 519630 3204 519636 3256
rect 519688 3244 519694 3256
rect 524230 3244 524236 3256
rect 519688 3216 524236 3244
rect 519688 3204 519694 3216
rect 524230 3204 524236 3216
rect 524288 3204 524294 3256
rect 56042 3136 56048 3188
rect 56100 3176 56106 3188
rect 68278 3176 68284 3188
rect 56100 3148 68284 3176
rect 56100 3136 56106 3148
rect 68278 3136 68284 3148
rect 68336 3136 68342 3188
rect 87598 3136 87604 3188
rect 87656 3176 87662 3188
rect 98638 3176 98644 3188
rect 87656 3148 98644 3176
rect 87656 3136 87662 3148
rect 98638 3136 98644 3148
rect 98696 3136 98702 3188
rect 102778 3136 102784 3188
rect 102836 3176 102842 3188
rect 110506 3176 110512 3188
rect 102836 3148 110512 3176
rect 102836 3136 102842 3148
rect 110506 3136 110512 3148
rect 110564 3136 110570 3188
rect 396718 3136 396724 3188
rect 396776 3176 396782 3188
rect 397730 3176 397736 3188
rect 396776 3148 397736 3176
rect 396776 3136 396782 3148
rect 397730 3136 397736 3148
rect 397788 3136 397794 3188
rect 443638 3136 443644 3188
rect 443696 3176 443702 3188
rect 449802 3176 449808 3188
rect 443696 3148 449808 3176
rect 443696 3136 443702 3148
rect 449802 3136 449808 3148
rect 449860 3136 449866 3188
rect 52546 3068 52552 3120
rect 52604 3108 52610 3120
rect 62758 3108 62764 3120
rect 52604 3080 62764 3108
rect 52604 3068 52610 3080
rect 62758 3068 62764 3080
rect 62816 3068 62822 3120
rect 86862 3068 86868 3120
rect 86920 3108 86926 3120
rect 103330 3108 103336 3120
rect 86920 3080 103336 3108
rect 86920 3068 86926 3080
rect 103330 3068 103336 3080
rect 103388 3068 103394 3120
rect 2866 3000 2872 3052
rect 2924 3040 2930 3052
rect 4798 3040 4804 3052
rect 2924 3012 4804 3040
rect 2924 3000 2930 3012
rect 4798 3000 4804 3012
rect 4856 3000 4862 3052
rect 48958 3000 48964 3052
rect 49016 3040 49022 3052
rect 57146 3040 57152 3052
rect 49016 3012 57152 3040
rect 49016 3000 49022 3012
rect 57146 3000 57152 3012
rect 57204 3000 57210 3052
rect 57238 3000 57244 3052
rect 57296 3040 57302 3052
rect 65610 3040 65616 3052
rect 57296 3012 65616 3040
rect 57296 3000 57302 3012
rect 65610 3000 65616 3012
rect 65668 3000 65674 3052
rect 84102 3000 84108 3052
rect 84160 3040 84166 3052
rect 95142 3040 95148 3052
rect 84160 3012 95148 3040
rect 84160 3000 84166 3012
rect 95142 3000 95148 3012
rect 95200 3000 95206 3052
rect 101398 3000 101404 3052
rect 101456 3040 101462 3052
rect 106918 3040 106924 3052
rect 101456 3012 106924 3040
rect 101456 3000 101462 3012
rect 106918 3000 106924 3012
rect 106976 3000 106982 3052
rect 425790 3000 425796 3052
rect 425848 3040 425854 3052
rect 427262 3040 427268 3052
rect 425848 3012 427268 3040
rect 425848 3000 425854 3012
rect 427262 3000 427268 3012
rect 427320 3000 427326 3052
rect 59630 2932 59636 2984
rect 59688 2972 59694 2984
rect 68370 2972 68376 2984
rect 59688 2944 68376 2972
rect 59688 2932 59694 2944
rect 68370 2932 68376 2944
rect 68428 2932 68434 2984
rect 86218 2932 86224 2984
rect 86276 2972 86282 2984
rect 96246 2972 96252 2984
rect 86276 2944 96252 2972
rect 86276 2932 86282 2944
rect 96246 2932 96252 2944
rect 96304 2932 96310 2984
rect 7650 2864 7656 2916
rect 7708 2904 7714 2916
rect 8202 2904 8208 2916
rect 7708 2876 8208 2904
rect 7708 2864 7714 2876
rect 8202 2864 8208 2876
rect 8260 2864 8266 2916
rect 57977 2907 58035 2913
rect 57977 2873 57989 2907
rect 58023 2904 58035 2907
rect 63770 2904 63776 2916
rect 58023 2876 63776 2904
rect 58023 2873 58035 2876
rect 57977 2867 58035 2873
rect 63770 2864 63776 2876
rect 63828 2864 63834 2916
rect 82722 2864 82728 2916
rect 82780 2904 82786 2916
rect 86862 2904 86868 2916
rect 82780 2876 86868 2904
rect 82780 2864 82786 2876
rect 86862 2864 86868 2876
rect 86920 2864 86926 2916
rect 421558 2864 421564 2916
rect 421616 2904 421622 2916
rect 423766 2904 423772 2916
rect 421616 2876 423772 2904
rect 421616 2864 421622 2876
rect 423766 2864 423772 2876
rect 423824 2864 423830 2916
rect 20622 2796 20628 2848
rect 20680 2836 20686 2848
rect 65058 2836 65064 2848
rect 20680 2808 65064 2836
rect 20680 2796 20686 2808
rect 65058 2796 65064 2808
rect 65116 2796 65122 2848
rect 83918 2796 83924 2848
rect 83976 2836 83982 2848
rect 92750 2836 92756 2848
rect 83976 2808 92756 2836
rect 83976 2796 83982 2808
rect 92750 2796 92756 2808
rect 92808 2796 92814 2848
rect 299474 1640 299480 1692
rect 299532 1680 299538 1692
rect 300762 1680 300768 1692
rect 299532 1652 300768 1680
rect 299532 1640 299538 1652
rect 300762 1640 300768 1652
rect 300820 1640 300826 1692
<< via1 >>
rect 201500 702992 201552 703044
rect 202788 702992 202840 703044
rect 204904 700680 204956 700732
rect 235172 700680 235224 700732
rect 206376 700612 206428 700664
rect 267648 700612 267700 700664
rect 213276 700544 213328 700596
rect 283840 700544 283892 700596
rect 377404 700544 377456 700596
rect 397460 700544 397512 700596
rect 446404 700544 446456 700596
rect 494796 700544 494848 700596
rect 198004 700476 198056 700528
rect 300124 700476 300176 700528
rect 376024 700476 376076 700528
rect 462320 700476 462372 700528
rect 215944 700408 215996 700460
rect 332508 700408 332560 700460
rect 388444 700408 388496 700460
rect 478512 700408 478564 700460
rect 40500 700340 40552 700392
rect 41328 700340 41380 700392
rect 170312 700340 170364 700392
rect 196532 700340 196584 700392
rect 209044 700340 209096 700392
rect 348792 700340 348844 700392
rect 374644 700340 374696 700392
rect 527180 700340 527232 700392
rect 24308 700272 24360 700324
rect 33784 700272 33836 700324
rect 59268 700272 59320 700324
rect 72976 700272 73028 700324
rect 154120 700272 154172 700324
rect 196624 700272 196676 700324
rect 214564 700272 214616 700324
rect 559656 700272 559708 700324
rect 88340 699660 88392 699712
rect 89168 699660 89220 699712
rect 104900 699660 104952 699712
rect 105452 699660 105504 699712
rect 214656 699660 214708 699712
rect 218980 699660 219032 699712
rect 360844 699660 360896 699712
rect 364984 699660 365036 699712
rect 371884 696940 371936 696992
rect 580172 696940 580224 696992
rect 138020 696872 138072 696924
rect 140044 696872 140096 696924
rect 140044 689596 140096 689648
rect 141148 689596 141200 689648
rect 141148 683612 141200 683664
rect 143540 683612 143592 683664
rect 3424 683136 3476 683188
rect 11704 683136 11756 683188
rect 385684 683136 385736 683188
rect 580172 683136 580224 683188
rect 143540 680484 143592 680536
rect 145564 680484 145616 680536
rect 3516 670692 3568 670744
rect 36544 670692 36596 670744
rect 213368 670692 213420 670744
rect 580172 670692 580224 670744
rect 145564 663212 145616 663264
rect 149704 663212 149756 663264
rect 3424 656888 3476 656940
rect 22744 656888 22796 656940
rect 149704 645872 149756 645924
rect 153200 645804 153252 645856
rect 370504 643084 370556 643136
rect 580172 643084 580224 643136
rect 153200 638868 153252 638920
rect 155224 638868 155276 638920
rect 3424 632068 3476 632120
rect 14464 632068 14516 632120
rect 382924 630640 382976 630692
rect 580172 630640 580224 630692
rect 155224 627920 155276 627972
rect 160468 627852 160520 627904
rect 160468 619624 160520 619676
rect 163504 619556 163556 619608
rect 3148 618264 3200 618316
rect 35164 618264 35216 618316
rect 209136 616836 209188 616888
rect 580172 616836 580224 616888
rect 163504 611940 163556 611992
rect 164884 611940 164936 611992
rect 3240 605820 3292 605872
rect 25504 605820 25556 605872
rect 367744 590656 367796 590708
rect 579804 590656 579856 590708
rect 164884 585692 164936 585744
rect 167552 585692 167604 585744
rect 3332 579640 3384 579692
rect 21364 579640 21416 579692
rect 167552 579572 167604 579624
rect 170404 579572 170456 579624
rect 449164 576852 449216 576904
rect 580172 576852 580224 576904
rect 170404 569100 170456 569152
rect 172428 569100 172480 569152
rect 3424 565836 3476 565888
rect 39304 565836 39356 565888
rect 172428 563048 172480 563100
rect 206284 563048 206336 563100
rect 579804 563048 579856 563100
rect 178040 562980 178092 563032
rect 178040 560192 178092 560244
rect 180708 560192 180760 560244
rect 3424 553392 3476 553444
rect 29644 553392 29696 553444
rect 180708 552032 180760 552084
rect 182824 551964 182876 552016
rect 182824 542308 182876 542360
rect 184204 542308 184256 542360
rect 431224 536800 431276 536852
rect 580172 536800 580224 536852
rect 184204 534080 184256 534132
rect 186136 534080 186188 534132
rect 186136 531292 186188 531344
rect 187700 531224 187752 531276
rect 187700 529184 187752 529236
rect 196808 529184 196860 529236
rect 3424 527144 3476 527196
rect 15844 527144 15896 527196
rect 381544 524424 381596 524476
rect 580172 524424 580224 524476
rect 3424 514768 3476 514820
rect 43444 514768 43496 514820
rect 204996 510620 205048 510672
rect 580172 510620 580224 510672
rect 89628 505724 89680 505776
rect 218888 505724 218940 505776
rect 114468 505656 114520 505708
rect 218704 505656 218756 505708
rect 144828 505588 144880 505640
rect 216312 505588 216364 505640
rect 142068 505520 142120 505572
rect 216128 505520 216180 505572
rect 143356 505452 143408 505504
rect 216496 505452 216548 505504
rect 219808 505452 219860 505504
rect 260840 505452 260892 505504
rect 133788 505384 133840 505436
rect 218796 505384 218848 505436
rect 219164 505384 219216 505436
rect 288440 505384 288492 505436
rect 129648 505316 129700 505368
rect 219256 505316 219308 505368
rect 219348 505316 219400 505368
rect 298100 505316 298152 505368
rect 117228 505248 117280 505300
rect 219072 505248 219124 505300
rect 219716 505248 219768 505300
rect 300860 505248 300912 505300
rect 217784 505180 217836 505232
rect 316040 505180 316092 505232
rect 218612 505112 218664 505164
rect 325700 505112 325752 505164
rect 56508 505044 56560 505096
rect 153200 505044 153252 505096
rect 158628 505044 158680 505096
rect 219992 505044 220044 505096
rect 57612 504976 57664 505028
rect 317420 504976 317472 505028
rect 53288 504908 53340 504960
rect 128636 504908 128688 504960
rect 58348 504840 58400 504892
rect 104900 504840 104952 504892
rect 108948 504840 109000 504892
rect 148508 504908 148560 504960
rect 164056 504908 164108 504960
rect 218980 504908 219032 504960
rect 219624 504908 219676 504960
rect 273260 504908 273312 504960
rect 197452 504840 197504 504892
rect 219440 504840 219492 504892
rect 277308 504840 277360 504892
rect 146576 504772 146628 504824
rect 215760 504772 215812 504824
rect 218428 504772 218480 504824
rect 277400 504772 277452 504824
rect 55036 504704 55088 504756
rect 149520 504704 149572 504756
rect 215300 504704 215352 504756
rect 219532 504704 219584 504756
rect 280160 504704 280212 504756
rect 98552 504636 98604 504688
rect 197360 504636 197412 504688
rect 218336 504636 218388 504688
rect 282920 504636 282972 504688
rect 57520 504568 57572 504620
rect 156052 504568 156104 504620
rect 219900 504568 219952 504620
rect 111708 504500 111760 504552
rect 215576 504500 215628 504552
rect 218520 504500 218572 504552
rect 295340 504500 295392 504552
rect 56416 504432 56468 504484
rect 165620 504432 165672 504484
rect 212448 504432 212500 504484
rect 307760 504432 307812 504484
rect 60004 504364 60056 504416
rect 88340 504364 88392 504416
rect 103888 504364 103940 504416
rect 215484 504364 215536 504416
rect 216588 504364 216640 504416
rect 313280 504364 313332 504416
rect 101312 504296 101364 504348
rect 215852 504296 215904 504348
rect 216404 504296 216456 504348
rect 320180 504296 320232 504348
rect 96528 504228 96580 504280
rect 215668 504228 215720 504280
rect 216220 504228 216272 504280
rect 322940 504228 322992 504280
rect 52276 504160 52328 504212
rect 176844 504160 176896 504212
rect 206468 504160 206520 504212
rect 339500 504160 339552 504212
rect 57796 504092 57848 504144
rect 270500 504092 270552 504144
rect 50804 504024 50856 504076
rect 265716 504024 265768 504076
rect 52184 503956 52236 504008
rect 267740 503956 267792 504008
rect 50620 503888 50672 503940
rect 302240 503888 302292 503940
rect 53196 503820 53248 503872
rect 305000 503820 305052 503872
rect 55128 503752 55180 503804
rect 310520 503752 310572 503804
rect 53380 503684 53432 503736
rect 129740 503684 129792 503736
rect 160100 503684 160152 503736
rect 180708 503684 180760 503736
rect 216036 503684 216088 503736
rect 218244 503684 218296 503736
rect 292580 503684 292632 503736
rect 53472 503616 53524 503668
rect 123760 503616 123812 503668
rect 220728 503616 220780 503668
rect 245844 503616 245896 503668
rect 53656 503548 53708 503600
rect 104072 503548 104124 503600
rect 93768 503480 93820 503532
rect 123576 503480 123628 503532
rect 201592 503548 201644 503600
rect 53564 503412 53616 503464
rect 113548 503412 113600 503464
rect 121368 503412 121420 503464
rect 200212 503480 200264 503532
rect 200764 503480 200816 503532
rect 263600 503548 263652 503600
rect 218152 503480 218204 503532
rect 285680 503480 285732 503532
rect 339408 503480 339460 503532
rect 356520 503480 356572 503532
rect 191748 503412 191800 503464
rect 218060 503412 218112 503464
rect 286876 503412 286928 503464
rect 350540 503412 350592 503464
rect 213184 503344 213236 503396
rect 196716 503276 196768 503328
rect 213184 502324 213236 502376
rect 2780 501032 2832 501084
rect 4804 501032 4856 501084
rect 196716 487339 196768 487348
rect 196716 487305 196725 487339
rect 196725 487305 196759 487339
rect 196759 487305 196768 487339
rect 196716 487296 196768 487305
rect 219808 486412 219860 486464
rect 196716 486344 196768 486396
rect 196716 486140 196768 486192
rect 363604 484372 363656 484424
rect 580172 484372 580224 484424
rect 196716 483871 196768 483880
rect 196716 483837 196725 483871
rect 196725 483837 196759 483871
rect 196759 483837 196768 483871
rect 196716 483828 196768 483837
rect 219808 483352 219860 483404
rect 219808 483259 219860 483268
rect 219808 483225 219817 483259
rect 219817 483225 219851 483259
rect 219851 483225 219860 483259
rect 219808 483216 219860 483225
rect 219808 481380 219860 481432
rect 219808 480700 219860 480752
rect 3424 474716 3476 474768
rect 17224 474716 17276 474768
rect 219808 470679 219860 470688
rect 219808 470645 219817 470679
rect 219817 470645 219851 470679
rect 219851 470645 219860 470679
rect 219808 470636 219860 470645
rect 443644 470568 443696 470620
rect 579988 470568 580040 470620
rect 219808 470543 219860 470552
rect 219808 470509 219817 470543
rect 219817 470509 219851 470543
rect 219851 470509 219860 470543
rect 219808 470500 219860 470509
rect 3240 462340 3292 462392
rect 47584 462340 47636 462392
rect 358084 456764 358136 456816
rect 580172 456764 580224 456816
rect 219808 451367 219860 451376
rect 219808 451333 219817 451367
rect 219817 451333 219851 451367
rect 219851 451333 219860 451367
rect 219808 451324 219860 451333
rect 219808 451231 219860 451240
rect 219808 451197 219817 451231
rect 219817 451197 219851 451231
rect 219851 451197 219860 451231
rect 219808 451188 219860 451197
rect 3148 448536 3200 448588
rect 32404 448536 32456 448588
rect 219808 432055 219860 432064
rect 219808 432021 219817 432055
rect 219817 432021 219851 432055
rect 219851 432021 219860 432055
rect 219808 432012 219860 432021
rect 219808 431919 219860 431928
rect 219808 431885 219817 431919
rect 219817 431885 219851 431919
rect 219851 431885 219860 431919
rect 219808 431876 219860 431885
rect 210516 430584 210568 430636
rect 216680 430584 216732 430636
rect 378784 430584 378836 430636
rect 580172 430584 580224 430636
rect 50712 429156 50764 429208
rect 57336 429156 57388 429208
rect 210608 429156 210660 429208
rect 216680 429156 216732 429208
rect 57336 426640 57388 426692
rect 57888 426640 57940 426692
rect 219808 422356 219860 422408
rect 3424 422288 3476 422340
rect 18604 422288 18656 422340
rect 219808 422220 219860 422272
rect 219808 412743 219860 412752
rect 219808 412709 219817 412743
rect 219817 412709 219851 412743
rect 219851 412709 219860 412743
rect 219808 412700 219860 412709
rect 219624 412632 219676 412684
rect 219808 412594 219860 412646
rect 219624 412496 219676 412548
rect 3148 409844 3200 409896
rect 50344 409844 50396 409896
rect 210424 407872 210476 407924
rect 213184 407872 213236 407924
rect 216680 407872 216732 407924
rect 210700 407124 210752 407176
rect 216772 407124 216824 407176
rect 219624 405832 219676 405884
rect 219716 405628 219768 405680
rect 425704 404336 425756 404388
rect 580172 404336 580224 404388
rect 219440 403087 219492 403096
rect 219440 403053 219449 403087
rect 219449 403053 219483 403087
rect 219483 403053 219492 403087
rect 219440 403044 219492 403053
rect 219532 402908 219584 402960
rect 219440 402883 219492 402892
rect 219440 402849 219449 402883
rect 219449 402849 219483 402883
rect 219483 402849 219492 402883
rect 219440 402840 219492 402849
rect 219532 402815 219584 402824
rect 219532 402781 219541 402815
rect 219541 402781 219575 402815
rect 219575 402781 219584 402815
rect 219532 402772 219584 402781
rect 197544 400052 197596 400104
rect 176568 399984 176620 400036
rect 187608 399984 187660 400036
rect 198832 399984 198884 400036
rect 184204 399916 184256 399968
rect 217416 399916 217468 399968
rect 115756 399848 115808 399900
rect 206376 399848 206428 399900
rect 217600 399848 217652 399900
rect 226340 399848 226392 399900
rect 119988 399780 120040 399832
rect 214656 399780 214708 399832
rect 217692 399780 217744 399832
rect 230480 399780 230532 399832
rect 113088 399712 113140 399764
rect 215944 399712 215996 399764
rect 217876 399712 217928 399764
rect 233240 399712 233292 399764
rect 52092 399644 52144 399696
rect 198924 399644 198976 399696
rect 199476 399644 199528 399696
rect 232044 399644 232096 399696
rect 56968 399576 57020 399628
rect 231952 399576 232004 399628
rect 59268 399508 59320 399560
rect 122932 399508 122984 399560
rect 180708 399508 180760 399560
rect 357624 399508 357676 399560
rect 52000 399440 52052 399492
rect 359004 399440 359056 399492
rect 57888 398760 57940 398812
rect 210424 398760 210476 398812
rect 218520 398760 218572 398812
rect 219532 398760 219584 398812
rect 224500 398760 224552 398812
rect 218152 398692 218204 398744
rect 219164 398556 219216 398608
rect 227720 398692 227772 398744
rect 219808 398624 219860 398676
rect 229284 398624 229336 398676
rect 226616 398556 226668 398608
rect 219348 398488 219400 398540
rect 226708 398488 226760 398540
rect 219716 398420 219768 398472
rect 229192 398420 229244 398472
rect 219624 398352 219676 398404
rect 229100 398352 229152 398404
rect 185584 398284 185636 398336
rect 196808 398284 196860 398336
rect 218336 398284 218388 398336
rect 227812 398284 227864 398336
rect 177948 398216 178000 398268
rect 210608 398216 210660 398268
rect 218244 398216 218296 398268
rect 228364 398216 228416 398268
rect 169668 398148 169720 398200
rect 210700 398148 210752 398200
rect 218060 398148 218112 398200
rect 228272 398148 228324 398200
rect 122748 398080 122800 398132
rect 196624 398080 196676 398132
rect 217784 398080 217836 398132
rect 228640 398080 228692 398132
rect 219440 398012 219492 398064
rect 226432 398012 226484 398064
rect 218428 397944 218480 397996
rect 226524 397944 226576 397996
rect 228088 397876 228140 397928
rect 218612 397808 218664 397860
rect 225420 397808 225472 397860
rect 228456 397740 228508 397792
rect 3424 397468 3476 397520
rect 143540 397468 143592 397520
rect 81992 397400 82044 397452
rect 224960 397400 225012 397452
rect 85488 397332 85540 397384
rect 229376 397332 229428 397384
rect 61476 397264 61528 397316
rect 278044 397264 278096 397316
rect 58808 397196 58860 397248
rect 109500 397196 109552 397248
rect 111248 397196 111300 397248
rect 137284 397196 137336 397248
rect 238024 397196 238076 397248
rect 239220 397196 239272 397248
rect 291844 397196 291896 397248
rect 298468 397196 298520 397248
rect 88800 397128 88852 397180
rect 94504 397128 94556 397180
rect 106464 397128 106516 397180
rect 134524 397128 134576 397180
rect 177304 397128 177356 397180
rect 237012 397128 237064 397180
rect 58992 397060 59044 397112
rect 99380 397060 99432 397112
rect 104072 397060 104124 397112
rect 113640 397060 113692 397112
rect 170404 397060 170456 397112
rect 184296 397060 184348 397112
rect 247684 397060 247736 397112
rect 80980 396992 81032 397044
rect 142804 396992 142856 397044
rect 173808 396992 173860 397044
rect 238116 396992 238168 397044
rect 90732 396924 90784 396976
rect 187792 396924 187844 396976
rect 196624 396924 196676 396976
rect 251272 396924 251324 396976
rect 58716 396856 58768 396908
rect 112076 396856 112128 396908
rect 115848 396856 115900 396908
rect 224776 396856 224828 396908
rect 58532 396788 58584 396840
rect 113180 396788 113232 396840
rect 118332 396788 118384 396840
rect 233424 396788 233476 396840
rect 58440 396720 58492 396772
rect 113732 396720 113784 396772
rect 117136 396720 117188 396772
rect 233332 396720 233384 396772
rect 240784 396720 240836 396772
rect 242900 396720 242952 396772
rect 249064 396720 249116 396772
rect 256884 396720 256936 396772
rect 268384 396720 268436 396772
rect 273260 396720 273312 396772
rect 287704 396720 287756 396772
rect 295892 396720 295944 396772
rect 307024 396720 307076 396772
rect 307852 396720 307904 396772
rect 96344 396652 96396 396704
rect 97264 396652 97316 396704
rect 105728 396652 105780 396704
rect 108304 396652 108356 396704
rect 231860 396652 231912 396704
rect 253204 396652 253256 396704
rect 254492 396652 254544 396704
rect 260104 396652 260156 396704
rect 260932 396652 260984 396704
rect 291936 396652 291988 396704
rect 292948 396652 293000 396704
rect 304264 396652 304316 396704
rect 305276 396652 305328 396704
rect 309784 396652 309836 396704
rect 315764 396652 315816 396704
rect 322204 396652 322256 396704
rect 323124 396652 323176 396704
rect 58900 396584 58952 396636
rect 95976 396584 96028 396636
rect 97356 396584 97408 396636
rect 102048 396584 102100 396636
rect 229468 396584 229520 396636
rect 92388 396516 92440 396568
rect 227904 396516 227956 396568
rect 246304 396516 246356 396568
rect 262036 396516 262088 396568
rect 59268 396448 59320 396500
rect 87604 396448 87656 396500
rect 100760 396448 100812 396500
rect 222108 396448 222160 396500
rect 276388 396448 276440 396500
rect 59084 396380 59136 396432
rect 94228 396380 94280 396432
rect 97632 396380 97684 396432
rect 106924 396380 106976 396432
rect 220084 396380 220136 396432
rect 273444 396380 273496 396432
rect 78312 396312 78364 396364
rect 222844 396312 222896 396364
rect 224868 396312 224920 396364
rect 278964 396312 279016 396364
rect 59728 396244 59780 396296
rect 236000 396244 236052 396296
rect 238208 396244 238260 396296
rect 272248 396244 272300 396296
rect 282184 396244 282236 396296
rect 325884 396244 325936 396296
rect 59452 396176 59504 396228
rect 240508 396176 240560 396228
rect 242256 396176 242308 396228
rect 259828 396176 259880 396228
rect 284944 396176 284996 396228
rect 289820 396176 289872 396228
rect 59544 396108 59596 396160
rect 252744 396108 252796 396160
rect 316684 396108 316736 396160
rect 343364 396108 343416 396160
rect 83372 396040 83424 396092
rect 87604 396040 87656 396092
rect 242164 395972 242216 396024
rect 247592 395972 247644 396024
rect 163872 395904 163924 395956
rect 222200 395904 222252 395956
rect 156420 395836 156472 395888
rect 215392 395836 215444 395888
rect 179328 395768 179380 395820
rect 241612 395768 241664 395820
rect 146024 395700 146076 395752
rect 209780 395700 209832 395752
rect 235264 395700 235316 395752
rect 249984 395700 250036 395752
rect 191748 395632 191800 395684
rect 268292 395632 268344 395684
rect 118608 395564 118660 395616
rect 197544 395564 197596 395616
rect 231124 395564 231176 395616
rect 265900 395564 265952 395616
rect 54852 395496 54904 395548
rect 138388 395496 138440 395548
rect 183284 395496 183336 395548
rect 185584 395496 185636 395548
rect 195888 395496 195940 395548
rect 276204 395496 276256 395548
rect 51908 395428 51960 395480
rect 91284 395428 91336 395480
rect 136272 395428 136324 395480
rect 227996 395428 228048 395480
rect 238116 395428 238168 395480
rect 273352 395428 273404 395480
rect 54944 395360 54996 395412
rect 123484 395360 123536 395412
rect 125968 395360 126020 395412
rect 228180 395360 228232 395412
rect 232504 395360 232556 395412
rect 270868 395360 270920 395412
rect 85028 395292 85080 395344
rect 233516 395292 233568 395344
rect 240876 395292 240928 395344
rect 283196 395292 283248 395344
rect 180524 393320 180576 393372
rect 183284 393320 183336 393372
rect 177396 388492 177448 388544
rect 180524 388492 180576 388544
rect 85488 378156 85540 378208
rect 580172 378156 580224 378208
rect 175280 377000 175332 377052
rect 177396 377000 177448 377052
rect 171140 375096 171192 375148
rect 175280 375096 175332 375148
rect 171140 372580 171192 372632
rect 164884 372512 164936 372564
rect 3424 371220 3476 371272
rect 144920 371220 144972 371272
rect 154488 367752 154540 367804
rect 228916 367752 228968 367804
rect 85396 364352 85448 364404
rect 579620 364352 579672 364404
rect 160100 359456 160152 359508
rect 164884 359456 164936 359508
rect 54760 358028 54812 358080
rect 147680 358028 147732 358080
rect 3148 357416 3200 357468
rect 147680 357416 147732 357468
rect 159364 357416 159416 357468
rect 160100 357416 160152 357468
rect 84108 351908 84160 351960
rect 580172 351908 580224 351960
rect 156604 346332 156656 346384
rect 159364 346332 159416 346384
rect 3332 345040 3384 345092
rect 146300 345040 146352 345092
rect 81348 324300 81400 324352
rect 580172 324300 580224 324352
rect 3424 318792 3476 318844
rect 147772 318792 147824 318844
rect 154580 311924 154632 311976
rect 156604 311924 156656 311976
rect 82728 311856 82780 311908
rect 579988 311856 580040 311908
rect 151084 306348 151136 306400
rect 154488 306348 154540 306400
rect 3240 304988 3292 305040
rect 150440 304988 150492 305040
rect 149704 299412 149756 299464
rect 151084 299412 151136 299464
rect 81256 298120 81308 298172
rect 580172 298120 580224 298172
rect 3424 292544 3476 292596
rect 149060 292544 149112 292596
rect 148324 282888 148376 282940
rect 149704 282888 149756 282940
rect 78588 271872 78640 271924
rect 580172 271872 580224 271924
rect 146944 271192 146996 271244
rect 148324 271192 148376 271244
rect 151728 266976 151780 267028
rect 212540 266976 212592 267028
rect 3056 266364 3108 266416
rect 150532 266432 150584 266484
rect 145564 266364 145616 266416
rect 146944 266364 146996 266416
rect 144184 262896 144236 262948
rect 145564 262896 145616 262948
rect 104716 261468 104768 261520
rect 229652 261468 229704 261520
rect 112996 258748 113048 258800
rect 360844 258748 360896 258800
rect 107476 258680 107528 258732
rect 376024 258680 376076 258732
rect 79968 258068 80020 258120
rect 580172 258068 580224 258120
rect 142804 256708 142856 256760
rect 144184 256708 144236 256760
rect 3424 253920 3476 253972
rect 153200 253920 153252 253972
rect 141424 251744 141476 251796
rect 142804 251744 142856 251796
rect 232688 250452 232740 250504
rect 317420 250452 317472 250504
rect 142896 249568 142948 249620
rect 226892 249568 226944 249620
rect 94504 249500 94556 249552
rect 180892 249500 180944 249552
rect 97356 249432 97408 249484
rect 195980 249432 196032 249484
rect 108304 249364 108356 249416
rect 207020 249364 207072 249416
rect 119896 249296 119948 249348
rect 223672 249296 223724 249348
rect 99196 249228 99248 249280
rect 225052 249228 225104 249280
rect 99288 249160 99340 249212
rect 230664 249160 230716 249212
rect 77116 249092 77168 249144
rect 233700 249092 233752 249144
rect 51816 249024 51868 249076
rect 259552 249024 259604 249076
rect 54208 248344 54260 248396
rect 129740 248344 129792 248396
rect 97264 248276 97316 248328
rect 176016 248276 176068 248328
rect 111708 248208 111760 248260
rect 193220 248208 193272 248260
rect 106924 248140 106976 248192
rect 198832 248140 198884 248192
rect 87604 248072 87656 248124
rect 171232 248072 171284 248124
rect 193128 248072 193180 248124
rect 316684 248072 316736 248124
rect 101956 248004 102008 248056
rect 229744 248004 229796 248056
rect 47584 247936 47636 247988
rect 142160 247936 142212 247988
rect 188988 247936 189040 247988
rect 342352 247936 342404 247988
rect 51724 247868 51776 247920
rect 265072 247868 265124 247920
rect 54576 247800 54628 247852
rect 277492 247800 277544 247852
rect 55864 247732 55916 247784
rect 310520 247732 310572 247784
rect 88248 247664 88300 247716
rect 580264 247664 580316 247716
rect 120724 247596 120776 247648
rect 196532 247596 196584 247648
rect 32404 246984 32456 247036
rect 140872 246984 140924 247036
rect 161388 246984 161440 247036
rect 233608 246984 233660 247036
rect 108856 246916 108908 246968
rect 229836 246916 229888 246968
rect 91008 246848 91060 246900
rect 228824 246848 228876 246900
rect 54484 246780 54536 246832
rect 280160 246780 280212 246832
rect 54300 246712 54352 246764
rect 287060 246712 287112 246764
rect 108856 246644 108908 246696
rect 388444 246644 388496 246696
rect 100668 246576 100720 246628
rect 382924 246576 382976 246628
rect 103336 246508 103388 246560
rect 385684 246508 385736 246560
rect 88156 246440 88208 246492
rect 378784 246440 378836 246492
rect 111708 246372 111760 246424
rect 412640 246372 412692 246424
rect 106188 246304 106240 246356
rect 542360 246304 542412 246356
rect 35164 246236 35216 246288
rect 132500 246236 132552 246288
rect 133788 246236 133840 246288
rect 228548 246236 228600 246288
rect 33784 246168 33836 246220
rect 126980 246168 127032 246220
rect 137284 246168 137336 246220
rect 212632 246168 212684 246220
rect 36544 246100 36596 246152
rect 129740 246100 129792 246152
rect 55956 246032 56008 246084
rect 140780 246032 140832 246084
rect 56048 245964 56100 246016
rect 120080 245964 120132 246016
rect 22744 245556 22796 245608
rect 129832 245556 129884 245608
rect 138572 245556 138624 245608
rect 141424 245624 141476 245676
rect 183468 245556 183520 245608
rect 232320 245556 232372 245608
rect 8208 245488 8260 245540
rect 127072 245488 127124 245540
rect 134524 245488 134576 245540
rect 208492 245488 208544 245540
rect 106096 245420 106148 245472
rect 228732 245420 228784 245472
rect 18604 245352 18656 245404
rect 142712 245352 142764 245404
rect 206928 245352 206980 245404
rect 287704 245352 287756 245404
rect 4804 245284 4856 245336
rect 138112 245284 138164 245336
rect 186228 245284 186280 245336
rect 357532 245284 357584 245336
rect 51632 245216 51684 245268
rect 266452 245216 266504 245268
rect 110328 245148 110380 245200
rect 377404 245148 377456 245200
rect 104808 245080 104860 245132
rect 374644 245080 374696 245132
rect 99288 245012 99340 245064
rect 370504 245012 370556 245064
rect 93584 244944 93636 244996
rect 381544 244944 381596 244996
rect 91008 244876 91060 244928
rect 443644 244876 443696 244928
rect 25504 244808 25556 244860
rect 132592 244808 132644 244860
rect 199384 244808 199436 244860
rect 232228 244808 232280 244860
rect 29644 244740 29696 244792
rect 135260 244740 135312 244792
rect 117136 244672 117188 244724
rect 213276 244672 213328 244724
rect 50344 244604 50396 244656
rect 145012 244604 145064 244656
rect 43444 244536 43496 244588
rect 138020 244536 138072 244588
rect 173716 244332 173768 244384
rect 177304 244332 177356 244384
rect 78496 244264 78548 244316
rect 579804 244264 579856 244316
rect 11704 244196 11756 244248
rect 128544 244196 128596 244248
rect 158628 244196 158680 244248
rect 218152 244196 218204 244248
rect 15844 244128 15896 244180
rect 137008 244128 137060 244180
rect 205548 244128 205600 244180
rect 291936 244128 291988 244180
rect 17224 244060 17276 244112
rect 139952 244060 140004 244112
rect 209688 244060 209740 244112
rect 302240 244060 302292 244112
rect 54392 243992 54444 244044
rect 285680 243992 285732 244044
rect 102048 243924 102100 243976
rect 371884 243924 371936 243976
rect 96528 243856 96580 243908
rect 367744 243856 367796 243908
rect 90916 243788 90968 243840
rect 363604 243788 363656 243840
rect 108764 243720 108816 243772
rect 429200 243720 429252 243772
rect 93492 243652 93544 243704
rect 431224 243652 431276 243704
rect 86776 243584 86828 243636
rect 425704 243584 425756 243636
rect 96436 243516 96488 243568
rect 449164 243516 449216 243568
rect 21364 243448 21416 243500
rect 134248 243448 134300 243500
rect 135904 243448 135956 243500
rect 138572 243448 138624 243500
rect 204168 243448 204220 243500
rect 242256 243448 242308 243500
rect 97908 243380 97960 243432
rect 209136 243380 209188 243432
rect 95148 243312 95200 243364
rect 206284 243312 206336 243364
rect 56324 243244 56376 243296
rect 165620 243244 165672 243296
rect 39304 243176 39356 243228
rect 135352 243176 135404 243228
rect 41328 243108 41380 243160
rect 125600 243108 125652 243160
rect 118608 243040 118660 243092
rect 201500 243040 201552 243092
rect 115756 242972 115808 243024
rect 198004 242972 198056 243024
rect 117044 242836 117096 242888
rect 226064 242836 226116 242888
rect 103244 242768 103296 242820
rect 214564 242768 214616 242820
rect 92388 242700 92440 242752
rect 204996 242700 205048 242752
rect 57060 242632 57112 242684
rect 169760 242632 169812 242684
rect 206836 242632 206888 242684
rect 263692 242632 263744 242684
rect 100576 242564 100628 242616
rect 213368 242564 213420 242616
rect 14464 242496 14516 242548
rect 131304 242496 131356 242548
rect 170404 242496 170456 242548
rect 194048 242496 194100 242548
rect 204076 242496 204128 242548
rect 284944 242496 284996 242548
rect 57152 242428 57204 242480
rect 183560 242428 183612 242480
rect 219348 242428 219400 242480
rect 320180 242428 320232 242480
rect 93676 242360 93728 242412
rect 230572 242360 230624 242412
rect 58164 242292 58216 242344
rect 266360 242292 266412 242344
rect 89628 242224 89680 242276
rect 358084 242224 358136 242276
rect 56232 242156 56284 242208
rect 88340 242156 88392 242208
rect 106096 242156 106148 242208
rect 446404 242156 446456 242208
rect 129648 242088 129700 242140
rect 225236 242088 225288 242140
rect 114468 242020 114520 242072
rect 209044 242020 209096 242072
rect 118516 241952 118568 242004
rect 204904 241952 204956 242004
rect 144828 241884 144880 241936
rect 225144 241884 225196 241936
rect 75828 241544 75880 241596
rect 242256 241544 242308 241596
rect 72332 241476 72384 241528
rect 240968 241476 241020 241528
rect 57888 241408 57940 241460
rect 58624 241408 58676 241460
rect 107568 241408 107620 241460
rect 230756 241408 230808 241460
rect 58256 241340 58308 241392
rect 181996 241340 182048 241392
rect 182088 241340 182140 241392
rect 184296 241340 184348 241392
rect 190368 241340 190420 241392
rect 196624 241340 196676 241392
rect 198648 241340 198700 241392
rect 249064 241340 249116 241392
rect 103428 241272 103480 241324
rect 229008 241272 229060 241324
rect 93768 241204 93820 241256
rect 225972 241204 226024 241256
rect 59176 241136 59228 241188
rect 198740 241136 198792 241188
rect 201408 241136 201460 241188
rect 258172 241136 258224 241188
rect 86868 241068 86920 241120
rect 232136 241068 232188 241120
rect 77208 241000 77260 241052
rect 226984 241000 227036 241052
rect 57152 240932 57204 240984
rect 210516 240932 210568 240984
rect 235356 240932 235408 240984
rect 270592 240932 270644 240984
rect 54668 240864 54720 240916
rect 244372 240864 244424 240916
rect 53104 240796 53156 240848
rect 249800 240796 249852 240848
rect 59636 240728 59688 240780
rect 274640 240728 274692 240780
rect 108948 240660 109000 240712
rect 226156 240660 226208 240712
rect 215208 240592 215260 240644
rect 238208 240592 238260 240644
rect 3424 240116 3476 240168
rect 106924 240116 106976 240168
rect 217232 240116 217284 240168
rect 226800 240116 226852 240168
rect 56140 227740 56192 227792
rect 59820 227740 59872 227792
rect 244924 225564 244976 225616
rect 255412 225564 255464 225616
rect 3516 215092 3568 215144
rect 7564 215092 7616 215144
rect 242256 206932 242308 206984
rect 580172 206932 580224 206984
rect 3056 202784 3108 202836
rect 29644 202784 29696 202836
rect 57336 201424 57388 201476
rect 58532 201424 58584 201476
rect 55036 198636 55088 198688
rect 57612 198636 57664 198688
rect 55128 195916 55180 195968
rect 57612 195916 57664 195968
rect 278044 193128 278096 193180
rect 580172 193128 580224 193180
rect 54760 190408 54812 190460
rect 57612 190408 57664 190460
rect 2780 188844 2832 188896
rect 4804 188844 4856 188896
rect 53196 184832 53248 184884
rect 57612 184832 57664 184884
rect 50620 183268 50672 183320
rect 57612 183268 57664 183320
rect 51632 180752 51684 180804
rect 56876 180752 56928 180804
rect 54852 172456 54904 172508
rect 57612 172456 57664 172508
rect 51724 169668 51776 169720
rect 57612 169668 57664 169720
rect 53288 166948 53340 167000
rect 57612 166948 57664 167000
rect 240968 166948 241020 167000
rect 580172 166948 580224 167000
rect 3240 164160 3292 164212
rect 11704 164160 11756 164212
rect 53380 163480 53432 163532
rect 57612 163480 57664 163532
rect 54208 161372 54260 161424
rect 57244 161372 57296 161424
rect 54300 158652 54352 158704
rect 57612 158652 57664 158704
rect 57428 155864 57480 155916
rect 58716 155864 58768 155916
rect 53472 153144 53524 153196
rect 57612 153144 57664 153196
rect 3516 150356 3568 150408
rect 18604 150356 18656 150408
rect 54392 150356 54444 150408
rect 57612 150356 57664 150408
rect 51816 144168 51868 144220
rect 57612 144168 57664 144220
rect 54944 142060 54996 142112
rect 57612 142060 57664 142112
rect 410524 139340 410576 139392
rect 580172 139340 580224 139392
rect 3516 137912 3568 137964
rect 15844 137912 15896 137964
rect 54484 136552 54536 136604
rect 57612 136552 57664 136604
rect 53564 133832 53616 133884
rect 57612 133832 57664 133884
rect 54576 132404 54628 132456
rect 57612 132404 57664 132456
rect 271144 126896 271196 126948
rect 580172 126896 580224 126948
rect 52184 118600 52236 118652
rect 57612 118600 57664 118652
rect 51908 115540 51960 115592
rect 57612 115540 57664 115592
rect 3148 111732 3200 111784
rect 14464 111732 14516 111784
rect 53656 110372 53708 110424
rect 57612 110372 57664 110424
rect 50804 107584 50856 107636
rect 57612 107584 57664 107636
rect 53104 104796 53156 104848
rect 57612 104796 57664 104848
rect 52000 102076 52052 102128
rect 57612 102076 57664 102128
rect 302884 100648 302936 100700
rect 580172 100648 580224 100700
rect 3516 97928 3568 97980
rect 25504 97928 25556 97980
rect 53748 90992 53800 91044
rect 57612 90992 57664 91044
rect 52092 88272 52144 88324
rect 57612 88272 57664 88324
rect 3516 85484 3568 85536
rect 17224 85484 17276 85536
rect 50896 85484 50948 85536
rect 57612 85484 57664 85536
rect 50988 79976 51040 80028
rect 57612 79976 57664 80028
rect 54668 78616 54720 78668
rect 57612 78616 57664 78668
rect 52276 75828 52328 75880
rect 57612 75828 57664 75880
rect 3516 71680 3568 71732
rect 21364 71680 21416 71732
rect 52368 70320 52420 70372
rect 57612 70320 57664 70372
rect 295984 60664 296036 60716
rect 580172 60664 580224 60716
rect 58624 60256 58676 60308
rect 59820 60256 59872 60308
rect 223672 59848 223724 59900
rect 224224 59848 224276 59900
rect 233240 59848 233292 59900
rect 233332 59848 233384 59900
rect 209688 59780 209740 59832
rect 252652 59780 252704 59832
rect 212632 59712 212684 59764
rect 258080 59712 258132 59764
rect 219164 59644 219216 59696
rect 291844 59644 291896 59696
rect 221004 59576 221056 59628
rect 304264 59576 304316 59628
rect 222476 59508 222528 59560
rect 309784 59508 309836 59560
rect 221832 59440 221884 59492
rect 313280 59440 313332 59492
rect 223948 59372 224000 59424
rect 322204 59372 322256 59424
rect 3056 59304 3108 59356
rect 36544 59304 36596 59356
rect 50712 59304 50764 59356
rect 211988 59304 212040 59356
rect 215944 59304 215996 59356
rect 227904 59304 227956 59356
rect 217140 59236 217192 59288
rect 227812 59236 227864 59288
rect 213184 59168 213236 59220
rect 221280 59168 221332 59220
rect 269120 59168 269172 59220
rect 218612 59100 218664 59152
rect 231860 59100 231912 59152
rect 222200 59032 222252 59084
rect 268384 59032 268436 59084
rect 219808 58964 219860 59016
rect 229100 58964 229152 59016
rect 214104 58896 214156 58948
rect 248420 58896 248472 58948
rect 211712 58828 211764 58880
rect 245660 58828 245712 58880
rect 207848 58760 207900 58812
rect 240784 58760 240836 58812
rect 217692 58692 217744 58744
rect 229468 58692 229520 58744
rect 211436 58624 211488 58676
rect 358912 58624 358964 58676
rect 209044 58556 209096 58608
rect 238024 58556 238076 58608
rect 208124 58488 208176 58540
rect 229284 58488 229336 58540
rect 210516 58420 210568 58472
rect 229376 58420 229428 58472
rect 260104 58352 260156 58404
rect 213552 58284 213604 58336
rect 229192 58284 229244 58336
rect 214380 58216 214432 58268
rect 263600 58216 263652 58268
rect 215576 58148 215628 58200
rect 251180 58148 251232 58200
rect 216772 58080 216824 58132
rect 227720 58080 227772 58132
rect 216220 58012 216272 58064
rect 224500 58012 224552 58064
rect 64512 57987 64564 57996
rect 64512 57953 64521 57987
rect 64521 57953 64555 57987
rect 64555 57953 64564 57987
rect 64512 57944 64564 57953
rect 28908 57808 28960 57860
rect 66904 57876 66956 57928
rect 68284 57876 68336 57928
rect 74080 57876 74132 57928
rect 58348 57808 58400 57860
rect 209320 57876 209372 57928
rect 220084 57876 220136 57928
rect 224684 57876 224736 57928
rect 87144 57808 87196 57860
rect 105452 57808 105504 57860
rect 106280 57808 106332 57860
rect 107568 57808 107620 57860
rect 109500 57808 109552 57860
rect 110328 57808 110380 57860
rect 133144 57808 133196 57860
rect 26148 57740 26200 57792
rect 66352 57740 66404 57792
rect 67088 57740 67140 57792
rect 70768 57740 70820 57792
rect 74356 57740 74408 57792
rect 101496 57740 101548 57792
rect 24768 57672 24820 57724
rect 65984 57672 66036 57724
rect 66076 57672 66128 57724
rect 66628 57672 66680 57724
rect 70308 57672 70360 57724
rect 77668 57672 77720 57724
rect 90548 57672 90600 57724
rect 91008 57672 91060 57724
rect 91652 57672 91704 57724
rect 19248 57604 19300 57656
rect 16488 57536 16540 57588
rect 63592 57536 63644 57588
rect 69572 57604 69624 57656
rect 70216 57604 70268 57656
rect 77300 57604 77352 57656
rect 78772 57604 78824 57656
rect 79508 57604 79560 57656
rect 92848 57604 92900 57656
rect 93584 57604 93636 57656
rect 94320 57672 94372 57724
rect 95148 57672 95200 57724
rect 95792 57672 95844 57724
rect 97540 57672 97592 57724
rect 99656 57672 99708 57724
rect 100576 57672 100628 57724
rect 101220 57672 101272 57724
rect 101864 57672 101916 57724
rect 124864 57740 124916 57792
rect 125600 57740 125652 57792
rect 126888 57740 126940 57792
rect 127440 57740 127492 57792
rect 128176 57740 128228 57792
rect 131580 57740 131632 57792
rect 136732 57808 136784 57860
rect 138112 57808 138164 57860
rect 135996 57740 136048 57792
rect 138756 57808 138808 57860
rect 149428 57808 149480 57860
rect 161572 57808 161624 57860
rect 161940 57808 161992 57860
rect 170312 57808 170364 57860
rect 170956 57808 171008 57860
rect 201868 57808 201920 57860
rect 202604 57808 202656 57860
rect 203708 57808 203760 57860
rect 204076 57808 204128 57860
rect 204536 57808 204588 57860
rect 205364 57808 205416 57860
rect 206100 57808 206152 57860
rect 206928 57808 206980 57860
rect 220360 57808 220412 57860
rect 225144 57808 225196 57860
rect 125876 57672 125928 57724
rect 126704 57672 126756 57724
rect 127716 57672 127768 57724
rect 128084 57672 128136 57724
rect 130108 57672 130160 57724
rect 130936 57672 130988 57724
rect 131304 57672 131356 57724
rect 132224 57672 132276 57724
rect 132500 57672 132552 57724
rect 123484 57604 123536 57656
rect 123944 57604 123996 57656
rect 126520 57604 126572 57656
rect 126796 57604 126848 57656
rect 127072 57604 127124 57656
rect 127900 57604 127952 57656
rect 128636 57604 128688 57656
rect 129556 57604 129608 57656
rect 130384 57604 130436 57656
rect 130844 57604 130896 57656
rect 131856 57604 131908 57656
rect 132408 57604 132460 57656
rect 132776 57604 132828 57656
rect 133696 57604 133748 57656
rect 65616 57536 65668 57588
rect 67548 57536 67600 57588
rect 13728 57468 13780 57520
rect 63316 57468 63368 57520
rect 64144 57468 64196 57520
rect 15108 57400 15160 57452
rect 63500 57400 63552 57452
rect 6828 57332 6880 57384
rect 61568 57332 61620 57384
rect 62764 57332 62816 57384
rect 66904 57468 66956 57520
rect 69020 57468 69072 57520
rect 72240 57468 72292 57520
rect 74724 57536 74776 57588
rect 75644 57536 75696 57588
rect 77208 57536 77260 57588
rect 79140 57536 79192 57588
rect 92572 57536 92624 57588
rect 93676 57536 93728 57588
rect 94044 57536 94096 57588
rect 94872 57536 94924 57588
rect 95240 57536 95292 57588
rect 96528 57536 96580 57588
rect 96712 57536 96764 57588
rect 97724 57536 97776 57588
rect 98184 57536 98236 57588
rect 99104 57536 99156 57588
rect 100024 57536 100076 57588
rect 100484 57536 100536 57588
rect 101772 57536 101824 57588
rect 102048 57536 102100 57588
rect 102692 57536 102744 57588
rect 103428 57536 103480 57588
rect 103888 57536 103940 57588
rect 104716 57536 104768 57588
rect 105360 57536 105412 57588
rect 106188 57536 106240 57588
rect 106556 57536 106608 57588
rect 107476 57536 107528 57588
rect 109776 57536 109828 57588
rect 110144 57536 110196 57588
rect 111892 57536 111944 57588
rect 112996 57536 113048 57588
rect 135260 57604 135312 57656
rect 134524 57536 134576 57588
rect 135168 57536 135220 57588
rect 135720 57536 135772 57588
rect 136456 57536 136508 57588
rect 136640 57672 136692 57724
rect 137836 57672 137888 57724
rect 140320 57740 140372 57792
rect 140504 57740 140556 57792
rect 145840 57672 145892 57724
rect 76748 57468 76800 57520
rect 90180 57468 90232 57520
rect 90916 57468 90968 57520
rect 64420 57400 64472 57452
rect 67824 57400 67876 57452
rect 71044 57400 71096 57452
rect 73068 57400 73120 57452
rect 65524 57332 65576 57384
rect 75000 57332 75052 57384
rect 75184 57400 75236 57452
rect 78496 57400 78548 57452
rect 88616 57400 88668 57452
rect 95516 57468 95568 57520
rect 96344 57468 96396 57520
rect 97264 57468 97316 57520
rect 100852 57400 100904 57452
rect 102048 57400 102100 57452
rect 102324 57468 102376 57520
rect 135444 57468 135496 57520
rect 136548 57468 136600 57520
rect 142804 57536 142856 57588
rect 147220 57604 147272 57656
rect 148600 57604 148652 57656
rect 162124 57672 162176 57724
rect 164608 57740 164660 57792
rect 170864 57740 170916 57792
rect 214564 57740 214616 57792
rect 220636 57740 220688 57792
rect 225696 57740 225748 57792
rect 166264 57672 166316 57724
rect 166448 57672 166500 57724
rect 213184 57672 213236 57724
rect 217416 57672 217468 57724
rect 225236 57672 225288 57724
rect 157524 57604 157576 57656
rect 167000 57604 167052 57656
rect 168196 57604 168248 57656
rect 213276 57604 213328 57656
rect 215300 57604 215352 57656
rect 147036 57468 147088 57520
rect 150348 57468 150400 57520
rect 103244 57400 103296 57452
rect 142620 57400 142672 57452
rect 143172 57400 143224 57452
rect 78220 57332 78272 57384
rect 10968 57264 11020 57316
rect 62396 57264 62448 57316
rect 63684 57264 63736 57316
rect 64604 57264 64656 57316
rect 73160 57264 73212 57316
rect 86868 57264 86920 57316
rect 101404 57332 101456 57384
rect 103520 57332 103572 57384
rect 104808 57332 104860 57384
rect 108580 57332 108632 57384
rect 108948 57332 109000 57384
rect 109224 57332 109276 57384
rect 110236 57332 110288 57384
rect 110696 57332 110748 57384
rect 111432 57332 111484 57384
rect 89812 57264 89864 57316
rect 90732 57264 90784 57316
rect 4068 57196 4120 57248
rect 60924 57196 60976 57248
rect 64236 57196 64288 57248
rect 33048 57128 33100 57180
rect 68100 57128 68152 57180
rect 70492 57196 70544 57248
rect 71688 57196 71740 57248
rect 77944 57196 77996 57248
rect 72608 57128 72660 57180
rect 75828 57128 75880 57180
rect 78864 57128 78916 57180
rect 85396 57128 85448 57180
rect 98644 57264 98696 57316
rect 100668 57264 100720 57316
rect 144184 57332 144236 57384
rect 145012 57332 145064 57384
rect 35808 57060 35860 57112
rect 68652 57060 68704 57112
rect 68928 57060 68980 57112
rect 77024 57060 77076 57112
rect 80244 57060 80296 57112
rect 80428 57060 80480 57112
rect 83556 57060 83608 57112
rect 94228 57196 94280 57248
rect 96620 57196 96672 57248
rect 144092 57264 144144 57316
rect 155500 57332 155552 57384
rect 156052 57468 156104 57520
rect 157156 57468 157208 57520
rect 167368 57536 167420 57588
rect 156880 57400 156932 57452
rect 157248 57400 157300 57452
rect 201040 57468 201092 57520
rect 201316 57468 201368 57520
rect 202512 57468 202564 57520
rect 202788 57468 202840 57520
rect 203064 57468 203116 57520
rect 203892 57468 203944 57520
rect 205180 57468 205232 57520
rect 205456 57468 205508 57520
rect 205732 57468 205784 57520
rect 206744 57468 206796 57520
rect 215944 57468 215996 57520
rect 218888 57536 218940 57588
rect 227996 57536 228048 57588
rect 217968 57468 218020 57520
rect 228548 57468 228600 57520
rect 220084 57400 220136 57452
rect 182548 57332 182600 57384
rect 183284 57332 183336 57384
rect 184020 57332 184072 57384
rect 184664 57332 184716 57384
rect 184940 57332 184992 57384
rect 185860 57332 185912 57384
rect 186504 57332 186556 57384
rect 187608 57332 187660 57384
rect 187792 57332 187844 57384
rect 188528 57332 188580 57384
rect 189080 57332 189132 57384
rect 190092 57332 190144 57384
rect 190552 57332 190604 57384
rect 191564 57332 191616 57384
rect 192392 57332 192444 57384
rect 193036 57332 193088 57384
rect 193220 57332 193272 57384
rect 193680 57332 193732 57384
rect 195336 57332 195388 57384
rect 195888 57332 195940 57384
rect 196532 57332 196584 57384
rect 197084 57332 197136 57384
rect 197452 57332 197504 57384
rect 198464 57332 198516 57384
rect 199200 57332 199252 57384
rect 199844 57332 199896 57384
rect 200120 57332 200172 57384
rect 201224 57332 201276 57384
rect 201592 57332 201644 57384
rect 202788 57332 202840 57384
rect 203432 57332 203484 57384
rect 204168 57332 204220 57384
rect 204260 57332 204312 57384
rect 205548 57332 205600 57384
rect 206376 57332 206428 57384
rect 391204 57332 391256 57384
rect 171232 57264 171284 57316
rect 172244 57264 172296 57316
rect 173992 57264 174044 57316
rect 174912 57264 174964 57316
rect 175372 57264 175424 57316
rect 176568 57264 176620 57316
rect 176844 57264 176896 57316
rect 177672 57264 177724 57316
rect 178960 57264 179012 57316
rect 179328 57264 179380 57316
rect 142252 57196 142304 57248
rect 142344 57196 142396 57248
rect 92204 57128 92256 57180
rect 105544 57128 105596 57180
rect 107752 57128 107804 57180
rect 108948 57128 109000 57180
rect 111340 57128 111392 57180
rect 111708 57128 111760 57180
rect 113364 57128 113416 57180
rect 114468 57128 114520 57180
rect 115480 57128 115532 57180
rect 115756 57128 115808 57180
rect 116032 57128 116084 57180
rect 116860 57128 116912 57180
rect 119252 57128 119304 57180
rect 119620 57128 119672 57180
rect 121736 57128 121788 57180
rect 122564 57128 122616 57180
rect 134064 57128 134116 57180
rect 136916 57128 136968 57180
rect 163780 57196 163832 57248
rect 171324 57196 171376 57248
rect 172428 57196 172480 57248
rect 173900 57196 173952 57248
rect 175096 57196 175148 57248
rect 177488 57196 177540 57248
rect 177856 57196 177908 57248
rect 178316 57196 178368 57248
rect 179236 57196 179288 57248
rect 179880 57196 179932 57248
rect 382924 57264 382976 57316
rect 180708 57196 180760 57248
rect 387064 57196 387116 57248
rect 91376 57060 91428 57112
rect 92388 57060 92440 57112
rect 98828 57060 98880 57112
rect 99288 57060 99340 57112
rect 108028 57060 108080 57112
rect 108672 57060 108724 57112
rect 39948 56992 40000 57044
rect 43444 56924 43496 56976
rect 66996 56992 67048 57044
rect 76104 56992 76156 57044
rect 94596 56992 94648 57044
rect 95056 56992 95108 57044
rect 102876 56992 102928 57044
rect 105084 56992 105136 57044
rect 53748 56856 53800 56908
rect 69848 56924 69900 56976
rect 50344 56788 50396 56840
rect 62948 56720 63000 56772
rect 64788 56720 64840 56772
rect 57244 56652 57296 56704
rect 64328 56652 64380 56704
rect 73436 56924 73488 56976
rect 82728 56924 82780 56976
rect 87696 56924 87748 56976
rect 87788 56924 87840 56976
rect 102784 56924 102836 56976
rect 105636 56924 105688 56976
rect 106096 56924 106148 56976
rect 106832 56992 106884 57044
rect 114560 57060 114612 57112
rect 115664 57060 115716 57112
rect 119068 57060 119120 57112
rect 119896 57060 119948 57112
rect 120540 57060 120592 57112
rect 137284 57060 137336 57112
rect 141332 57060 141384 57112
rect 143080 57060 143132 57112
rect 144368 57060 144420 57112
rect 146760 57060 146812 57112
rect 110420 56992 110472 57044
rect 111708 56992 111760 57044
rect 116952 56992 117004 57044
rect 117136 56992 117188 57044
rect 120264 56992 120316 57044
rect 121276 56992 121328 57044
rect 121460 56992 121512 57044
rect 142712 56992 142764 57044
rect 152096 56992 152148 57044
rect 117596 56924 117648 56976
rect 133512 56924 133564 56976
rect 84476 56856 84528 56908
rect 88892 56856 88944 56908
rect 96988 56856 97040 56908
rect 97908 56856 97960 56908
rect 104164 56856 104216 56908
rect 116400 56856 116452 56908
rect 116952 56856 117004 56908
rect 118424 56856 118476 56908
rect 129004 56856 129056 56908
rect 130016 56856 130068 56908
rect 141424 56924 141476 56976
rect 150900 56924 150952 56976
rect 151268 56924 151320 56976
rect 137928 56856 137980 56908
rect 70400 56788 70452 56840
rect 74540 56788 74592 56840
rect 80888 56788 80940 56840
rect 83188 56788 83240 56840
rect 84752 56788 84804 56840
rect 87604 56788 87656 56840
rect 122012 56788 122064 56840
rect 122748 56788 122800 56840
rect 129740 56788 129792 56840
rect 68376 56720 68428 56772
rect 74908 56720 74960 56772
rect 82084 56720 82136 56772
rect 83464 56720 83516 56772
rect 84200 56720 84252 56772
rect 86224 56720 86276 56772
rect 114008 56720 114060 56772
rect 122932 56720 122984 56772
rect 124036 56720 124088 56772
rect 124404 56720 124456 56772
rect 125324 56720 125376 56772
rect 129188 56720 129240 56772
rect 129648 56720 129700 56772
rect 62856 56584 62908 56636
rect 29644 56516 29696 56568
rect 63040 56516 63092 56568
rect 64604 56516 64656 56568
rect 65708 56584 65760 56636
rect 65984 56584 66036 56636
rect 67456 56584 67508 56636
rect 71504 56652 71556 56704
rect 81808 56652 81860 56704
rect 82728 56652 82780 56704
rect 83004 56652 83056 56704
rect 84016 56652 84068 56704
rect 85948 56652 86000 56704
rect 86868 56652 86920 56704
rect 88340 56652 88392 56704
rect 89444 56652 89496 56704
rect 123024 56652 123076 56704
rect 124128 56652 124180 56704
rect 124220 56652 124272 56704
rect 125048 56652 125100 56704
rect 70952 56584 71004 56636
rect 71044 56584 71096 56636
rect 75552 56584 75604 56636
rect 80612 56584 80664 56636
rect 81256 56584 81308 56636
rect 81532 56584 81584 56636
rect 82544 56584 82596 56636
rect 83280 56584 83332 56636
rect 83924 56584 83976 56636
rect 85672 56584 85724 56636
rect 86776 56584 86828 56636
rect 87512 56584 87564 56636
rect 88248 56584 88300 56636
rect 88984 56584 89036 56636
rect 89536 56584 89588 56636
rect 133972 56788 134024 56840
rect 135076 56788 135128 56840
rect 140044 56788 140096 56840
rect 151912 56856 151964 56908
rect 153936 56856 153988 56908
rect 146944 56788 146996 56840
rect 139676 56720 139728 56772
rect 147680 56720 147732 56772
rect 134248 56652 134300 56704
rect 134432 56652 134484 56704
rect 150532 56788 150584 56840
rect 153016 56788 153068 56840
rect 155224 56788 155276 56840
rect 147864 56720 147916 56772
rect 133328 56584 133380 56636
rect 136732 56584 136784 56636
rect 137928 56584 137980 56636
rect 138388 56584 138440 56636
rect 139124 56584 139176 56636
rect 139584 56584 139636 56636
rect 140872 56584 140924 56636
rect 141148 56584 141200 56636
rect 141976 56584 142028 56636
rect 143816 56584 143868 56636
rect 144460 56584 144512 56636
rect 145288 56584 145340 56636
rect 146208 56584 146260 56636
rect 148324 56652 148376 56704
rect 151820 56652 151872 56704
rect 153016 56652 153068 56704
rect 147956 56584 148008 56636
rect 148968 56584 149020 56636
rect 150624 56584 150676 56636
rect 151728 56584 151780 56636
rect 152464 56584 152516 56636
rect 153108 56584 153160 56636
rect 153292 56720 153344 56772
rect 156604 56856 156656 56908
rect 157708 56856 157760 56908
rect 173164 57128 173216 57180
rect 173624 57128 173676 57180
rect 175924 57128 175976 57180
rect 176292 57128 176344 57180
rect 169116 57060 169168 57112
rect 177120 57128 177172 57180
rect 177948 57128 178000 57180
rect 216036 57128 216088 57180
rect 223396 57128 223448 57180
rect 233608 57128 233660 57180
rect 172520 56992 172572 57044
rect 172704 56992 172756 57044
rect 178040 56992 178092 57044
rect 170036 56924 170088 56976
rect 174544 56924 174596 56976
rect 174636 56924 174688 56976
rect 217324 57060 217376 57112
rect 230480 57060 230532 57112
rect 220176 56992 220228 57044
rect 185768 56924 185820 56976
rect 186136 56924 186188 56976
rect 186320 56924 186372 56976
rect 186688 56924 186740 56976
rect 187884 56924 187936 56976
rect 188896 56924 188948 56976
rect 154212 56652 154264 56704
rect 154488 56652 154540 56704
rect 158996 56720 159048 56772
rect 159824 56720 159876 56772
rect 169024 56788 169076 56840
rect 173256 56788 173308 56840
rect 174820 56788 174872 56840
rect 175188 56788 175240 56840
rect 180156 56788 180208 56840
rect 180708 56788 180760 56840
rect 182272 56856 182324 56908
rect 183376 56856 183428 56908
rect 210424 56924 210476 56976
rect 215024 56924 215076 56976
rect 228732 56924 228784 56976
rect 192116 56856 192168 56908
rect 192944 56856 192996 56908
rect 193496 56856 193548 56908
rect 194140 56856 194192 56908
rect 194784 56856 194836 56908
rect 195704 56856 195756 56908
rect 196256 56856 196308 56908
rect 196900 56856 196952 56908
rect 197636 56856 197688 56908
rect 198648 56856 198700 56908
rect 198924 56856 198976 56908
rect 199936 56856 199988 56908
rect 207020 56856 207072 56908
rect 242164 56856 242216 56908
rect 184204 56788 184256 56840
rect 189540 56788 189592 56840
rect 190368 56788 190420 56840
rect 190828 56788 190880 56840
rect 191380 56788 191432 56840
rect 193312 56788 193364 56840
rect 194416 56788 194468 56840
rect 209136 56788 209188 56840
rect 210884 56788 210936 56840
rect 233240 56788 233292 56840
rect 170496 56720 170548 56772
rect 175648 56720 175700 56772
rect 176476 56720 176528 56772
rect 188344 56720 188396 56772
rect 207572 56720 207624 56772
rect 229560 56720 229612 56772
rect 157800 56652 157852 56704
rect 158628 56652 158680 56704
rect 158904 56652 158956 56704
rect 159640 56652 159692 56704
rect 160468 56652 160520 56704
rect 161388 56652 161440 56704
rect 34428 56448 34480 56500
rect 68192 56448 68244 56500
rect 156328 56584 156380 56636
rect 156972 56584 157024 56636
rect 158076 56584 158128 56636
rect 158536 56584 158588 56636
rect 159548 56584 159600 56636
rect 159916 56584 159968 56636
rect 160744 56584 160796 56636
rect 161296 56584 161348 56636
rect 161664 56584 161716 56636
rect 162584 56584 162636 56636
rect 162860 56584 162912 56636
rect 164056 56584 164108 56636
rect 154488 56516 154540 56568
rect 166356 56652 166408 56704
rect 164332 56584 164384 56636
rect 165160 56584 165212 56636
rect 165252 56584 165304 56636
rect 165436 56584 165488 56636
rect 166172 56584 166224 56636
rect 166908 56584 166960 56636
rect 170404 56652 170456 56704
rect 169116 56584 169168 56636
rect 172980 56652 173032 56704
rect 173808 56652 173860 56704
rect 179788 56652 179840 56704
rect 180616 56652 180668 56704
rect 186964 56652 187016 56704
rect 209044 56652 209096 56704
rect 209964 56652 210016 56704
rect 230572 56652 230624 56704
rect 179512 56584 179564 56636
rect 185216 56584 185268 56636
rect 185952 56584 186004 56636
rect 212908 56584 212960 56636
rect 225052 56584 225104 56636
rect 171508 56516 171560 56568
rect 436744 56516 436796 56568
rect 181076 56448 181128 56500
rect 454684 56448 454736 56500
rect 30288 56380 30340 56432
rect 21364 56312 21416 56364
rect 60372 56312 60424 56364
rect 183744 56380 183796 56432
rect 468484 56380 468536 56432
rect 65984 56312 66036 56364
rect 182824 56312 182876 56364
rect 461584 56312 461636 56364
rect 27528 56244 27580 56296
rect 66076 56244 66128 56296
rect 184848 56244 184900 56296
rect 472624 56244 472676 56296
rect 22836 56176 22888 56228
rect 65432 56176 65484 56228
rect 185492 56176 185544 56228
rect 475384 56176 475436 56228
rect 17868 56108 17920 56160
rect 64052 56108 64104 56160
rect 187332 56108 187384 56160
rect 479524 56108 479576 56160
rect 8208 56040 8260 56092
rect 61844 56040 61896 56092
rect 182088 56040 182140 56092
rect 483020 56040 483072 56092
rect 4804 55972 4856 56024
rect 60648 55972 60700 56024
rect 93124 55972 93176 56024
rect 112444 55972 112496 56024
rect 186596 55972 186648 56024
rect 500960 55972 501012 56024
rect 56140 55904 56192 55956
rect 580264 55904 580316 55956
rect 11704 55836 11756 55888
rect 60096 55836 60148 55888
rect 99380 55836 99432 55888
rect 152464 55836 152516 55888
rect 189356 55836 189408 55888
rect 512644 55836 512696 55888
rect 41328 55768 41380 55820
rect 69940 55768 69992 55820
rect 167644 55768 167696 55820
rect 425704 55768 425756 55820
rect 48228 55700 48280 55752
rect 71964 55700 72016 55752
rect 163136 55700 163188 55752
rect 407764 55700 407816 55752
rect 52368 55632 52420 55684
rect 72884 55632 72936 55684
rect 116676 55632 116728 55684
rect 224960 55632 225012 55684
rect 55128 55564 55180 55616
rect 73804 55564 73856 55616
rect 114928 55564 114980 55616
rect 218060 55564 218112 55616
rect 59268 55496 59320 55548
rect 70400 55496 70452 55548
rect 113088 55496 113140 55548
rect 209780 55496 209832 55548
rect 133512 55428 133564 55480
rect 227720 55428 227772 55480
rect 112168 55360 112220 55412
rect 207020 55360 207072 55412
rect 129740 55292 129792 55344
rect 213920 55292 213972 55344
rect 139952 55156 140004 55208
rect 316040 55156 316092 55208
rect 140780 55088 140832 55140
rect 320180 55088 320232 55140
rect 141700 55020 141752 55072
rect 324320 55020 324372 55072
rect 142528 54952 142580 55004
rect 327080 54952 327132 55004
rect 162308 54884 162360 54936
rect 405740 54884 405792 54936
rect 164148 54816 164200 54868
rect 412640 54816 412692 54868
rect 164976 54748 165028 54800
rect 414664 54748 414716 54800
rect 167736 54680 167788 54732
rect 427820 54680 427872 54732
rect 189540 54612 189592 54664
rect 485044 54612 485096 54664
rect 187976 54544 188028 54596
rect 507860 54544 507912 54596
rect 37188 54476 37240 54528
rect 69204 54476 69256 54528
rect 193404 54476 193456 54528
rect 530584 54476 530636 54528
rect 139032 54408 139084 54460
rect 313280 54408 313332 54460
rect 140320 54340 140372 54392
rect 309140 54340 309192 54392
rect 137192 54272 137244 54324
rect 306380 54272 306432 54324
rect 136640 54204 136692 54256
rect 302240 54204 302292 54256
rect 134064 54136 134116 54188
rect 231860 54136 231912 54188
rect 155868 54068 155920 54120
rect 222844 54068 222896 54120
rect 155500 53932 155552 53984
rect 155868 53932 155920 53984
rect 149152 53728 149204 53780
rect 353300 53728 353352 53780
rect 165804 53660 165856 53712
rect 418804 53660 418856 53712
rect 166724 53592 166776 53644
rect 421564 53592 421616 53644
rect 187792 53524 187844 53576
rect 447784 53524 447836 53576
rect 168380 53456 168432 53508
rect 430580 53456 430632 53508
rect 186504 53388 186556 53440
rect 450544 53388 450596 53440
rect 171324 53320 171376 53372
rect 445760 53320 445812 53372
rect 186320 53252 186372 53304
rect 502340 53252 502392 53304
rect 191932 53184 191984 53236
rect 519544 53184 519596 53236
rect 190920 53116 190972 53168
rect 520280 53116 520332 53168
rect 192116 53048 192168 53100
rect 526444 53048 526496 53100
rect 143448 52980 143500 53032
rect 331220 52980 331272 53032
rect 124220 52912 124272 52964
rect 258080 52912 258132 52964
rect 123208 52844 123260 52896
rect 251180 52844 251232 52896
rect 118884 52776 118936 52828
rect 233240 52776 233292 52828
rect 117688 52708 117740 52760
rect 229100 52708 229152 52760
rect 144644 52368 144696 52420
rect 335360 52368 335412 52420
rect 145564 52300 145616 52352
rect 339500 52300 339552 52352
rect 146484 52232 146536 52284
rect 342260 52232 342312 52284
rect 147404 52164 147456 52216
rect 346400 52164 346452 52216
rect 148232 52096 148284 52148
rect 349160 52096 349212 52148
rect 150072 52028 150124 52080
rect 357440 52028 357492 52080
rect 168748 51960 168800 52012
rect 431960 51960 432012 52012
rect 169944 51892 169996 51944
rect 434720 51892 434772 51944
rect 174084 51824 174136 51876
rect 452660 51824 452712 51876
rect 193680 51756 193732 51808
rect 528560 51756 528612 51808
rect 97540 51688 97592 51740
rect 142160 51688 142212 51740
rect 200396 51688 200448 51740
rect 544384 51688 544436 51740
rect 144368 51620 144420 51672
rect 328460 51620 328512 51672
rect 123024 51552 123076 51604
rect 253940 51552 253992 51604
rect 119252 51484 119304 51536
rect 236000 51484 236052 51536
rect 142252 51416 142304 51468
rect 240140 51416 240192 51468
rect 159088 51008 159140 51060
rect 393320 51008 393372 51060
rect 170312 50940 170364 50992
rect 438860 50940 438912 50992
rect 173072 50872 173124 50924
rect 443644 50872 443696 50924
rect 173992 50804 174044 50856
rect 456892 50804 456944 50856
rect 193496 50736 193548 50788
rect 489184 50736 489236 50788
rect 197636 50668 197688 50720
rect 533344 50668 533396 50720
rect 199292 50600 199344 50652
rect 537484 50600 537536 50652
rect 194876 50532 194928 50584
rect 535460 50532 535512 50584
rect 196164 50464 196216 50516
rect 539600 50464 539652 50516
rect 196624 50396 196676 50448
rect 542360 50396 542412 50448
rect 197728 50328 197780 50380
rect 546500 50328 546552 50380
rect 150900 50260 150952 50312
rect 322940 50260 322992 50312
rect 137928 50192 137980 50244
rect 284300 50192 284352 50244
rect 150624 49648 150676 49700
rect 291200 49648 291252 49700
rect 151820 49580 151872 49632
rect 298100 49580 298152 49632
rect 139676 49512 139728 49564
rect 293960 49512 294012 49564
rect 155868 49444 155920 49496
rect 311900 49444 311952 49496
rect 147956 49376 148008 49428
rect 305000 49376 305052 49428
rect 172520 49308 172572 49360
rect 340880 49308 340932 49360
rect 161572 49240 161624 49292
rect 329840 49240 329892 49292
rect 140872 49172 140924 49224
rect 316132 49172 316184 49224
rect 154856 49104 154908 49156
rect 375380 49104 375432 49156
rect 157800 49036 157852 49088
rect 382280 49036 382332 49088
rect 160376 48968 160428 49020
rect 396724 48968 396776 49020
rect 147404 48900 147456 48952
rect 276020 48900 276072 48952
rect 158444 47948 158496 48000
rect 388444 47948 388496 48000
rect 179512 47880 179564 47932
rect 411260 47880 411312 47932
rect 161112 47812 161164 47864
rect 400220 47812 400272 47864
rect 164056 47744 164108 47796
rect 407120 47744 407172 47796
rect 188344 47676 188396 47728
rect 432052 47676 432104 47728
rect 210424 47608 210476 47660
rect 460940 47608 460992 47660
rect 165344 47540 165396 47592
rect 418160 47540 418212 47592
rect 287704 46860 287756 46912
rect 580172 46860 580224 46912
rect 3516 45500 3568 45552
rect 40684 45500 40736 45552
rect 3516 33056 3568 33108
rect 22744 33056 22796 33108
rect 55772 33056 55824 33108
rect 580172 33056 580224 33108
rect 216036 24148 216088 24200
rect 447140 24148 447192 24200
rect 220176 24080 220228 24132
rect 467840 24080 467892 24132
rect 86592 22720 86644 22772
rect 103520 22720 103572 22772
rect 217324 22720 217376 22772
rect 454040 22720 454092 22772
rect 214564 21360 214616 21412
rect 440240 21360 440292 21412
rect 3516 20612 3568 20664
rect 33784 20612 33836 20664
rect 55680 20612 55732 20664
rect 580172 20612 580224 20664
rect 186964 20204 187016 20256
rect 357532 20204 357584 20256
rect 213276 20136 213328 20188
rect 404360 20136 404412 20188
rect 184204 20068 184256 20120
rect 386420 20068 386472 20120
rect 220084 20000 220136 20052
rect 425060 20000 425112 20052
rect 213184 19932 213236 19984
rect 422300 19932 422352 19984
rect 147036 19252 147088 19304
rect 287060 19252 287112 19304
rect 209136 19184 209188 19236
rect 365720 19184 365772 19236
rect 173256 19116 173308 19168
rect 336740 19116 336792 19168
rect 162124 19048 162176 19100
rect 332600 19048 332652 19100
rect 169116 18980 169168 19032
rect 343640 18980 343692 19032
rect 169024 18912 169076 18964
rect 347780 18912 347832 18964
rect 170496 18844 170548 18896
rect 350540 18844 350592 18896
rect 166356 18776 166408 18828
rect 354680 18776 354732 18828
rect 173164 18708 173216 18760
rect 361580 18708 361632 18760
rect 155224 18640 155276 18692
rect 368480 18640 368532 18692
rect 88984 18572 89036 18624
rect 96620 18572 96672 18624
rect 97632 18572 97684 18624
rect 147128 18572 147180 18624
rect 161204 18572 161256 18624
rect 401600 18572 401652 18624
rect 122472 18504 122524 18556
rect 247040 18504 247092 18556
rect 115572 18436 115624 18488
rect 220820 18436 220872 18488
rect 126520 17892 126572 17944
rect 262220 17892 262272 17944
rect 127900 17824 127952 17876
rect 266360 17824 266412 17876
rect 127992 17756 128044 17808
rect 269120 17756 269172 17808
rect 129372 17688 129424 17740
rect 273260 17688 273312 17740
rect 130752 17620 130804 17672
rect 280160 17620 280212 17672
rect 166264 17552 166316 17604
rect 318800 17552 318852 17604
rect 170404 17484 170456 17536
rect 325700 17484 325752 17536
rect 142988 17416 143040 17468
rect 300860 17416 300912 17468
rect 146944 17348 146996 17400
rect 307760 17348 307812 17400
rect 97724 17280 97776 17332
rect 119344 17280 119396 17332
rect 144736 17280 144788 17332
rect 332692 17280 332744 17332
rect 94872 17212 94924 17264
rect 122104 17212 122156 17264
rect 209044 17212 209096 17264
rect 415492 17212 415544 17264
rect 125416 17144 125468 17196
rect 259460 17144 259512 17196
rect 125324 17076 125376 17128
rect 255320 17076 255372 17128
rect 142896 17008 142948 17060
rect 242900 17008 242952 17060
rect 119804 16532 119856 16584
rect 238116 16532 238168 16584
rect 121184 16464 121236 16516
rect 241704 16464 241756 16516
rect 122564 16396 122616 16448
rect 245200 16396 245252 16448
rect 122656 16328 122708 16380
rect 248788 16328 248840 16380
rect 123944 16260 123996 16312
rect 252376 16260 252428 16312
rect 201132 16192 201184 16244
rect 560852 16192 560904 16244
rect 202420 16124 202472 16176
rect 564440 16124 564492 16176
rect 203892 16056 203944 16108
rect 568028 16056 568080 16108
rect 99012 15988 99064 16040
rect 116584 15988 116636 16040
rect 203984 15988 204036 16040
rect 571524 15988 571576 16040
rect 94964 15920 95016 15972
rect 115204 15920 115256 15972
rect 205180 15920 205232 15972
rect 575112 15920 575164 15972
rect 112996 15852 113048 15904
rect 206192 15852 206244 15904
rect 206744 15852 206796 15904
rect 578608 15852 578660 15904
rect 119896 15784 119948 15836
rect 234620 15784 234672 15836
rect 118608 15716 118660 15768
rect 231032 15716 231084 15768
rect 117044 15648 117096 15700
rect 226340 15648 226392 15700
rect 116952 15580 117004 15632
rect 223948 15580 224000 15632
rect 115756 15512 115808 15564
rect 220452 15512 220504 15564
rect 115664 15444 115716 15496
rect 216864 15444 216916 15496
rect 114284 15376 114336 15428
rect 213368 15376 213420 15428
rect 112904 15308 112956 15360
rect 209872 15308 209924 15360
rect 183192 15104 183244 15156
rect 489920 15104 489972 15156
rect 184756 15036 184808 15088
rect 493508 15036 493560 15088
rect 185952 14968 186004 15020
rect 497096 14968 497148 15020
rect 186044 14900 186096 14952
rect 500592 14900 500644 14952
rect 187332 14832 187384 14884
rect 504180 14832 504232 14884
rect 188896 14764 188948 14816
rect 507676 14764 507728 14816
rect 188712 14696 188764 14748
rect 511264 14696 511316 14748
rect 190184 14628 190236 14680
rect 514760 14628 514812 14680
rect 191564 14560 191616 14612
rect 518348 14560 518400 14612
rect 191472 14492 191524 14544
rect 521844 14492 521896 14544
rect 106004 14424 106056 14476
rect 182548 14424 182600 14476
rect 193036 14424 193088 14476
rect 525432 14424 525484 14476
rect 183284 14356 183336 14408
rect 486424 14356 486476 14408
rect 181996 14288 182048 14340
rect 481640 14288 481692 14340
rect 180524 14220 180576 14272
rect 478144 14220 478196 14272
rect 180616 14152 180668 14204
rect 473360 14152 473412 14204
rect 179052 14084 179104 14136
rect 471060 14084 471112 14136
rect 177764 14016 177816 14068
rect 467472 14016 467524 14068
rect 177672 13948 177724 14000
rect 463976 13948 464028 14000
rect 176292 13880 176344 13932
rect 460388 13880 460440 13932
rect 158536 13744 158588 13796
rect 389456 13744 389508 13796
rect 159824 13676 159876 13728
rect 393044 13676 393096 13728
rect 159732 13608 159784 13660
rect 396540 13608 396592 13660
rect 161296 13540 161348 13592
rect 398840 13540 398892 13592
rect 162584 13472 162636 13524
rect 403624 13472 403676 13524
rect 162676 13404 162728 13456
rect 407212 13404 407264 13456
rect 163964 13336 164016 13388
rect 410800 13336 410852 13388
rect 165252 13268 165304 13320
rect 414296 13268 414348 13320
rect 165436 13200 165488 13252
rect 417884 13200 417936 13252
rect 166908 13132 166960 13184
rect 421380 13132 421432 13184
rect 168196 13064 168248 13116
rect 423772 13064 423824 13116
rect 157064 12996 157116 13048
rect 385960 12996 386012 13048
rect 156972 12928 157024 12980
rect 382372 12928 382424 12980
rect 155776 12860 155828 12912
rect 378876 12860 378928 12912
rect 154212 12792 154264 12844
rect 374000 12792 374052 12844
rect 154304 12724 154356 12776
rect 371700 12724 371752 12776
rect 152924 12656 152976 12708
rect 368204 12656 368256 12708
rect 153016 12588 153068 12640
rect 364616 12588 364668 12640
rect 151544 12520 151596 12572
rect 361120 12520 361172 12572
rect 133604 12384 133656 12436
rect 290188 12384 290240 12436
rect 135076 12316 135128 12368
rect 293684 12316 293736 12368
rect 134984 12248 135036 12300
rect 297272 12248 297324 12300
rect 136456 12180 136508 12232
rect 299480 12180 299532 12232
rect 137836 12112 137888 12164
rect 304356 12112 304408 12164
rect 137744 12044 137796 12096
rect 307944 12044 307996 12096
rect 139124 11976 139176 12028
rect 311440 11976 311492 12028
rect 139216 11908 139268 11960
rect 315028 11908 315080 11960
rect 140688 11840 140740 11892
rect 318524 11840 318576 11892
rect 141976 11772 142028 11824
rect 322112 11772 322164 11824
rect 141792 11704 141844 11756
rect 325608 11704 325660 11756
rect 357532 11704 357584 11756
rect 358728 11704 358780 11756
rect 432052 11704 432104 11756
rect 433248 11704 433300 11756
rect 132316 11636 132368 11688
rect 286600 11636 286652 11688
rect 132224 11568 132276 11620
rect 283104 11568 283156 11620
rect 130844 11500 130896 11552
rect 279516 11500 279568 11552
rect 129464 11432 129516 11484
rect 276112 11432 276164 11484
rect 129556 11364 129608 11416
rect 272432 11364 272484 11416
rect 128084 11296 128136 11348
rect 268844 11296 268896 11348
rect 126612 11228 126664 11280
rect 265348 11228 265400 11280
rect 126704 11160 126756 11212
rect 261760 11160 261812 11212
rect 107292 10956 107344 11008
rect 187332 10956 187384 11008
rect 197084 10956 197136 11008
rect 541992 10956 542044 11008
rect 107384 10888 107436 10940
rect 188528 10888 188580 10940
rect 198464 10888 198516 10940
rect 545488 10888 545540 10940
rect 108672 10820 108724 10872
rect 190828 10820 190880 10872
rect 198556 10820 198608 10872
rect 547880 10820 547932 10872
rect 108764 10752 108816 10804
rect 192024 10752 192076 10804
rect 199844 10752 199896 10804
rect 552664 10752 552716 10804
rect 110236 10684 110288 10736
rect 195612 10684 195664 10736
rect 201224 10684 201276 10736
rect 556160 10684 556212 10736
rect 108580 10616 108632 10668
rect 193220 10616 193272 10668
rect 201316 10616 201368 10668
rect 559748 10616 559800 10668
rect 110144 10548 110196 10600
rect 197912 10548 197964 10600
rect 202512 10548 202564 10600
rect 202604 10548 202656 10600
rect 563244 10548 563296 10600
rect 110052 10480 110104 10532
rect 199108 10480 199160 10532
rect 566832 10480 566884 10532
rect 111524 10412 111576 10464
rect 202512 10412 202564 10464
rect 204076 10412 204128 10464
rect 570328 10412 570380 10464
rect 111432 10344 111484 10396
rect 201500 10344 201552 10396
rect 205364 10344 205416 10396
rect 572720 10344 572772 10396
rect 88156 10276 88208 10328
rect 106924 10276 106976 10328
rect 111340 10276 111392 10328
rect 205088 10276 205140 10328
rect 205272 10276 205324 10328
rect 577412 10276 577464 10328
rect 195796 10208 195848 10260
rect 538404 10208 538456 10260
rect 195704 10140 195756 10192
rect 534908 10140 534960 10192
rect 114376 10072 114428 10124
rect 215668 10072 215720 10124
rect 215944 10072 215996 10124
rect 372896 10072 372948 10124
rect 117136 10004 117188 10056
rect 226432 10004 226484 10056
rect 116860 9936 116912 9988
rect 222752 9936 222804 9988
rect 115480 9868 115532 9920
rect 219256 9868 219308 9920
rect 114468 9800 114520 9852
rect 212172 9800 212224 9852
rect 112812 9732 112864 9784
rect 208584 9732 208636 9784
rect 176384 9596 176436 9648
rect 462780 9596 462832 9648
rect 101864 9528 101916 9580
rect 163688 9528 163740 9580
rect 177856 9528 177908 9580
rect 466276 9528 466328 9580
rect 101772 9460 101824 9512
rect 167184 9460 167236 9512
rect 179236 9460 179288 9512
rect 469864 9460 469916 9512
rect 103336 9392 103388 9444
rect 170772 9392 170824 9444
rect 179144 9392 179196 9444
rect 473452 9392 473504 9444
rect 104716 9324 104768 9376
rect 174268 9324 174320 9376
rect 180708 9324 180760 9376
rect 476948 9324 477000 9376
rect 104624 9256 104676 9308
rect 177856 9256 177908 9308
rect 181904 9256 181956 9308
rect 481732 9256 481784 9308
rect 104532 9188 104584 9240
rect 176660 9188 176712 9240
rect 183376 9188 183428 9240
rect 485228 9188 485280 9240
rect 106188 9120 106240 9172
rect 180248 9120 180300 9172
rect 183100 9120 183152 9172
rect 488816 9120 488868 9172
rect 106096 9052 106148 9104
rect 181444 9052 181496 9104
rect 184664 9052 184716 9104
rect 492312 9052 492364 9104
rect 107568 8984 107620 9036
rect 183744 8984 183796 9036
rect 185860 8984 185912 9036
rect 495900 8984 495952 9036
rect 107476 8916 107528 8968
rect 184940 8916 184992 8968
rect 186136 8916 186188 8968
rect 499396 8916 499448 8968
rect 176476 8848 176528 8900
rect 459192 8848 459244 8900
rect 175188 8780 175240 8832
rect 455696 8780 455748 8832
rect 175096 8712 175148 8764
rect 452108 8712 452160 8764
rect 173808 8644 173860 8696
rect 448612 8644 448664 8696
rect 172336 8576 172388 8628
rect 445024 8576 445076 8628
rect 172244 8508 172296 8560
rect 441528 8508 441580 8560
rect 171048 8440 171100 8492
rect 437940 8440 437992 8492
rect 169668 8372 169720 8424
rect 434444 8372 434496 8424
rect 151636 8236 151688 8288
rect 363512 8236 363564 8288
rect 153108 8168 153160 8220
rect 367008 8168 367060 8220
rect 154488 8100 154540 8152
rect 370596 8100 370648 8152
rect 154396 8032 154448 8084
rect 374092 8032 374144 8084
rect 155592 7964 155644 8016
rect 377680 7964 377732 8016
rect 157156 7896 157208 7948
rect 381176 7896 381228 7948
rect 95056 7828 95108 7880
rect 137652 7828 137704 7880
rect 157248 7828 157300 7880
rect 384764 7828 384816 7880
rect 96344 7760 96396 7812
rect 141240 7760 141292 7812
rect 158628 7760 158680 7812
rect 388260 7760 388312 7812
rect 99104 7692 99156 7744
rect 151820 7692 151872 7744
rect 159640 7692 159692 7744
rect 391848 7692 391900 7744
rect 99196 7624 99248 7676
rect 155408 7624 155460 7676
rect 159916 7624 159968 7676
rect 395344 7624 395396 7676
rect 100484 7556 100536 7608
rect 158904 7556 158956 7608
rect 161388 7556 161440 7608
rect 398932 7556 398984 7608
rect 151728 7488 151780 7540
rect 359924 7488 359976 7540
rect 150348 7420 150400 7472
rect 356336 7420 356388 7472
rect 148876 7352 148928 7404
rect 352840 7352 352892 7404
rect 148968 7284 149020 7336
rect 349252 7284 349304 7336
rect 147588 7216 147640 7268
rect 345756 7216 345808 7268
rect 146116 7148 146168 7200
rect 342168 7148 342220 7200
rect 146208 7080 146260 7132
rect 338672 7080 338724 7132
rect 144828 7012 144880 7064
rect 335084 7012 335136 7064
rect 126796 6808 126848 6860
rect 264152 6808 264204 6860
rect 128176 6740 128228 6792
rect 267740 6740 267792 6792
rect 128268 6672 128320 6724
rect 271236 6672 271288 6724
rect 129648 6604 129700 6656
rect 274824 6604 274876 6656
rect 130936 6536 130988 6588
rect 278320 6536 278372 6588
rect 131028 6468 131080 6520
rect 281908 6468 281960 6520
rect 132408 6400 132460 6452
rect 285404 6400 285456 6452
rect 133696 6332 133748 6384
rect 288992 6332 289044 6384
rect 105636 6264 105688 6316
rect 128176 6264 128228 6316
rect 133788 6264 133840 6316
rect 292580 6264 292632 6316
rect 93584 6196 93636 6248
rect 130568 6196 130620 6248
rect 135168 6196 135220 6248
rect 296076 6196 296128 6248
rect 93492 6128 93544 6180
rect 134156 6128 134208 6180
rect 136548 6128 136600 6180
rect 299664 6128 299716 6180
rect 126888 6060 126940 6112
rect 260656 6060 260708 6112
rect 125232 5992 125284 6044
rect 257068 5992 257120 6044
rect 123760 5924 123812 5976
rect 253480 5924 253532 5976
rect 124036 5856 124088 5908
rect 249984 5856 250036 5908
rect 122748 5788 122800 5840
rect 246396 5788 246448 5840
rect 121368 5720 121420 5772
rect 242992 5720 243044 5772
rect 121276 5652 121328 5704
rect 239312 5652 239364 5704
rect 119620 5584 119672 5636
rect 235816 5584 235868 5636
rect 99288 5448 99340 5500
rect 154212 5448 154264 5500
rect 196900 5448 196952 5500
rect 540796 5448 540848 5500
rect 100576 5380 100628 5432
rect 157800 5380 157852 5432
rect 197176 5380 197228 5432
rect 544292 5380 544344 5432
rect 102048 5312 102100 5364
rect 162492 5312 162544 5364
rect 198280 5312 198332 5364
rect 547972 5312 548024 5364
rect 101956 5244 102008 5296
rect 166080 5244 166132 5296
rect 199936 5244 199988 5296
rect 551468 5244 551520 5296
rect 103428 5176 103480 5228
rect 169576 5176 169628 5228
rect 200028 5176 200080 5228
rect 554964 5176 555016 5228
rect 104808 5108 104860 5160
rect 173164 5108 173216 5160
rect 202604 5108 202656 5160
rect 558552 5108 558604 5160
rect 108948 5040 109000 5092
rect 189724 5040 189776 5092
rect 202788 5040 202840 5092
rect 562048 5040 562100 5092
rect 108856 4972 108908 5024
rect 193312 4972 193364 5024
rect 194140 4972 194192 5024
rect 565636 4972 565688 5024
rect 110328 4904 110380 4956
rect 196808 4904 196860 4956
rect 204168 4904 204220 4956
rect 569132 4904 569184 4956
rect 111708 4836 111760 4888
rect 201040 4836 201092 4888
rect 205548 4836 205600 4888
rect 572812 4836 572864 4888
rect 62028 4768 62080 4820
rect 71044 4768 71096 4820
rect 111616 4768 111668 4820
rect 203892 4768 203944 4820
rect 205456 4768 205508 4820
rect 576308 4768 576360 4820
rect 97816 4700 97868 4752
rect 150624 4700 150676 4752
rect 200304 4700 200356 4752
rect 93400 4632 93452 4684
rect 132960 4632 133012 4684
rect 133144 4632 133196 4684
rect 186136 4632 186188 4684
rect 195888 4632 195940 4684
rect 537208 4700 537260 4752
rect 533712 4632 533764 4684
rect 97908 4564 97960 4616
rect 147036 4564 147088 4616
rect 148324 4564 148376 4616
rect 175464 4564 175516 4616
rect 194508 4564 194560 4616
rect 530124 4564 530176 4616
rect 96436 4496 96488 4548
rect 143540 4496 143592 4548
rect 192852 4496 192904 4548
rect 526628 4496 526680 4548
rect 96528 4428 96580 4480
rect 140044 4428 140096 4480
rect 140136 4428 140188 4480
rect 179052 4428 179104 4480
rect 191656 4428 191708 4480
rect 523040 4428 523092 4480
rect 95148 4360 95200 4412
rect 136456 4360 136508 4412
rect 191380 4360 191432 4412
rect 519544 4360 519596 4412
rect 92296 4292 92348 4344
rect 126980 4292 127032 4344
rect 190276 4292 190328 4344
rect 515956 4292 516008 4344
rect 93676 4224 93728 4276
rect 129372 4224 129424 4276
rect 190092 4224 190144 4276
rect 512460 4224 512512 4276
rect 43076 4088 43128 4140
rect 38384 4020 38436 4072
rect 87696 4156 87748 4208
rect 90364 4156 90416 4208
rect 98644 4156 98696 4208
rect 101036 4156 101088 4208
rect 105544 4156 105596 4208
rect 108120 4156 108172 4208
rect 64144 4088 64196 4140
rect 65524 4088 65576 4140
rect 89444 4088 89496 4140
rect 67088 4020 67140 4072
rect 89536 4020 89588 4072
rect 112444 4088 112496 4140
rect 131764 4088 131816 4140
rect 141424 4088 141476 4140
rect 144736 4088 144788 4140
rect 222844 4088 222896 4140
rect 112812 4020 112864 4072
rect 115204 4020 115256 4072
rect 138848 4020 138900 4072
rect 209780 4020 209832 4072
rect 210976 4020 211028 4072
rect 226340 4020 226392 4072
rect 227536 4020 227588 4072
rect 276020 4088 276072 4140
rect 277124 4088 277176 4140
rect 387064 4088 387116 4140
rect 479340 4088 479392 4140
rect 379980 4020 380032 4072
rect 391204 4020 391256 4072
rect 582196 4020 582248 4072
rect 35992 3952 36044 4004
rect 12348 3884 12400 3936
rect 29644 3884 29696 3936
rect 31300 3884 31352 3936
rect 28816 3816 28868 3868
rect 1676 3748 1728 3800
rect 21364 3748 21416 3800
rect 23020 3748 23072 3800
rect 60832 3952 60884 4004
rect 64328 3952 64380 4004
rect 90916 3952 90968 4004
rect 119896 3952 119948 4004
rect 168104 3952 168156 4004
rect 429660 3952 429712 4004
rect 436836 3952 436888 4004
rect 442632 3952 442684 4004
rect 447784 3952 447836 4004
rect 63684 3884 63736 3936
rect 63776 3884 63828 3936
rect 89628 3884 89680 3936
rect 117596 3884 117648 3936
rect 144184 3884 144236 3936
rect 161296 3884 161348 3936
rect 174544 3884 174596 3936
rect 436744 3884 436796 3936
rect 64328 3816 64380 3868
rect 66996 3816 67048 3868
rect 82544 3816 82596 3868
rect 85672 3816 85724 3868
rect 90732 3816 90784 3868
rect 118792 3816 118844 3868
rect 119344 3816 119396 3868
rect 145932 3816 145984 3868
rect 172152 3816 172204 3868
rect 443828 3816 443880 3868
rect 450544 3816 450596 3868
rect 479524 3952 479576 4004
rect 505376 3952 505428 4004
rect 454684 3884 454736 3936
rect 480536 3884 480588 3936
rect 19432 3680 19484 3732
rect 66904 3748 66956 3800
rect 90824 3748 90876 3800
rect 121092 3748 121144 3800
rect 122104 3748 122156 3800
rect 62948 3680 63000 3732
rect 91008 3680 91060 3732
rect 122288 3680 122340 3732
rect 129004 3748 129056 3800
rect 148324 3748 148376 3800
rect 175924 3748 175976 3800
rect 450912 3748 450964 3800
rect 510068 3816 510120 3868
rect 506480 3748 506532 3800
rect 135260 3680 135312 3732
rect 142804 3680 142856 3732
rect 171968 3680 172020 3732
rect 176568 3680 176620 3732
rect 458088 3680 458140 3732
rect 461676 3680 461728 3732
rect 487620 3680 487672 3732
rect 544384 3680 544436 3732
rect 557356 3680 557408 3732
rect 8760 3612 8812 3664
rect 9956 3544 10008 3596
rect 10968 3544 11020 3596
rect 11152 3612 11204 3664
rect 62488 3612 62540 3664
rect 84016 3612 84068 3664
rect 91560 3612 91612 3664
rect 92388 3612 92440 3664
rect 124680 3612 124732 3664
rect 134524 3612 134576 3664
rect 164884 3612 164936 3664
rect 177948 3612 178000 3664
rect 465172 3612 465224 3664
rect 472624 3612 472676 3664
rect 485044 3612 485096 3664
rect 517152 3612 517204 3664
rect 62120 3544 62172 3596
rect 5264 3476 5316 3528
rect 572 3408 624 3460
rect 11704 3408 11756 3460
rect 15936 3408 15988 3460
rect 16488 3408 16540 3460
rect 17040 3408 17092 3460
rect 17868 3408 17920 3460
rect 18236 3408 18288 3460
rect 19248 3408 19300 3460
rect 21824 3408 21876 3460
rect 22836 3408 22888 3460
rect 24216 3408 24268 3460
rect 24768 3408 24820 3460
rect 25320 3408 25372 3460
rect 26148 3408 26200 3460
rect 26516 3408 26568 3460
rect 27528 3408 27580 3460
rect 27712 3408 27764 3460
rect 28908 3408 28960 3460
rect 32404 3408 32456 3460
rect 33048 3408 33100 3460
rect 33600 3408 33652 3460
rect 34428 3408 34480 3460
rect 34796 3408 34848 3460
rect 35808 3408 35860 3460
rect 40684 3408 40736 3460
rect 41328 3408 41380 3460
rect 41880 3408 41932 3460
rect 43444 3408 43496 3460
rect 46664 3408 46716 3460
rect 50344 3408 50396 3460
rect 51356 3408 51408 3460
rect 52368 3408 52420 3460
rect 45468 3340 45520 3392
rect 58440 3476 58492 3528
rect 59268 3476 59320 3528
rect 64144 3544 64196 3596
rect 81348 3544 81400 3596
rect 63224 3476 63276 3528
rect 74724 3476 74776 3528
rect 75000 3476 75052 3528
rect 75828 3476 75880 3528
rect 76196 3476 76248 3528
rect 77208 3476 77260 3528
rect 80336 3476 80388 3528
rect 80888 3476 80940 3528
rect 81256 3476 81308 3528
rect 82084 3476 82136 3528
rect 83464 3544 83516 3596
rect 87972 3544 88024 3596
rect 90640 3544 90692 3596
rect 123484 3544 123536 3596
rect 124864 3544 124916 3596
rect 125876 3544 125928 3596
rect 137284 3544 137336 3596
rect 168380 3544 168432 3596
rect 179328 3544 179380 3596
rect 472256 3544 472308 3596
rect 473360 3544 473412 3596
rect 474556 3544 474608 3596
rect 481640 3544 481692 3596
rect 482836 3544 482888 3596
rect 489184 3544 489236 3596
rect 532516 3612 532568 3664
rect 537484 3612 537536 3664
rect 553768 3612 553820 3664
rect 530584 3544 530636 3596
rect 531320 3544 531372 3596
rect 533344 3544 533396 3596
rect 550272 3544 550324 3596
rect 572720 3544 572772 3596
rect 573916 3544 573968 3596
rect 84476 3476 84528 3528
rect 85488 3476 85540 3528
rect 66444 3408 66496 3460
rect 66720 3408 66772 3460
rect 67548 3408 67600 3460
rect 67916 3408 67968 3460
rect 68928 3408 68980 3460
rect 69112 3408 69164 3460
rect 70216 3408 70268 3460
rect 72608 3408 72660 3460
rect 73068 3408 73120 3460
rect 73804 3408 73856 3460
rect 75184 3408 75236 3460
rect 77392 3408 77444 3460
rect 78956 3408 79008 3460
rect 79692 3408 79744 3460
rect 80428 3408 80480 3460
rect 82636 3408 82688 3460
rect 89168 3408 89220 3460
rect 89352 3476 89404 3528
rect 116400 3476 116452 3528
rect 116584 3476 116636 3528
rect 153016 3476 153068 3528
rect 193220 3476 193272 3528
rect 194416 3476 194468 3528
rect 206928 3476 206980 3528
rect 581000 3476 581052 3528
rect 99840 3408 99892 3460
rect 100392 3408 100444 3460
rect 61016 3340 61068 3392
rect 65524 3340 65576 3392
rect 76104 3340 76156 3392
rect 88248 3340 88300 3392
rect 109316 3340 109368 3392
rect 147128 3408 147180 3460
rect 149520 3408 149572 3460
rect 152464 3408 152516 3460
rect 156604 3408 156656 3460
rect 206836 3408 206888 3460
rect 583392 3408 583444 3460
rect 160100 3340 160152 3392
rect 242900 3340 242952 3392
rect 244096 3340 244148 3392
rect 307760 3340 307812 3392
rect 309048 3340 309100 3392
rect 316040 3340 316092 3392
rect 317328 3340 317380 3392
rect 332600 3340 332652 3392
rect 333888 3340 333940 3392
rect 349160 3340 349212 3392
rect 350448 3340 350500 3392
rect 374000 3340 374052 3392
rect 375288 3340 375340 3392
rect 382924 3340 382976 3392
rect 475752 3340 475804 3392
rect 44272 3272 44324 3324
rect 50160 3204 50212 3256
rect 64420 3272 64472 3324
rect 86684 3272 86736 3324
rect 105728 3272 105780 3324
rect 106924 3272 106976 3324
rect 111616 3272 111668 3324
rect 115204 3272 115256 3324
rect 382280 3272 382332 3324
rect 383568 3272 383620 3324
rect 398840 3272 398892 3324
rect 400128 3272 400180 3324
rect 407764 3272 407816 3324
rect 409604 3272 409656 3324
rect 414664 3272 414716 3324
rect 416688 3272 416740 3324
rect 423772 3272 423824 3324
rect 424968 3272 425020 3324
rect 475384 3272 475436 3324
rect 498200 3340 498252 3392
rect 512644 3340 512696 3392
rect 513564 3340 513616 3392
rect 526444 3340 526496 3392
rect 527824 3340 527876 3392
rect 547880 3340 547932 3392
rect 549076 3340 549128 3392
rect 494704 3272 494756 3324
rect 62856 3204 62908 3256
rect 86776 3204 86828 3256
rect 102232 3204 102284 3256
rect 102876 3204 102928 3256
rect 114008 3204 114060 3256
rect 388444 3204 388496 3256
rect 390652 3204 390704 3256
rect 407120 3204 407172 3256
rect 408408 3204 408460 3256
rect 418804 3204 418856 3256
rect 420184 3204 420236 3256
rect 468484 3204 468536 3256
rect 491116 3204 491168 3256
rect 519636 3204 519688 3256
rect 524236 3204 524288 3256
rect 56048 3136 56100 3188
rect 68284 3136 68336 3188
rect 87604 3136 87656 3188
rect 98644 3136 98696 3188
rect 102784 3136 102836 3188
rect 110512 3136 110564 3188
rect 396724 3136 396776 3188
rect 397736 3136 397788 3188
rect 443644 3136 443696 3188
rect 449808 3136 449860 3188
rect 52552 3068 52604 3120
rect 62764 3068 62816 3120
rect 86868 3068 86920 3120
rect 103336 3068 103388 3120
rect 2872 3000 2924 3052
rect 4804 3000 4856 3052
rect 48964 3000 49016 3052
rect 57152 3000 57204 3052
rect 57244 3000 57296 3052
rect 65616 3000 65668 3052
rect 84108 3000 84160 3052
rect 95148 3000 95200 3052
rect 101404 3000 101456 3052
rect 106924 3000 106976 3052
rect 425796 3000 425848 3052
rect 427268 3000 427320 3052
rect 59636 2932 59688 2984
rect 68376 2932 68428 2984
rect 86224 2932 86276 2984
rect 96252 2932 96304 2984
rect 7656 2864 7708 2916
rect 8208 2864 8260 2916
rect 63776 2864 63828 2916
rect 82728 2864 82780 2916
rect 86868 2864 86920 2916
rect 421564 2864 421616 2916
rect 423772 2864 423824 2916
rect 20628 2796 20680 2848
rect 65064 2796 65116 2848
rect 83924 2796 83976 2848
rect 92756 2796 92808 2848
rect 299480 1640 299532 1692
rect 300768 1640 300820 1692
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 412652 703582 413508 703610
rect 8128 702434 8156 703520
rect 8128 702406 8248 702434
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3436 683194 3464 684247
rect 3424 683188 3476 683194
rect 3424 683130 3476 683136
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3528 670750 3556 671191
rect 3516 670744 3568 670750
rect 3516 670686 3568 670692
rect 3422 658200 3478 658209
rect 3422 658135 3478 658144
rect 3436 656946 3464 658135
rect 3424 656940 3476 656946
rect 3424 656882 3476 656888
rect 3424 632120 3476 632126
rect 3422 632088 3424 632097
rect 3476 632088 3478 632097
rect 3422 632023 3478 632032
rect 3146 619168 3202 619177
rect 3146 619103 3202 619112
rect 3160 618322 3188 619103
rect 3148 618316 3200 618322
rect 3148 618258 3200 618264
rect 3238 606112 3294 606121
rect 3238 606047 3294 606056
rect 3252 605878 3280 606047
rect 3240 605872 3292 605878
rect 3240 605814 3292 605820
rect 3330 580000 3386 580009
rect 3330 579935 3386 579944
rect 3344 579698 3372 579935
rect 3332 579692 3384 579698
rect 3332 579634 3384 579640
rect 3422 566944 3478 566953
rect 3422 566879 3478 566888
rect 3436 565894 3464 566879
rect 3424 565888 3476 565894
rect 3424 565830 3476 565836
rect 3422 553888 3478 553897
rect 3422 553823 3478 553832
rect 3436 553450 3464 553823
rect 3424 553444 3476 553450
rect 3424 553386 3476 553392
rect 3422 527912 3478 527921
rect 3422 527847 3478 527856
rect 3436 527202 3464 527847
rect 3424 527196 3476 527202
rect 3424 527138 3476 527144
rect 3422 514856 3478 514865
rect 3422 514791 3424 514800
rect 3476 514791 3478 514800
rect 3424 514762 3476 514768
rect 2778 501800 2834 501809
rect 2778 501735 2834 501744
rect 2792 501090 2820 501735
rect 2780 501084 2832 501090
rect 2780 501026 2832 501032
rect 4804 501084 4856 501090
rect 4804 501026 4856 501032
rect 3422 475688 3478 475697
rect 3422 475623 3478 475632
rect 3436 474774 3464 475623
rect 3424 474768 3476 474774
rect 3424 474710 3476 474716
rect 3238 462632 3294 462641
rect 3238 462567 3294 462576
rect 3252 462398 3280 462567
rect 3240 462392 3292 462398
rect 3240 462334 3292 462340
rect 3146 449576 3202 449585
rect 3146 449511 3202 449520
rect 3160 448594 3188 449511
rect 3148 448588 3200 448594
rect 3148 448530 3200 448536
rect 3422 423600 3478 423609
rect 3422 423535 3478 423544
rect 3436 422346 3464 423535
rect 3424 422340 3476 422346
rect 3424 422282 3476 422288
rect 3146 410544 3202 410553
rect 3146 410479 3202 410488
rect 3160 409902 3188 410479
rect 3148 409896 3200 409902
rect 3148 409838 3200 409844
rect 3424 397520 3476 397526
rect 3422 397488 3424 397497
rect 3476 397488 3478 397497
rect 3422 397423 3478 397432
rect 3422 371376 3478 371385
rect 3422 371311 3478 371320
rect 3436 371278 3464 371311
rect 3424 371272 3476 371278
rect 3424 371214 3476 371220
rect 3146 358456 3202 358465
rect 3146 358391 3202 358400
rect 3160 357474 3188 358391
rect 3148 357468 3200 357474
rect 3148 357410 3200 357416
rect 3330 345400 3386 345409
rect 3330 345335 3386 345344
rect 3344 345098 3372 345335
rect 3332 345092 3384 345098
rect 3332 345034 3384 345040
rect 3422 319288 3478 319297
rect 3422 319223 3478 319232
rect 3436 318850 3464 319223
rect 3424 318844 3476 318850
rect 3424 318786 3476 318792
rect 3238 306232 3294 306241
rect 3238 306167 3294 306176
rect 3252 305046 3280 306167
rect 3240 305040 3292 305046
rect 3240 304982 3292 304988
rect 3422 293176 3478 293185
rect 3422 293111 3478 293120
rect 3436 292602 3464 293111
rect 3424 292596 3476 292602
rect 3424 292538 3476 292544
rect 3054 267200 3110 267209
rect 3054 267135 3110 267144
rect 3068 266422 3096 267135
rect 3056 266416 3108 266422
rect 3056 266358 3108 266364
rect 3422 254144 3478 254153
rect 3422 254079 3478 254088
rect 3436 253978 3464 254079
rect 3424 253972 3476 253978
rect 3424 253914 3476 253920
rect 4816 245342 4844 501026
rect 8220 245546 8248 702406
rect 24320 700330 24348 703520
rect 40512 700398 40540 703520
rect 40500 700392 40552 700398
rect 40500 700334 40552 700340
rect 41328 700392 41380 700398
rect 41328 700334 41380 700340
rect 24308 700324 24360 700330
rect 24308 700266 24360 700272
rect 33784 700324 33836 700330
rect 33784 700266 33836 700272
rect 11704 683188 11756 683194
rect 11704 683130 11756 683136
rect 8208 245540 8260 245546
rect 8208 245482 8260 245488
rect 4804 245336 4856 245342
rect 4804 245278 4856 245284
rect 11716 244254 11744 683130
rect 22744 656940 22796 656946
rect 22744 656882 22796 656888
rect 14464 632120 14516 632126
rect 14464 632062 14516 632068
rect 11704 244248 11756 244254
rect 11704 244190 11756 244196
rect 14476 242554 14504 632062
rect 21364 579692 21416 579698
rect 21364 579634 21416 579640
rect 15844 527196 15896 527202
rect 15844 527138 15896 527144
rect 15856 244186 15884 527138
rect 17224 474768 17276 474774
rect 17224 474710 17276 474716
rect 15844 244180 15896 244186
rect 15844 244122 15896 244128
rect 17236 244118 17264 474710
rect 18604 422340 18656 422346
rect 18604 422282 18656 422288
rect 18616 245410 18644 422282
rect 18604 245404 18656 245410
rect 18604 245346 18656 245352
rect 17224 244112 17276 244118
rect 17224 244054 17276 244060
rect 21376 243506 21404 579634
rect 22756 245614 22784 656882
rect 25504 605872 25556 605878
rect 25504 605814 25556 605820
rect 22744 245608 22796 245614
rect 22744 245550 22796 245556
rect 25516 244866 25544 605814
rect 29644 553444 29696 553450
rect 29644 553386 29696 553392
rect 25504 244860 25556 244866
rect 25504 244802 25556 244808
rect 29656 244798 29684 553386
rect 32404 448588 32456 448594
rect 32404 448530 32456 448536
rect 32416 247042 32444 448530
rect 32404 247036 32456 247042
rect 32404 246978 32456 246984
rect 33796 246226 33824 700266
rect 36544 670744 36596 670750
rect 36544 670686 36596 670692
rect 35164 618316 35216 618322
rect 35164 618258 35216 618264
rect 35176 246294 35204 618258
rect 35164 246288 35216 246294
rect 35164 246230 35216 246236
rect 33784 246220 33836 246226
rect 33784 246162 33836 246168
rect 36556 246158 36584 670686
rect 39304 565888 39356 565894
rect 39304 565830 39356 565836
rect 36544 246152 36596 246158
rect 36544 246094 36596 246100
rect 29644 244792 29696 244798
rect 29644 244734 29696 244740
rect 21364 243500 21416 243506
rect 21364 243442 21416 243448
rect 39316 243234 39344 565830
rect 39304 243228 39356 243234
rect 39304 243170 39356 243176
rect 41340 243166 41368 700334
rect 72988 700330 73016 703520
rect 59268 700324 59320 700330
rect 59268 700266 59320 700272
rect 72976 700324 73028 700330
rect 72976 700266 73028 700272
rect 43444 514820 43496 514826
rect 43444 514762 43496 514768
rect 43456 244594 43484 514762
rect 56508 505096 56560 505102
rect 56508 505038 56560 505044
rect 53288 504960 53340 504966
rect 53288 504902 53340 504908
rect 52366 504248 52422 504257
rect 52276 504212 52328 504218
rect 52366 504183 52422 504192
rect 52276 504154 52328 504160
rect 50986 504112 51042 504121
rect 50804 504076 50856 504082
rect 50986 504047 51042 504056
rect 50804 504018 50856 504024
rect 50620 503940 50672 503946
rect 50620 503882 50672 503888
rect 47584 462392 47636 462398
rect 47584 462334 47636 462340
rect 47596 247994 47624 462334
rect 50344 409896 50396 409902
rect 50344 409838 50396 409844
rect 47584 247988 47636 247994
rect 47584 247930 47636 247936
rect 50356 244662 50384 409838
rect 50344 244656 50396 244662
rect 50344 244598 50396 244604
rect 43444 244588 43496 244594
rect 43444 244530 43496 244536
rect 41328 243160 41380 243166
rect 41328 243102 41380 243108
rect 14464 242548 14516 242554
rect 14464 242490 14516 242496
rect 3422 241088 3478 241097
rect 3422 241023 3478 241032
rect 3436 240174 3464 241023
rect 3424 240168 3476 240174
rect 3424 240110 3476 240116
rect 33782 234832 33838 234841
rect 33782 234767 33838 234776
rect 15842 232384 15898 232393
rect 15842 232319 15898 232328
rect 14462 230888 14518 230897
rect 14462 230823 14518 230832
rect 11702 229528 11758 229537
rect 11702 229463 11758 229472
rect 7562 229392 7618 229401
rect 7562 229327 7618 229336
rect 3422 226944 3478 226953
rect 3422 226879 3478 226888
rect 3056 202836 3108 202842
rect 3056 202778 3108 202784
rect 3068 201929 3096 202778
rect 3054 201920 3110 201929
rect 3054 201855 3110 201864
rect 2780 188896 2832 188902
rect 2778 188864 2780 188873
rect 2832 188864 2834 188873
rect 2778 188799 2834 188808
rect 3240 164212 3292 164218
rect 3240 164154 3292 164160
rect 3252 162897 3280 164154
rect 3238 162888 3294 162897
rect 3238 162823 3294 162832
rect 3148 111784 3200 111790
rect 3148 111726 3200 111732
rect 3160 110673 3188 111726
rect 3146 110664 3202 110673
rect 3146 110599 3202 110608
rect 3056 59356 3108 59362
rect 3056 59298 3108 59304
rect 3068 58585 3096 59298
rect 3054 58576 3110 58585
rect 3054 58511 3110 58520
rect 3436 6497 3464 226879
rect 4802 226672 4858 226681
rect 4802 226607 4858 226616
rect 3516 215144 3568 215150
rect 3516 215086 3568 215092
rect 3528 214985 3556 215086
rect 3514 214976 3570 214985
rect 3514 214911 3570 214920
rect 4816 188902 4844 226607
rect 7576 215150 7604 229327
rect 7564 215144 7616 215150
rect 7564 215086 7616 215092
rect 4804 188896 4856 188902
rect 4804 188838 4856 188844
rect 11716 164218 11744 229463
rect 11704 164212 11756 164218
rect 11704 164154 11756 164160
rect 3516 150408 3568 150414
rect 3516 150350 3568 150356
rect 3528 149841 3556 150350
rect 3514 149832 3570 149841
rect 3514 149767 3570 149776
rect 3516 137964 3568 137970
rect 3516 137906 3568 137912
rect 3528 136785 3556 137906
rect 3514 136776 3570 136785
rect 3514 136711 3570 136720
rect 14476 111790 14504 230823
rect 15856 137970 15884 232319
rect 17222 232248 17278 232257
rect 17222 232183 17278 232192
rect 15844 137964 15896 137970
rect 15844 137906 15896 137912
rect 14464 111784 14516 111790
rect 14464 111726 14516 111732
rect 3516 97980 3568 97986
rect 3516 97922 3568 97928
rect 3528 97617 3556 97922
rect 3514 97608 3570 97617
rect 3514 97543 3570 97552
rect 17236 85542 17264 232183
rect 22742 231024 22798 231033
rect 22742 230959 22798 230968
rect 21362 229664 21418 229673
rect 21362 229599 21418 229608
rect 18602 228576 18658 228585
rect 18602 228511 18658 228520
rect 18616 150414 18644 228511
rect 18604 150408 18656 150414
rect 18604 150350 18656 150356
rect 3516 85536 3568 85542
rect 3516 85478 3568 85484
rect 17224 85536 17276 85542
rect 17224 85478 17276 85484
rect 3528 84697 3556 85478
rect 3514 84688 3570 84697
rect 3514 84623 3570 84632
rect 21376 71738 21404 229599
rect 3516 71732 3568 71738
rect 3516 71674 3568 71680
rect 21364 71732 21416 71738
rect 21364 71674 21416 71680
rect 3528 71641 3556 71674
rect 3514 71632 3570 71641
rect 3514 71567 3570 71576
rect 19248 57656 19300 57662
rect 19248 57598 19300 57604
rect 16488 57588 16540 57594
rect 16488 57530 16540 57536
rect 13728 57520 13780 57526
rect 13728 57462 13780 57468
rect 6828 57384 6880 57390
rect 6828 57326 6880 57332
rect 4068 57248 4120 57254
rect 4068 57190 4120 57196
rect 3516 45552 3568 45558
rect 3514 45520 3516 45529
rect 3568 45520 3570 45529
rect 3514 45455 3570 45464
rect 3516 33108 3568 33114
rect 3516 33050 3568 33056
rect 3528 32473 3556 33050
rect 3514 32464 3570 32473
rect 3514 32399 3570 32408
rect 3516 20664 3568 20670
rect 3516 20606 3568 20612
rect 3528 19417 3556 20606
rect 3514 19408 3570 19417
rect 3514 19343 3570 19352
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 1676 3800 1728 3806
rect 1676 3742 1728 3748
rect 572 3460 624 3466
rect 572 3402 624 3408
rect 584 480 612 3402
rect 1688 480 1716 3742
rect 2872 3052 2924 3058
rect 2872 2994 2924 3000
rect 2884 480 2912 2994
rect 4080 480 4108 57190
rect 4804 56024 4856 56030
rect 4804 55966 4856 55972
rect 4816 3058 4844 55966
rect 6840 6914 6868 57326
rect 10968 57316 11020 57322
rect 10968 57258 11020 57264
rect 8208 56092 8260 56098
rect 8208 56034 8260 56040
rect 6472 6886 6868 6914
rect 5264 3528 5316 3534
rect 5264 3470 5316 3476
rect 4804 3052 4856 3058
rect 4804 2994 4856 3000
rect 5276 480 5304 3470
rect 6472 480 6500 6886
rect 8220 2922 8248 56034
rect 8760 3664 8812 3670
rect 8760 3606 8812 3612
rect 7656 2916 7708 2922
rect 7656 2858 7708 2864
rect 8208 2916 8260 2922
rect 8208 2858 8260 2864
rect 7668 480 7696 2858
rect 8772 480 8800 3606
rect 10980 3602 11008 57258
rect 11704 55888 11756 55894
rect 11704 55830 11756 55836
rect 11152 3664 11204 3670
rect 11152 3606 11204 3612
rect 9956 3596 10008 3602
rect 9956 3538 10008 3544
rect 10968 3596 11020 3602
rect 10968 3538 11020 3544
rect 9968 480 9996 3538
rect 11164 480 11192 3606
rect 11716 3466 11744 55830
rect 13740 6914 13768 57462
rect 15108 57452 15160 57458
rect 15108 57394 15160 57400
rect 15120 6914 15148 57394
rect 13556 6886 13768 6914
rect 14752 6886 15148 6914
rect 12348 3936 12400 3942
rect 12348 3878 12400 3884
rect 11704 3460 11756 3466
rect 11704 3402 11756 3408
rect 12360 480 12388 3878
rect 13556 480 13584 6886
rect 14752 480 14780 6886
rect 16500 3466 16528 57530
rect 17868 56160 17920 56166
rect 17868 56102 17920 56108
rect 17880 3466 17908 56102
rect 19260 3466 19288 57598
rect 21364 56364 21416 56370
rect 21364 56306 21416 56312
rect 21376 3806 21404 56306
rect 22756 33114 22784 230959
rect 25502 228032 25558 228041
rect 25502 227967 25558 227976
rect 25516 97986 25544 227967
rect 29642 226808 29698 226817
rect 29642 226743 29698 226752
rect 29656 202842 29684 226743
rect 29644 202836 29696 202842
rect 29644 202778 29696 202784
rect 25504 97980 25556 97986
rect 25504 97922 25556 97928
rect 28908 57860 28960 57866
rect 28908 57802 28960 57808
rect 26148 57792 26200 57798
rect 26148 57734 26200 57740
rect 24768 57724 24820 57730
rect 24768 57666 24820 57672
rect 22836 56228 22888 56234
rect 22836 56170 22888 56176
rect 22744 33108 22796 33114
rect 22744 33050 22796 33056
rect 21364 3800 21416 3806
rect 21364 3742 21416 3748
rect 19432 3732 19484 3738
rect 19432 3674 19484 3680
rect 15936 3460 15988 3466
rect 15936 3402 15988 3408
rect 16488 3460 16540 3466
rect 16488 3402 16540 3408
rect 17040 3460 17092 3466
rect 17040 3402 17092 3408
rect 17868 3460 17920 3466
rect 17868 3402 17920 3408
rect 18236 3460 18288 3466
rect 18236 3402 18288 3408
rect 19248 3460 19300 3466
rect 19248 3402 19300 3408
rect 15948 480 15976 3402
rect 17052 480 17080 3402
rect 18248 480 18276 3402
rect 19444 480 19472 3674
rect 22848 3466 22876 56170
rect 23020 3800 23072 3806
rect 23020 3742 23072 3748
rect 21824 3460 21876 3466
rect 21824 3402 21876 3408
rect 22836 3460 22888 3466
rect 22836 3402 22888 3408
rect 20628 2848 20680 2854
rect 20628 2790 20680 2796
rect 20640 480 20668 2790
rect 21836 480 21864 3402
rect 23032 480 23060 3742
rect 24780 3466 24808 57666
rect 26160 3466 26188 57734
rect 27528 56296 27580 56302
rect 27528 56238 27580 56244
rect 27540 3466 27568 56238
rect 28816 3868 28868 3874
rect 28816 3810 28868 3816
rect 24216 3460 24268 3466
rect 24216 3402 24268 3408
rect 24768 3460 24820 3466
rect 24768 3402 24820 3408
rect 25320 3460 25372 3466
rect 25320 3402 25372 3408
rect 26148 3460 26200 3466
rect 26148 3402 26200 3408
rect 26516 3460 26568 3466
rect 26516 3402 26568 3408
rect 27528 3460 27580 3466
rect 27528 3402 27580 3408
rect 27712 3460 27764 3466
rect 27712 3402 27764 3408
rect 24228 480 24256 3402
rect 25332 480 25360 3402
rect 26528 480 26556 3402
rect 27724 480 27752 3402
rect 28828 1986 28856 3810
rect 28920 3466 28948 57802
rect 33048 57180 33100 57186
rect 33048 57122 33100 57128
rect 29644 56568 29696 56574
rect 29644 56510 29696 56516
rect 29656 3942 29684 56510
rect 30288 56432 30340 56438
rect 30288 56374 30340 56380
rect 30300 6914 30328 56374
rect 30116 6886 30328 6914
rect 29644 3936 29696 3942
rect 29644 3878 29696 3884
rect 28908 3460 28960 3466
rect 28908 3402 28960 3408
rect 28828 1958 28948 1986
rect 28920 480 28948 1958
rect 30116 480 30144 6886
rect 31300 3936 31352 3942
rect 31300 3878 31352 3884
rect 31312 480 31340 3878
rect 33060 3466 33088 57122
rect 33796 20670 33824 234767
rect 40682 228304 40738 228313
rect 40682 228239 40738 228248
rect 36542 228168 36598 228177
rect 36542 228103 36598 228112
rect 36556 59362 36584 228103
rect 36544 59356 36596 59362
rect 36544 59298 36596 59304
rect 35808 57112 35860 57118
rect 35808 57054 35860 57060
rect 34428 56500 34480 56506
rect 34428 56442 34480 56448
rect 33784 20664 33836 20670
rect 33784 20606 33836 20612
rect 34440 3466 34468 56442
rect 35820 3466 35848 57054
rect 39948 57044 40000 57050
rect 39948 56986 40000 56992
rect 37188 54528 37240 54534
rect 37188 54470 37240 54476
rect 35992 4004 36044 4010
rect 35992 3946 36044 3952
rect 32404 3460 32456 3466
rect 32404 3402 32456 3408
rect 33048 3460 33100 3466
rect 33048 3402 33100 3408
rect 33600 3460 33652 3466
rect 33600 3402 33652 3408
rect 34428 3460 34480 3466
rect 34428 3402 34480 3408
rect 34796 3460 34848 3466
rect 34796 3402 34848 3408
rect 35808 3460 35860 3466
rect 35808 3402 35860 3408
rect 32416 480 32444 3402
rect 33612 480 33640 3402
rect 34808 480 34836 3402
rect 36004 480 36032 3946
rect 37200 480 37228 54470
rect 39960 6914 39988 56986
rect 40696 45558 40724 228239
rect 50632 183326 50660 503882
rect 50712 429208 50764 429214
rect 50712 429150 50764 429156
rect 50620 183320 50672 183326
rect 50620 183262 50672 183268
rect 50724 59362 50752 429150
rect 50816 107642 50844 504018
rect 50894 503840 50950 503849
rect 50894 503775 50950 503784
rect 50804 107636 50856 107642
rect 50804 107578 50856 107584
rect 50908 85542 50936 503775
rect 50896 85536 50948 85542
rect 50896 85478 50948 85484
rect 51000 80034 51028 504047
rect 52184 504008 52236 504014
rect 52184 503950 52236 503956
rect 52092 399696 52144 399702
rect 52092 399638 52144 399644
rect 52000 399492 52052 399498
rect 52000 399434 52052 399440
rect 51908 395480 51960 395486
rect 51908 395422 51960 395428
rect 51816 249076 51868 249082
rect 51816 249018 51868 249024
rect 51724 247920 51776 247926
rect 51724 247862 51776 247868
rect 51632 245268 51684 245274
rect 51632 245210 51684 245216
rect 51644 180810 51672 245210
rect 51632 180804 51684 180810
rect 51632 180746 51684 180752
rect 51736 169726 51764 247862
rect 51724 169720 51776 169726
rect 51724 169662 51776 169668
rect 51828 144226 51856 249018
rect 51816 144220 51868 144226
rect 51816 144162 51868 144168
rect 51920 115598 51948 395422
rect 51908 115592 51960 115598
rect 51908 115534 51960 115540
rect 52012 102134 52040 399434
rect 52000 102128 52052 102134
rect 52000 102070 52052 102076
rect 52104 88330 52132 399638
rect 52196 118658 52224 503950
rect 52184 118652 52236 118658
rect 52184 118594 52236 118600
rect 52092 88324 52144 88330
rect 52092 88266 52144 88272
rect 50988 80028 51040 80034
rect 50988 79970 51040 79976
rect 52288 75886 52316 504154
rect 52276 75880 52328 75886
rect 52276 75822 52328 75828
rect 52380 70378 52408 504183
rect 53196 503872 53248 503878
rect 53196 503814 53248 503820
rect 53104 240848 53156 240854
rect 53104 240790 53156 240796
rect 53116 104854 53144 240790
rect 53208 184890 53236 503814
rect 53196 184884 53248 184890
rect 53196 184826 53248 184832
rect 53300 167006 53328 504902
rect 55036 504756 55088 504762
rect 55036 504698 55088 504704
rect 53746 503976 53802 503985
rect 53746 503911 53802 503920
rect 53380 503736 53432 503742
rect 53380 503678 53432 503684
rect 53288 167000 53340 167006
rect 53288 166942 53340 166948
rect 53392 163538 53420 503678
rect 53472 503668 53524 503674
rect 53472 503610 53524 503616
rect 53380 163532 53432 163538
rect 53380 163474 53432 163480
rect 53484 153202 53512 503610
rect 53656 503600 53708 503606
rect 53656 503542 53708 503548
rect 53564 503464 53616 503470
rect 53564 503406 53616 503412
rect 53472 153196 53524 153202
rect 53472 153138 53524 153144
rect 53576 133890 53604 503406
rect 53564 133884 53616 133890
rect 53564 133826 53616 133832
rect 53668 110430 53696 503542
rect 53656 110424 53708 110430
rect 53656 110366 53708 110372
rect 53104 104848 53156 104854
rect 53104 104790 53156 104796
rect 53760 91050 53788 503911
rect 54852 395548 54904 395554
rect 54852 395490 54904 395496
rect 54760 358080 54812 358086
rect 54760 358022 54812 358028
rect 54208 248396 54260 248402
rect 54208 248338 54260 248344
rect 54220 161430 54248 248338
rect 54576 247852 54628 247858
rect 54576 247794 54628 247800
rect 54484 246832 54536 246838
rect 54484 246774 54536 246780
rect 54300 246764 54352 246770
rect 54300 246706 54352 246712
rect 54208 161424 54260 161430
rect 54208 161366 54260 161372
rect 54312 158710 54340 246706
rect 54392 244044 54444 244050
rect 54392 243986 54444 243992
rect 54300 158704 54352 158710
rect 54300 158646 54352 158652
rect 54404 150414 54432 243986
rect 54392 150408 54444 150414
rect 54392 150350 54444 150356
rect 54496 136610 54524 246774
rect 54484 136604 54536 136610
rect 54484 136546 54536 136552
rect 54588 132462 54616 247794
rect 54668 240916 54720 240922
rect 54668 240858 54720 240864
rect 54576 132456 54628 132462
rect 54576 132398 54628 132404
rect 53748 91044 53800 91050
rect 53748 90986 53800 90992
rect 54680 78674 54708 240858
rect 54772 190466 54800 358022
rect 54760 190460 54812 190466
rect 54760 190402 54812 190408
rect 54864 172514 54892 395490
rect 54944 395412 54996 395418
rect 54944 395354 54996 395360
rect 54852 172508 54904 172514
rect 54852 172450 54904 172456
rect 54956 142118 54984 395354
rect 55048 198694 55076 504698
rect 56416 504484 56468 504490
rect 56416 504426 56468 504432
rect 55128 503804 55180 503810
rect 55128 503746 55180 503752
rect 55036 198688 55088 198694
rect 55036 198630 55088 198636
rect 55140 195974 55168 503746
rect 55864 247784 55916 247790
rect 55864 247726 55916 247732
rect 55678 226400 55734 226409
rect 55678 226335 55734 226344
rect 55128 195968 55180 195974
rect 55128 195910 55180 195916
rect 54944 142112 54996 142118
rect 54944 142054 54996 142060
rect 54668 78668 54720 78674
rect 54668 78610 54720 78616
rect 52368 70372 52420 70378
rect 52368 70314 52420 70320
rect 50712 59356 50764 59362
rect 50712 59298 50764 59304
rect 43444 56976 43496 56982
rect 43444 56918 43496 56924
rect 41328 55820 41380 55826
rect 41328 55762 41380 55768
rect 40684 45552 40736 45558
rect 40684 45494 40736 45500
rect 39592 6886 39988 6914
rect 38384 4072 38436 4078
rect 38384 4014 38436 4020
rect 38396 480 38424 4014
rect 39592 480 39620 6886
rect 41340 3466 41368 55762
rect 43076 4140 43128 4146
rect 43076 4082 43128 4088
rect 40684 3460 40736 3466
rect 40684 3402 40736 3408
rect 41328 3460 41380 3466
rect 41328 3402 41380 3408
rect 41880 3460 41932 3466
rect 41880 3402 41932 3408
rect 40696 480 40724 3402
rect 41892 480 41920 3402
rect 43088 480 43116 4082
rect 43456 3466 43484 56918
rect 53748 56908 53800 56914
rect 53748 56850 53800 56856
rect 50344 56840 50396 56846
rect 50344 56782 50396 56788
rect 48228 55752 48280 55758
rect 48228 55694 48280 55700
rect 48240 6914 48268 55694
rect 47872 6886 48268 6914
rect 43444 3460 43496 3466
rect 43444 3402 43496 3408
rect 46664 3460 46716 3466
rect 46664 3402 46716 3408
rect 45468 3392 45520 3398
rect 45468 3334 45520 3340
rect 44272 3324 44324 3330
rect 44272 3266 44324 3272
rect 44284 480 44312 3266
rect 45480 480 45508 3334
rect 46676 480 46704 3402
rect 47872 480 47900 6886
rect 50356 3466 50384 56782
rect 52368 55684 52420 55690
rect 52368 55626 52420 55632
rect 52380 3466 52408 55626
rect 50344 3460 50396 3466
rect 50344 3402 50396 3408
rect 51356 3460 51408 3466
rect 51356 3402 51408 3408
rect 52368 3460 52420 3466
rect 52368 3402 52420 3408
rect 50160 3256 50212 3262
rect 50160 3198 50212 3204
rect 48964 3052 49016 3058
rect 48964 2994 49016 3000
rect 48976 480 49004 2994
rect 50172 480 50200 3198
rect 51368 480 51396 3402
rect 52552 3120 52604 3126
rect 52552 3062 52604 3068
rect 52564 480 52592 3062
rect 53760 480 53788 56850
rect 55128 55616 55180 55622
rect 55128 55558 55180 55564
rect 55140 6914 55168 55558
rect 55692 20670 55720 226335
rect 55770 226128 55826 226137
rect 55770 226063 55826 226072
rect 55784 33114 55812 226063
rect 55876 192953 55904 247726
rect 55956 246084 56008 246090
rect 55956 246026 56008 246032
rect 55862 192944 55918 192953
rect 55862 192879 55918 192888
rect 55968 176905 55996 246026
rect 56048 246016 56100 246022
rect 56048 245958 56100 245964
rect 55954 176896 56010 176905
rect 55954 176831 56010 176840
rect 56060 139233 56088 245958
rect 56324 243296 56376 243302
rect 56324 243238 56376 243244
rect 56232 242208 56284 242214
rect 56232 242150 56284 242156
rect 56140 227792 56192 227798
rect 56140 227734 56192 227740
rect 56046 139224 56102 139233
rect 56046 139159 56102 139168
rect 56152 55962 56180 227734
rect 56244 66609 56272 242150
rect 56336 222601 56364 243238
rect 56428 225321 56456 504426
rect 56414 225312 56470 225321
rect 56414 225247 56470 225256
rect 56322 222592 56378 222601
rect 56322 222527 56378 222536
rect 56520 203833 56548 505038
rect 57612 505028 57664 505034
rect 57612 504970 57664 504976
rect 57520 504620 57572 504626
rect 57520 504562 57572 504568
rect 57242 435976 57298 435985
rect 57242 435911 57298 435920
rect 57150 432848 57206 432857
rect 57150 432783 57206 432792
rect 57058 410000 57114 410009
rect 57058 409935 57114 409944
rect 56966 407552 57022 407561
rect 56966 407487 57022 407496
rect 56980 399634 57008 407487
rect 56968 399628 57020 399634
rect 56968 399570 57020 399576
rect 57072 242690 57100 409935
rect 57060 242684 57112 242690
rect 57060 242626 57112 242632
rect 57164 242486 57192 432783
rect 57152 242480 57204 242486
rect 57152 242422 57204 242428
rect 57256 242185 57284 435911
rect 57426 433800 57482 433809
rect 57426 433735 57482 433744
rect 57334 429992 57390 430001
rect 57334 429927 57390 429936
rect 57348 429214 57376 429927
rect 57336 429208 57388 429214
rect 57336 429150 57388 429156
rect 57336 426692 57388 426698
rect 57336 426634 57388 426640
rect 57242 242176 57298 242185
rect 57242 242111 57298 242120
rect 57152 240984 57204 240990
rect 57152 240926 57204 240932
rect 56506 203824 56562 203833
rect 56506 203759 56562 203768
rect 56876 180804 56928 180810
rect 56876 180746 56928 180752
rect 56888 179625 56916 180746
rect 56874 179616 56930 179625
rect 56874 179551 56930 179560
rect 57164 96257 57192 240926
rect 57348 201482 57376 426634
rect 57336 201476 57388 201482
rect 57336 201418 57388 201424
rect 57244 161424 57296 161430
rect 57244 161366 57296 161372
rect 57256 160721 57284 161366
rect 57242 160712 57298 160721
rect 57242 160647 57298 160656
rect 57440 155922 57468 433735
rect 57532 217161 57560 504562
rect 57518 217152 57574 217161
rect 57518 217087 57574 217096
rect 57624 211857 57652 504970
rect 58348 504892 58400 504898
rect 58348 504834 58400 504840
rect 57796 504144 57848 504150
rect 57796 504086 57848 504092
rect 57702 436928 57758 436937
rect 57702 436863 57758 436872
rect 57610 211848 57666 211857
rect 57610 211783 57666 211792
rect 57612 198688 57664 198694
rect 57612 198630 57664 198636
rect 57624 198393 57652 198630
rect 57610 198384 57666 198393
rect 57610 198319 57666 198328
rect 57612 195968 57664 195974
rect 57612 195910 57664 195916
rect 57624 195673 57652 195910
rect 57610 195664 57666 195673
rect 57610 195599 57666 195608
rect 57612 190460 57664 190466
rect 57612 190402 57664 190408
rect 57624 190369 57652 190402
rect 57610 190360 57666 190369
rect 57610 190295 57666 190304
rect 57610 184920 57666 184929
rect 57610 184855 57612 184864
rect 57664 184855 57666 184864
rect 57612 184826 57664 184832
rect 57612 183320 57664 183326
rect 57612 183262 57664 183268
rect 57624 182209 57652 183262
rect 57610 182200 57666 182209
rect 57610 182135 57666 182144
rect 57612 172508 57664 172514
rect 57612 172450 57664 172456
rect 57624 171465 57652 172450
rect 57610 171456 57666 171465
rect 57610 171391 57666 171400
rect 57612 169720 57664 169726
rect 57612 169662 57664 169668
rect 57624 168745 57652 169662
rect 57610 168736 57666 168745
rect 57610 168671 57666 168680
rect 57612 167000 57664 167006
rect 57612 166942 57664 166948
rect 57624 166161 57652 166942
rect 57610 166152 57666 166161
rect 57610 166087 57666 166096
rect 57612 163532 57664 163538
rect 57612 163474 57664 163480
rect 57624 163441 57652 163474
rect 57610 163432 57666 163441
rect 57610 163367 57666 163376
rect 57612 158704 57664 158710
rect 57612 158646 57664 158652
rect 57624 158001 57652 158646
rect 57610 157992 57666 158001
rect 57610 157927 57666 157936
rect 57428 155916 57480 155922
rect 57428 155858 57480 155864
rect 57612 153196 57664 153202
rect 57612 153138 57664 153144
rect 57624 152697 57652 153138
rect 57610 152688 57666 152697
rect 57610 152623 57666 152632
rect 57612 150408 57664 150414
rect 57612 150350 57664 150356
rect 57624 149977 57652 150350
rect 57610 149968 57666 149977
rect 57610 149903 57666 149912
rect 57610 144664 57666 144673
rect 57610 144599 57666 144608
rect 57624 144226 57652 144599
rect 57612 144220 57664 144226
rect 57612 144162 57664 144168
rect 57612 142112 57664 142118
rect 57612 142054 57664 142060
rect 57624 141953 57652 142054
rect 57610 141944 57666 141953
rect 57610 141879 57666 141888
rect 57612 136604 57664 136610
rect 57612 136546 57664 136552
rect 57624 136513 57652 136546
rect 57610 136504 57666 136513
rect 57610 136439 57666 136448
rect 57612 133884 57664 133890
rect 57612 133826 57664 133832
rect 57624 133793 57652 133826
rect 57610 133784 57666 133793
rect 57610 133719 57666 133728
rect 57612 132456 57664 132462
rect 57612 132398 57664 132404
rect 57624 131209 57652 132398
rect 57610 131200 57666 131209
rect 57610 131135 57666 131144
rect 57716 120465 57744 436863
rect 57808 123049 57836 504086
rect 57886 431080 57942 431089
rect 57886 431015 57942 431024
rect 57900 426698 57928 431015
rect 57888 426692 57940 426698
rect 57888 426634 57940 426640
rect 57886 408232 57942 408241
rect 57886 408167 57942 408176
rect 57900 398818 57928 408167
rect 57888 398812 57940 398818
rect 57888 398754 57940 398760
rect 57900 241466 57928 398754
rect 58164 242344 58216 242350
rect 58164 242286 58216 242292
rect 57888 241460 57940 241466
rect 57888 241402 57940 241408
rect 57886 225992 57942 226001
rect 57886 225927 57942 225936
rect 57900 219881 57928 225927
rect 57886 219872 57942 219881
rect 57886 219807 57942 219816
rect 58176 174185 58204 242286
rect 58256 241392 58308 241398
rect 58256 241334 58308 241340
rect 58162 174176 58218 174185
rect 58162 174111 58218 174120
rect 57794 123040 57850 123049
rect 57794 122975 57850 122984
rect 57702 120456 57758 120465
rect 57702 120391 57758 120400
rect 57612 118652 57664 118658
rect 57612 118594 57664 118600
rect 57624 117745 57652 118594
rect 57610 117736 57666 117745
rect 57610 117671 57666 117680
rect 57612 115592 57664 115598
rect 57612 115534 57664 115540
rect 57624 115025 57652 115534
rect 57610 115016 57666 115025
rect 57610 114951 57666 114960
rect 58268 112305 58296 241334
rect 58360 228449 58388 504834
rect 59082 428224 59138 428233
rect 59082 428159 59138 428168
rect 59096 398041 59124 428159
rect 59280 399566 59308 700266
rect 89180 699718 89208 703520
rect 105464 699718 105492 703520
rect 88340 699712 88392 699718
rect 88340 699654 88392 699660
rect 89168 699712 89220 699718
rect 89168 699654 89220 699660
rect 104900 699712 104952 699718
rect 104900 699654 104952 699660
rect 105452 699712 105504 699718
rect 105452 699654 105504 699660
rect 88352 504422 88380 699654
rect 89628 505776 89680 505782
rect 89628 505718 89680 505724
rect 60004 504416 60056 504422
rect 60004 504358 60056 504364
rect 88340 504416 88392 504422
rect 88340 504358 88392 504364
rect 59268 399560 59320 399566
rect 59268 399502 59320 399508
rect 59082 398032 59138 398041
rect 59082 397967 59138 397976
rect 58808 397248 58860 397254
rect 58808 397190 58860 397196
rect 58716 396908 58768 396914
rect 58716 396850 58768 396856
rect 58532 396840 58584 396846
rect 58532 396782 58584 396788
rect 58440 396772 58492 396778
rect 58440 396714 58492 396720
rect 58346 228440 58402 228449
rect 58346 228375 58402 228384
rect 58346 225584 58402 225593
rect 58346 225519 58402 225528
rect 58254 112296 58310 112305
rect 58254 112231 58310 112240
rect 57612 110424 57664 110430
rect 57612 110366 57664 110372
rect 57624 109585 57652 110366
rect 57610 109576 57666 109585
rect 57610 109511 57666 109520
rect 57612 107636 57664 107642
rect 57612 107578 57664 107584
rect 57624 107001 57652 107578
rect 57610 106992 57666 107001
rect 57610 106927 57666 106936
rect 57612 104848 57664 104854
rect 57612 104790 57664 104796
rect 57624 104281 57652 104790
rect 57610 104272 57666 104281
rect 57610 104207 57666 104216
rect 57612 102128 57664 102134
rect 57612 102070 57664 102076
rect 57624 101561 57652 102070
rect 57610 101552 57666 101561
rect 57610 101487 57666 101496
rect 57150 96248 57206 96257
rect 57150 96183 57206 96192
rect 57612 91044 57664 91050
rect 57612 90986 57664 90992
rect 57624 90817 57652 90986
rect 57610 90808 57666 90817
rect 57610 90743 57666 90752
rect 57612 88324 57664 88330
rect 57612 88266 57664 88272
rect 57624 88097 57652 88266
rect 57610 88088 57666 88097
rect 57610 88023 57666 88032
rect 57612 85536 57664 85542
rect 57612 85478 57664 85484
rect 57624 85377 57652 85478
rect 57610 85368 57666 85377
rect 57610 85303 57666 85312
rect 57610 80064 57666 80073
rect 57610 79999 57612 80008
rect 57664 79999 57666 80008
rect 57612 79970 57664 79976
rect 57612 78668 57664 78674
rect 57612 78610 57664 78616
rect 57624 77353 57652 78610
rect 57610 77344 57666 77353
rect 57610 77279 57666 77288
rect 57612 75880 57664 75886
rect 57612 75822 57664 75828
rect 57624 74633 57652 75822
rect 57610 74624 57666 74633
rect 57610 74559 57666 74568
rect 57612 70372 57664 70378
rect 57612 70314 57664 70320
rect 57624 69329 57652 70314
rect 57610 69320 57666 69329
rect 57610 69255 57666 69264
rect 56230 66600 56286 66609
rect 56230 66535 56286 66544
rect 58360 57866 58388 225519
rect 58452 209137 58480 396714
rect 58438 209128 58494 209137
rect 58438 209063 58494 209072
rect 58544 206417 58572 396782
rect 58624 241460 58676 241466
rect 58624 241402 58676 241408
rect 58530 206408 58586 206417
rect 58530 206343 58586 206352
rect 58532 201476 58584 201482
rect 58532 201418 58584 201424
rect 58544 98841 58572 201418
rect 58530 98832 58586 98841
rect 58530 98767 58586 98776
rect 58636 60314 58664 241402
rect 58728 201113 58756 396850
rect 58714 201104 58770 201113
rect 58714 201039 58770 201048
rect 58820 187649 58848 397190
rect 58992 397112 59044 397118
rect 58992 397054 59044 397060
rect 58900 396636 58952 396642
rect 58900 396578 58952 396584
rect 58806 187640 58862 187649
rect 58806 187575 58862 187584
rect 58716 155916 58768 155922
rect 58716 155858 58768 155864
rect 58624 60308 58676 60314
rect 58624 60250 58676 60256
rect 58728 57905 58756 155858
rect 58912 155417 58940 396578
rect 58898 155408 58954 155417
rect 58898 155343 58954 155352
rect 59004 147257 59032 397054
rect 59268 396500 59320 396506
rect 59268 396442 59320 396448
rect 59084 396432 59136 396438
rect 59084 396374 59136 396380
rect 58990 147248 59046 147257
rect 58990 147183 59046 147192
rect 59096 128489 59124 396374
rect 59176 241188 59228 241194
rect 59176 241130 59228 241136
rect 59082 128480 59138 128489
rect 59082 128415 59138 128424
rect 59188 61305 59216 241130
rect 59280 93537 59308 396442
rect 59728 396296 59780 396302
rect 59728 396238 59780 396244
rect 59452 396228 59504 396234
rect 59452 396170 59504 396176
rect 59266 93528 59322 93537
rect 59266 93463 59322 93472
rect 59464 82793 59492 396170
rect 59544 396160 59596 396166
rect 59544 396102 59596 396108
rect 59556 125769 59584 396102
rect 59636 240780 59688 240786
rect 59636 240722 59688 240728
rect 59648 214577 59676 240722
rect 59634 214568 59690 214577
rect 59634 214503 59690 214512
rect 59542 125760 59598 125769
rect 59542 125695 59598 125704
rect 59450 82784 59506 82793
rect 59450 82719 59506 82728
rect 59740 72049 59768 396238
rect 60016 232529 60044 504358
rect 89640 503577 89668 505718
rect 91006 505200 91062 505209
rect 91006 505135 91062 505144
rect 89626 503568 89682 503577
rect 89626 503503 89682 503512
rect 91020 495434 91048 505135
rect 104912 504898 104940 699654
rect 137848 698306 137876 703520
rect 154132 700330 154160 703520
rect 170324 700398 170352 703520
rect 202800 703050 202828 703520
rect 201500 703044 201552 703050
rect 201500 702986 201552 702992
rect 202788 703044 202840 703050
rect 202788 702986 202840 702992
rect 198004 700528 198056 700534
rect 198004 700470 198056 700476
rect 170312 700392 170364 700398
rect 170312 700334 170364 700340
rect 196532 700392 196584 700398
rect 196532 700334 196584 700340
rect 154120 700324 154172 700330
rect 154120 700266 154172 700272
rect 137848 698278 138060 698306
rect 138032 696930 138060 698278
rect 138020 696924 138072 696930
rect 138020 696866 138072 696872
rect 140044 696924 140096 696930
rect 140044 696866 140096 696872
rect 140056 689654 140084 696866
rect 140044 689648 140096 689654
rect 140044 689590 140096 689596
rect 141148 689648 141200 689654
rect 141148 689590 141200 689596
rect 141160 683670 141188 689590
rect 141148 683664 141200 683670
rect 141148 683606 141200 683612
rect 143540 683664 143592 683670
rect 143540 683606 143592 683612
rect 143552 680542 143580 683606
rect 143540 680536 143592 680542
rect 143540 680478 143592 680484
rect 145564 680536 145616 680542
rect 145564 680478 145616 680484
rect 145576 663270 145604 680478
rect 145564 663264 145616 663270
rect 145564 663206 145616 663212
rect 149704 663264 149756 663270
rect 149704 663206 149756 663212
rect 149716 645930 149744 663206
rect 149704 645924 149756 645930
rect 149704 645866 149756 645872
rect 153200 645856 153252 645862
rect 153200 645798 153252 645804
rect 153212 638926 153240 645798
rect 153200 638920 153252 638926
rect 153200 638862 153252 638868
rect 155224 638920 155276 638926
rect 155224 638862 155276 638868
rect 155236 627978 155264 638862
rect 155224 627972 155276 627978
rect 155224 627914 155276 627920
rect 160468 627904 160520 627910
rect 160468 627846 160520 627852
rect 160480 619682 160508 627846
rect 160468 619676 160520 619682
rect 160468 619618 160520 619624
rect 163504 619608 163556 619614
rect 163504 619550 163556 619556
rect 163516 611998 163544 619550
rect 163504 611992 163556 611998
rect 163504 611934 163556 611940
rect 164884 611992 164936 611998
rect 164884 611934 164936 611940
rect 164896 585750 164924 611934
rect 164884 585744 164936 585750
rect 164884 585686 164936 585692
rect 167552 585744 167604 585750
rect 167552 585686 167604 585692
rect 167564 579630 167592 585686
rect 167552 579624 167604 579630
rect 167552 579566 167604 579572
rect 170404 579624 170456 579630
rect 170404 579566 170456 579572
rect 170416 569158 170444 579566
rect 170404 569152 170456 569158
rect 170404 569094 170456 569100
rect 172428 569152 172480 569158
rect 172428 569094 172480 569100
rect 172440 563106 172468 569094
rect 172428 563100 172480 563106
rect 172428 563042 172480 563048
rect 178040 563032 178092 563038
rect 178040 562974 178092 562980
rect 178052 560250 178080 562974
rect 178040 560244 178092 560250
rect 178040 560186 178092 560192
rect 180708 560244 180760 560250
rect 180708 560186 180760 560192
rect 180720 552090 180748 560186
rect 180708 552084 180760 552090
rect 180708 552026 180760 552032
rect 182824 552016 182876 552022
rect 182824 551958 182876 551964
rect 182836 542366 182864 551958
rect 182824 542360 182876 542366
rect 182824 542302 182876 542308
rect 184204 542360 184256 542366
rect 184204 542302 184256 542308
rect 184216 534138 184244 542302
rect 184204 534132 184256 534138
rect 184204 534074 184256 534080
rect 186136 534132 186188 534138
rect 186136 534074 186188 534080
rect 186148 531350 186176 534074
rect 186136 531344 186188 531350
rect 186136 531286 186188 531292
rect 187700 531276 187752 531282
rect 187700 531218 187752 531224
rect 187712 529242 187740 531218
rect 187700 529236 187752 529242
rect 187700 529178 187752 529184
rect 114468 505708 114520 505714
rect 114468 505650 114520 505656
rect 104900 504892 104952 504898
rect 104900 504834 104952 504840
rect 108948 504892 109000 504898
rect 108948 504834 109000 504840
rect 98552 504688 98604 504694
rect 98552 504630 98604 504636
rect 96528 504280 96580 504286
rect 96528 504222 96580 504228
rect 96540 503577 96568 504222
rect 98564 503577 98592 504630
rect 103888 504416 103940 504422
rect 103888 504358 103940 504364
rect 101312 504348 101364 504354
rect 101312 504290 101364 504296
rect 101324 503577 101352 504290
rect 103900 503577 103928 504358
rect 104072 503600 104124 503606
rect 96526 503568 96582 503577
rect 93768 503532 93820 503538
rect 96526 503503 96582 503512
rect 98550 503568 98606 503577
rect 98550 503503 98606 503512
rect 101310 503568 101366 503577
rect 101310 503503 101366 503512
rect 103886 503568 103942 503577
rect 103886 503503 103942 503512
rect 104070 503568 104072 503577
rect 104124 503568 104126 503577
rect 104070 503503 104126 503512
rect 93768 503474 93820 503480
rect 93780 500954 93808 503474
rect 108960 502334 108988 504834
rect 111708 504552 111760 504558
rect 111708 504494 111760 504500
rect 111720 502334 111748 504494
rect 113546 503568 113602 503577
rect 113546 503503 113602 503512
rect 113560 503470 113588 503503
rect 113548 503464 113600 503470
rect 113548 503406 113600 503412
rect 114480 502334 114508 505650
rect 144828 505640 144880 505646
rect 144828 505582 144880 505588
rect 142068 505572 142120 505578
rect 142068 505514 142120 505520
rect 133788 505436 133840 505442
rect 133788 505378 133840 505384
rect 129648 505368 129700 505374
rect 129648 505310 129700 505316
rect 117228 505300 117280 505306
rect 117228 505242 117280 505248
rect 117240 503713 117268 505242
rect 128636 504960 128688 504966
rect 128636 504902 128688 504908
rect 128648 503713 128676 504902
rect 129660 504393 129688 505310
rect 129646 504384 129702 504393
rect 129646 504319 129702 504328
rect 129740 503736 129792 503742
rect 117226 503704 117282 503713
rect 128634 503704 128690 503713
rect 117226 503639 117282 503648
rect 123760 503668 123812 503674
rect 129740 503678 129792 503684
rect 128634 503639 128690 503648
rect 123760 503610 123812 503616
rect 123772 503577 123800 503610
rect 129752 503577 129780 503678
rect 123574 503568 123630 503577
rect 123574 503503 123576 503512
rect 123628 503503 123630 503512
rect 123758 503568 123814 503577
rect 123758 503503 123814 503512
rect 129738 503568 129794 503577
rect 129738 503503 129794 503512
rect 123576 503474 123628 503480
rect 121368 503464 121420 503470
rect 121368 503406 121420 503412
rect 108684 502306 108988 502334
rect 111260 502306 111748 502334
rect 111996 502306 114508 502334
rect 108684 500954 108712 502306
rect 89824 495406 91048 495434
rect 91572 500926 93808 500954
rect 108500 500926 108712 500954
rect 89824 494054 89852 495406
rect 89548 494026 89852 494054
rect 89548 490385 89576 494026
rect 91572 490385 91600 500926
rect 108500 495434 108528 500926
rect 108408 495406 108528 495434
rect 108408 494054 108436 495406
rect 108316 494026 108436 494054
rect 108316 491065 108344 494026
rect 111260 493354 111288 502306
rect 110984 493326 111288 493354
rect 110984 492674 111012 493326
rect 110892 492646 111012 492674
rect 108302 491056 108358 491065
rect 108302 490991 108358 491000
rect 89534 490376 89590 490385
rect 89534 490311 89590 490320
rect 91558 490376 91614 490385
rect 91558 490311 91614 490320
rect 110892 489914 110920 492646
rect 110800 489886 110920 489914
rect 110800 488534 110828 489886
rect 110800 488506 110920 488534
rect 110892 487154 110920 488506
rect 111996 488345 112024 502306
rect 121380 499574 121408 503406
rect 133800 502334 133828 505378
rect 133708 502306 133828 502334
rect 142080 502334 142108 505514
rect 143356 505504 143408 505510
rect 143356 505446 143408 505452
rect 143368 503577 143396 505446
rect 143354 503568 143410 503577
rect 143354 503503 143410 503512
rect 144458 503568 144514 503577
rect 144458 503503 144514 503512
rect 144472 502334 144500 503503
rect 144840 502334 144868 505582
rect 153200 505096 153252 505102
rect 153200 505038 153252 505044
rect 158628 505096 158680 505102
rect 158628 505038 158680 505044
rect 148508 504960 148560 504966
rect 148508 504902 148560 504908
rect 146576 504824 146628 504830
rect 146576 504766 146628 504772
rect 146588 503577 146616 504766
rect 148520 503713 148548 504902
rect 149520 504756 149572 504762
rect 149520 504698 149572 504704
rect 148506 503704 148562 503713
rect 148506 503639 148562 503648
rect 149532 503577 149560 504698
rect 146574 503568 146630 503577
rect 146574 503503 146630 503512
rect 149518 503568 149574 503577
rect 149518 503503 149574 503512
rect 142080 502306 144500 502334
rect 144564 502306 144868 502334
rect 133708 500954 133736 502306
rect 120828 499546 121408 499574
rect 133616 500926 133736 500954
rect 144564 500954 144592 502306
rect 144564 500926 145052 500954
rect 120828 498194 120856 499546
rect 118528 498166 120856 498194
rect 111982 488336 112038 488345
rect 111982 488271 112038 488280
rect 110800 487126 110920 487154
rect 110800 485774 110828 487126
rect 110616 485746 110828 485774
rect 110616 484394 110644 485746
rect 118528 485217 118556 498166
rect 133616 491881 133644 500926
rect 145024 499574 145052 500926
rect 153212 499574 153240 505038
rect 156052 504620 156104 504626
rect 156052 504562 156104 504568
rect 156064 503577 156092 504562
rect 158640 503577 158668 505038
rect 164056 504960 164108 504966
rect 164056 504902 164108 504908
rect 160100 503736 160152 503742
rect 160100 503678 160152 503684
rect 160112 503577 160140 503678
rect 164068 503577 164096 504902
rect 165620 504484 165672 504490
rect 165620 504426 165672 504432
rect 165632 503577 165660 504426
rect 176844 504212 176896 504218
rect 176844 504154 176896 504160
rect 176856 503713 176884 504154
rect 180708 503736 180760 503742
rect 176842 503704 176898 503713
rect 180708 503678 180760 503684
rect 176842 503639 176898 503648
rect 156050 503568 156106 503577
rect 156050 503503 156106 503512
rect 158626 503568 158682 503577
rect 158626 503503 158682 503512
rect 160098 503568 160154 503577
rect 160098 503503 160154 503512
rect 164054 503568 164110 503577
rect 164054 503503 164110 503512
rect 165618 503568 165674 503577
rect 165618 503503 165674 503512
rect 144748 499546 145052 499574
rect 153028 499546 153240 499574
rect 144748 496814 144776 499546
rect 144748 496786 144960 496814
rect 144932 492674 144960 496786
rect 144932 492646 145236 492674
rect 133602 491872 133658 491881
rect 133602 491807 133658 491816
rect 145208 491294 145236 492646
rect 153028 491745 153056 499546
rect 180720 495434 180748 503678
rect 191748 503464 191800 503470
rect 191748 503406 191800 503412
rect 180628 495406 180748 495434
rect 180628 494054 180656 495406
rect 179616 494026 180656 494054
rect 153014 491736 153070 491745
rect 153014 491671 153070 491680
rect 143552 491266 145236 491294
rect 179616 491294 179644 494026
rect 179616 491266 179736 491294
rect 143552 489914 143580 491266
rect 179708 489914 179736 491266
rect 191760 490906 191788 503406
rect 196544 495434 196572 700334
rect 196624 700324 196676 700330
rect 196624 700266 196676 700272
rect 196360 495406 196572 495434
rect 196360 494054 196388 495406
rect 195900 494026 196388 494054
rect 191760 490878 194732 490906
rect 143460 489886 143580 489914
rect 179616 489886 179736 489914
rect 143460 488534 143488 489886
rect 143368 488506 143488 488534
rect 179616 488534 179644 489886
rect 194704 488534 194732 490878
rect 179616 488506 179736 488534
rect 194704 488506 195836 488534
rect 143368 487154 143396 488506
rect 179708 487154 179736 488506
rect 143368 487126 143488 487154
rect 143460 485774 143488 487126
rect 179524 487126 179736 487154
rect 179524 485774 179552 487126
rect 195808 486282 195836 488506
rect 195900 487234 195928 494026
rect 196636 487370 196664 700266
rect 196808 529236 196860 529242
rect 196808 529178 196860 529184
rect 196716 503328 196768 503334
rect 196716 503270 196768 503276
rect 196728 488534 196756 503270
rect 196820 489914 196848 529178
rect 197452 504892 197504 504898
rect 197452 504834 197504 504840
rect 197360 504688 197412 504694
rect 197360 504630 197412 504636
rect 196820 489886 197032 489914
rect 196728 488506 196848 488534
rect 196636 487354 196756 487370
rect 196636 487348 196768 487354
rect 196636 487342 196716 487348
rect 196716 487290 196768 487296
rect 195900 487206 196756 487234
rect 196728 486402 196756 487206
rect 196716 486396 196768 486402
rect 196716 486338 196768 486344
rect 196714 486296 196770 486305
rect 195808 486254 196714 486282
rect 196714 486231 196770 486240
rect 196716 486192 196768 486198
rect 143460 485746 143764 485774
rect 118514 485208 118570 485217
rect 118514 485143 118570 485152
rect 143736 484394 143764 485746
rect 110616 484366 111472 484394
rect 111444 483721 111472 484366
rect 143092 484366 143764 484394
rect 179340 485746 179552 485774
rect 196544 486140 196716 486146
rect 196544 486134 196768 486140
rect 196544 486118 196756 486134
rect 179340 484394 179368 485746
rect 179340 484366 180288 484394
rect 143092 484129 143120 484366
rect 180260 484129 180288 484366
rect 143078 484120 143134 484129
rect 143078 484055 143134 484064
rect 180246 484120 180302 484129
rect 180246 484055 180302 484064
rect 111430 483712 111486 483721
rect 111430 483647 111486 483656
rect 176568 400036 176620 400042
rect 176568 399978 176620 399984
rect 187608 400036 187660 400042
rect 187608 399978 187660 399984
rect 115756 399900 115808 399906
rect 115756 399842 115808 399848
rect 113088 399764 113140 399770
rect 113088 399706 113140 399712
rect 85486 398168 85542 398177
rect 85486 398103 85542 398112
rect 92386 398168 92442 398177
rect 92386 398103 92442 398112
rect 95974 398168 96030 398177
rect 95974 398103 96030 398112
rect 99378 398168 99434 398177
rect 99378 398103 99434 398112
rect 81992 397452 82044 397458
rect 81992 397394 82044 397400
rect 82004 397361 82032 397394
rect 85500 397390 85528 398103
rect 85488 397384 85540 397390
rect 78310 397352 78366 397361
rect 61476 397316 61528 397322
rect 78310 397287 78366 397296
rect 80978 397352 81034 397361
rect 80978 397287 81034 397296
rect 81990 397352 82046 397361
rect 81990 397287 82046 397296
rect 83370 397352 83426 397361
rect 83370 397287 83426 397296
rect 85026 397352 85082 397361
rect 85488 397326 85540 397332
rect 87602 397352 87658 397361
rect 85026 397287 85082 397296
rect 87602 397287 87658 397296
rect 88798 397352 88854 397361
rect 88798 397287 88854 397296
rect 90730 397352 90786 397361
rect 90730 397287 90786 397296
rect 91282 397352 91338 397361
rect 91282 397287 91338 397296
rect 61476 397258 61528 397264
rect 61488 248414 61516 397258
rect 77206 396808 77262 396817
rect 77206 396743 77262 396752
rect 77114 396672 77170 396681
rect 77114 396607 77170 396616
rect 77128 249150 77156 396607
rect 77116 249144 77168 249150
rect 77116 249086 77168 249092
rect 61488 248386 61792 248414
rect 60002 232520 60058 232529
rect 60002 232455 60058 232464
rect 59820 227792 59872 227798
rect 59820 227734 59872 227740
rect 59832 226658 59860 227734
rect 59832 226630 60490 226658
rect 61106 226128 61162 226137
rect 61162 226086 61410 226114
rect 61106 226063 61162 226072
rect 61764 226001 61792 248386
rect 75828 241596 75880 241602
rect 75828 241538 75880 241544
rect 72332 241528 72384 241534
rect 72332 241470 72384 241476
rect 70306 233472 70362 233481
rect 70306 233407 70362 233416
rect 67546 233336 67602 233345
rect 67546 233271 67602 233280
rect 64602 232112 64658 232121
rect 64602 232047 64658 232056
rect 63314 230616 63370 230625
rect 63314 230551 63370 230560
rect 63328 226644 63356 230551
rect 64616 226658 64644 232047
rect 66166 229120 66222 229129
rect 66166 229055 66222 229064
rect 64262 226630 64644 226658
rect 66180 226644 66208 229055
rect 67560 226658 67588 233271
rect 69018 229256 69074 229265
rect 69018 229191 69074 229200
rect 68006 227760 68062 227769
rect 68006 227695 68062 227704
rect 67114 226630 67588 226658
rect 68020 226644 68048 227695
rect 69032 226644 69060 229191
rect 70320 226658 70348 233407
rect 72344 226658 72372 241470
rect 74170 234696 74226 234705
rect 74170 234631 74226 234640
rect 72790 230752 72846 230761
rect 72790 230687 72846 230696
rect 69966 226630 70348 226658
rect 71898 226630 72372 226658
rect 72804 226644 72832 230687
rect 74184 226658 74212 234631
rect 75734 231976 75790 231985
rect 75734 231911 75790 231920
rect 74998 227488 75054 227497
rect 74998 227423 75054 227432
rect 75012 226658 75040 227423
rect 75748 226658 75776 231911
rect 75840 227497 75868 241538
rect 77220 241058 77248 396743
rect 78324 396370 78352 397287
rect 80992 397050 81020 397287
rect 80980 397044 81032 397050
rect 80980 396986 81032 396992
rect 78770 396808 78826 396817
rect 78770 396743 78826 396752
rect 78312 396364 78364 396370
rect 78312 396306 78364 396312
rect 78588 271924 78640 271930
rect 78588 271866 78640 271872
rect 78496 244316 78548 244322
rect 78496 244258 78548 244264
rect 77208 241052 77260 241058
rect 77208 240994 77260 241000
rect 76930 236056 76986 236065
rect 76930 235991 76986 236000
rect 75826 227488 75882 227497
rect 75826 227423 75882 227432
rect 76944 226658 76972 235991
rect 78508 229094 78536 244258
rect 78048 229066 78536 229094
rect 78048 226658 78076 229066
rect 78600 226658 78628 271866
rect 78784 248414 78812 396743
rect 83384 396098 83412 397287
rect 83372 396092 83424 396098
rect 83372 396034 83424 396040
rect 85040 395350 85068 397287
rect 86866 396808 86922 396817
rect 86866 396743 86922 396752
rect 85028 395344 85080 395350
rect 85028 395286 85080 395292
rect 85488 378208 85540 378214
rect 85488 378150 85540 378156
rect 85396 364404 85448 364410
rect 85396 364346 85448 364352
rect 84108 351960 84160 351966
rect 84108 351902 84160 351908
rect 81348 324352 81400 324358
rect 81348 324294 81400 324300
rect 81256 298172 81308 298178
rect 81256 298114 81308 298120
rect 79968 258120 80020 258126
rect 79968 258062 80020 258068
rect 78784 248386 78904 248414
rect 73738 226630 74212 226658
rect 74750 226630 75040 226658
rect 75670 226630 75776 226658
rect 76590 226630 76972 226658
rect 77602 226630 78076 226658
rect 78522 226630 78628 226658
rect 65430 226536 65486 226545
rect 65182 226494 65430 226522
rect 65430 226471 65486 226480
rect 62118 226400 62174 226409
rect 71134 226400 71190 226409
rect 62174 226358 62330 226386
rect 70886 226358 71134 226386
rect 62118 226335 62174 226344
rect 71134 226335 71190 226344
rect 78876 226001 78904 248386
rect 79980 229094 80008 258062
rect 81268 229094 81296 298114
rect 79888 229066 80008 229094
rect 80808 229066 81296 229094
rect 79888 226658 79916 229066
rect 80808 226658 80836 229066
rect 79442 226630 79916 226658
rect 80454 226630 80836 226658
rect 81360 226644 81388 324294
rect 82728 311908 82780 311914
rect 82728 311850 82780 311856
rect 82740 229094 82768 311850
rect 84120 229094 84148 351902
rect 82648 229066 82768 229094
rect 83752 229066 84148 229094
rect 82648 226658 82676 229066
rect 83752 226658 83780 229066
rect 84566 227488 84622 227497
rect 84566 227423 84622 227432
rect 84580 226658 84608 227423
rect 85408 226658 85436 364346
rect 85500 227497 85528 378150
rect 86776 243636 86828 243642
rect 86776 243578 86828 243584
rect 86788 229094 86816 243578
rect 86880 241126 86908 396743
rect 87616 396506 87644 397287
rect 88812 397186 88840 397287
rect 88800 397180 88852 397186
rect 88800 397122 88852 397128
rect 90744 396982 90772 397287
rect 90732 396976 90784 396982
rect 90732 396918 90784 396924
rect 88338 396808 88394 396817
rect 88338 396743 88394 396752
rect 91006 396808 91062 396817
rect 91006 396743 91062 396752
rect 87604 396500 87656 396506
rect 87604 396442 87656 396448
rect 87604 396092 87656 396098
rect 87604 396034 87656 396040
rect 87616 248130 87644 396034
rect 87604 248124 87656 248130
rect 87604 248066 87656 248072
rect 88248 247716 88300 247722
rect 88248 247658 88300 247664
rect 88156 246492 88208 246498
rect 88156 246434 88208 246440
rect 86868 241120 86920 241126
rect 86868 241062 86920 241068
rect 88168 229094 88196 246434
rect 86512 229066 86816 229094
rect 87432 229066 88196 229094
rect 85486 227488 85542 227497
rect 85486 227423 85542 227432
rect 86512 226658 86540 229066
rect 87432 226658 87460 229066
rect 88260 226658 88288 247658
rect 88352 242214 88380 396743
rect 91020 246906 91048 396743
rect 91296 395486 91324 397287
rect 92400 396574 92428 398103
rect 94226 397352 94282 397361
rect 94226 397287 94282 397296
rect 93674 396808 93730 396817
rect 93674 396743 93730 396752
rect 92388 396568 92440 396574
rect 92388 396510 92440 396516
rect 91284 395480 91336 395486
rect 91284 395422 91336 395428
rect 91008 246900 91060 246906
rect 91008 246842 91060 246848
rect 93584 244996 93636 245002
rect 93584 244938 93636 244944
rect 91008 244928 91060 244934
rect 91008 244870 91060 244876
rect 90916 243840 90968 243846
rect 90916 243782 90968 243788
rect 89628 242276 89680 242282
rect 89628 242218 89680 242224
rect 88340 242208 88392 242214
rect 88340 242150 88392 242156
rect 89640 229094 89668 242218
rect 90928 234614 90956 243782
rect 89456 229066 89668 229094
rect 90376 234586 90956 234614
rect 89456 226658 89484 229066
rect 90376 226658 90404 234586
rect 91020 226658 91048 244870
rect 93492 243704 93544 243710
rect 93492 243646 93544 243652
rect 92388 242752 92440 242758
rect 92388 242694 92440 242700
rect 92400 234614 92428 242694
rect 93504 234614 93532 243646
rect 92216 234586 92428 234614
rect 93136 234586 93532 234614
rect 92216 226658 92244 234586
rect 93136 226658 93164 234586
rect 82294 226630 82676 226658
rect 83306 226630 83780 226658
rect 84226 226630 84608 226658
rect 85146 226630 85436 226658
rect 86158 226630 86540 226658
rect 87078 226630 87460 226658
rect 87998 226630 88288 226658
rect 89010 226630 89484 226658
rect 89930 226630 90404 226658
rect 90850 226630 91048 226658
rect 91862 226630 92244 226658
rect 92782 226630 93164 226658
rect 93596 226658 93624 244938
rect 93688 242418 93716 396743
rect 93766 396672 93822 396681
rect 93766 396607 93822 396616
rect 93676 242412 93728 242418
rect 93676 242354 93728 242360
rect 93780 241262 93808 396607
rect 94240 396438 94268 397287
rect 94504 397180 94556 397186
rect 94504 397122 94556 397128
rect 94228 396432 94280 396438
rect 94228 396374 94280 396380
rect 94516 249558 94544 397122
rect 95988 396642 96016 398103
rect 97630 397352 97686 397361
rect 97630 397287 97686 397296
rect 96342 396808 96398 396817
rect 96342 396743 96398 396752
rect 96356 396710 96384 396743
rect 96344 396704 96396 396710
rect 96344 396646 96396 396652
rect 97264 396704 97316 396710
rect 97264 396646 97316 396652
rect 95976 396636 96028 396642
rect 95976 396578 96028 396584
rect 94504 249552 94556 249558
rect 94504 249494 94556 249500
rect 97276 248334 97304 396646
rect 97356 396636 97408 396642
rect 97356 396578 97408 396584
rect 97368 249490 97396 396578
rect 97644 396438 97672 397287
rect 99392 397118 99420 398103
rect 100758 397352 100814 397361
rect 100758 397287 100814 397296
rect 102046 397352 102102 397361
rect 102046 397287 102102 397296
rect 104070 397352 104126 397361
rect 104070 397287 104126 397296
rect 106462 397352 106518 397361
rect 106462 397287 106518 397296
rect 109498 397352 109554 397361
rect 109498 397287 109554 397296
rect 111246 397352 111302 397361
rect 111246 397287 111302 397296
rect 112074 397352 112130 397361
rect 112074 397287 112130 397296
rect 99380 397112 99432 397118
rect 99380 397054 99432 397060
rect 99194 396808 99250 396817
rect 99194 396743 99250 396752
rect 97632 396432 97684 396438
rect 97632 396374 97684 396380
rect 97356 249484 97408 249490
rect 97356 249426 97408 249432
rect 99208 249286 99236 396743
rect 99286 396672 99342 396681
rect 99286 396607 99342 396616
rect 99196 249280 99248 249286
rect 99196 249222 99248 249228
rect 99300 249218 99328 396607
rect 100772 396506 100800 397287
rect 101954 396808 102010 396817
rect 101954 396743 102010 396752
rect 100760 396500 100812 396506
rect 100760 396442 100812 396448
rect 99288 249212 99340 249218
rect 99288 249154 99340 249160
rect 97264 248328 97316 248334
rect 97264 248270 97316 248276
rect 101968 248062 101996 396743
rect 102060 396642 102088 397287
rect 104084 397118 104112 397287
rect 106476 397186 106504 397287
rect 109512 397254 109540 397287
rect 111260 397254 111288 397287
rect 109500 397248 109552 397254
rect 109500 397190 109552 397196
rect 111248 397248 111300 397254
rect 111248 397190 111300 397196
rect 106464 397180 106516 397186
rect 106464 397122 106516 397128
rect 104072 397112 104124 397118
rect 104072 397054 104124 397060
rect 112088 396914 112116 397287
rect 112076 396908 112128 396914
rect 112076 396850 112128 396856
rect 103426 396808 103482 396817
rect 103426 396743 103482 396752
rect 104714 396808 104770 396817
rect 104714 396743 104770 396752
rect 105726 396808 105782 396817
rect 105726 396743 105782 396752
rect 106094 396808 106150 396817
rect 106094 396743 106150 396752
rect 107566 396808 107622 396817
rect 107566 396743 107622 396752
rect 108946 396808 109002 396817
rect 108946 396743 109002 396752
rect 111706 396808 111762 396817
rect 111706 396743 111762 396752
rect 102048 396636 102100 396642
rect 102048 396578 102100 396584
rect 101956 248056 102008 248062
rect 101956 247998 102008 248004
rect 100668 246628 100720 246634
rect 100668 246570 100720 246576
rect 99288 245064 99340 245070
rect 99288 245006 99340 245012
rect 96528 243908 96580 243914
rect 96528 243850 96580 243856
rect 96436 243568 96488 243574
rect 96436 243510 96488 243516
rect 95148 243364 95200 243370
rect 95148 243306 95200 243312
rect 93768 241256 93820 241262
rect 93768 241198 93820 241204
rect 95160 226658 95188 243306
rect 96448 234614 96476 243510
rect 96356 234586 96476 234614
rect 95974 230344 96030 230353
rect 95974 230279 96030 230288
rect 95988 226658 96016 230279
rect 93596 226630 93702 226658
rect 94714 226630 95188 226658
rect 95634 226630 96016 226658
rect 96356 226658 96384 234586
rect 96540 230353 96568 243850
rect 97908 243432 97960 243438
rect 97908 243374 97960 243380
rect 96526 230344 96582 230353
rect 96526 230279 96582 230288
rect 97920 226658 97948 243374
rect 99300 234614 99328 245006
rect 100576 242616 100628 242622
rect 100576 242558 100628 242564
rect 98840 234586 99328 234614
rect 98840 226658 98868 234586
rect 99654 230344 99710 230353
rect 99654 230279 99710 230288
rect 99668 226658 99696 230279
rect 100588 226658 100616 242558
rect 100680 230353 100708 246570
rect 103336 246560 103388 246566
rect 103336 246502 103388 246508
rect 102048 243976 102100 243982
rect 102048 243918 102100 243924
rect 102060 234614 102088 243918
rect 103244 242820 103296 242826
rect 103244 242762 103296 242768
rect 103256 234614 103284 242762
rect 101784 234586 102088 234614
rect 103164 234586 103284 234614
rect 100666 230344 100722 230353
rect 100666 230279 100722 230288
rect 101784 226658 101812 234586
rect 102230 228984 102286 228993
rect 102230 228919 102286 228928
rect 96356 226630 96554 226658
rect 97566 226630 97948 226658
rect 98486 226630 98868 226658
rect 99406 226630 99696 226658
rect 100418 226630 100616 226658
rect 101338 226630 101812 226658
rect 102244 226644 102272 228919
rect 103164 226658 103192 234586
rect 103348 228993 103376 246502
rect 103440 241330 103468 396743
rect 104728 261526 104756 396743
rect 105740 396710 105768 396743
rect 105728 396704 105780 396710
rect 105728 396646 105780 396652
rect 104716 261520 104768 261526
rect 104716 261462 104768 261468
rect 106108 245478 106136 396743
rect 106924 396432 106976 396438
rect 106924 396374 106976 396380
rect 106936 248198 106964 396374
rect 107476 258732 107528 258738
rect 107476 258674 107528 258680
rect 106924 248192 106976 248198
rect 106924 248134 106976 248140
rect 106188 246356 106240 246362
rect 106188 246298 106240 246304
rect 106096 245472 106148 245478
rect 106096 245414 106148 245420
rect 104808 245132 104860 245138
rect 104808 245074 104860 245080
rect 103428 241324 103480 241330
rect 103428 241266 103480 241272
rect 104820 234614 104848 245074
rect 106096 242208 106148 242214
rect 106096 242150 106148 242156
rect 104544 234586 104848 234614
rect 103334 228984 103390 228993
rect 103334 228919 103390 228928
rect 104544 226658 104572 234586
rect 105358 230344 105414 230353
rect 105358 230279 105414 230288
rect 105372 226658 105400 230279
rect 103164 226630 103270 226658
rect 104190 226630 104572 226658
rect 105110 226630 105400 226658
rect 106108 226644 106136 242150
rect 106200 230353 106228 246298
rect 106924 240168 106976 240174
rect 106924 240110 106976 240116
rect 106936 233889 106964 240110
rect 106922 233880 106978 233889
rect 106922 233815 106978 233824
rect 106186 230344 106242 230353
rect 106186 230279 106242 230288
rect 107488 226658 107516 258674
rect 107580 241466 107608 396743
rect 108304 396704 108356 396710
rect 108304 396646 108356 396652
rect 108854 396672 108910 396681
rect 108316 249422 108344 396646
rect 108854 396607 108910 396616
rect 108304 249416 108356 249422
rect 108304 249358 108356 249364
rect 108868 246974 108896 396607
rect 108856 246968 108908 246974
rect 108856 246910 108908 246916
rect 108856 246696 108908 246702
rect 108856 246638 108908 246644
rect 108764 243772 108816 243778
rect 108764 243714 108816 243720
rect 107568 241460 107620 241466
rect 107568 241402 107620 241408
rect 108776 231169 108804 243714
rect 108762 231160 108818 231169
rect 108762 231095 108818 231104
rect 108868 228993 108896 246638
rect 108960 240718 108988 396743
rect 111720 248266 111748 396743
rect 112996 258800 113048 258806
rect 112996 258742 113048 258748
rect 111708 248260 111760 248266
rect 111708 248202 111760 248208
rect 111708 246424 111760 246430
rect 111708 246366 111760 246372
rect 110328 245200 110380 245206
rect 110328 245142 110380 245148
rect 108948 240712 109000 240718
rect 108948 240654 109000 240660
rect 108946 231160 109002 231169
rect 108946 231095 109002 231104
rect 107934 228984 107990 228993
rect 107934 228919 107990 228928
rect 108854 228984 108910 228993
rect 108854 228919 108910 228928
rect 107042 226630 107516 226658
rect 107948 226644 107976 228919
rect 108960 226644 108988 231095
rect 110340 229094 110368 245142
rect 111720 229094 111748 246366
rect 113008 229094 113036 258742
rect 110248 229066 110368 229094
rect 111168 229066 111748 229094
rect 112272 229066 113036 229094
rect 110248 226658 110276 229066
rect 111168 226658 111196 229066
rect 112272 226658 112300 229066
rect 113100 226658 113128 399706
rect 113638 398168 113694 398177
rect 113638 398103 113694 398112
rect 113178 397352 113234 397361
rect 113178 397287 113234 397296
rect 113192 396846 113220 397287
rect 113652 397118 113680 398103
rect 113730 397352 113786 397361
rect 113730 397287 113786 397296
rect 113640 397112 113692 397118
rect 113640 397054 113692 397060
rect 113180 396840 113232 396846
rect 113180 396782 113232 396788
rect 113744 396778 113772 397287
rect 113732 396772 113784 396778
rect 113732 396714 113784 396720
rect 115768 393314 115796 399842
rect 119988 399832 120040 399838
rect 119988 399774 120040 399780
rect 115846 397352 115902 397361
rect 115846 397287 115902 397296
rect 117134 397352 117190 397361
rect 117134 397287 117190 397296
rect 118330 397352 118386 397361
rect 118330 397287 118386 397296
rect 118606 397352 118662 397361
rect 118606 397287 118662 397296
rect 115860 396914 115888 397287
rect 115848 396908 115900 396914
rect 115848 396850 115900 396856
rect 117042 396808 117098 396817
rect 117148 396778 117176 397287
rect 118344 396846 118372 397287
rect 118332 396840 118384 396846
rect 118332 396782 118384 396788
rect 117042 396743 117098 396752
rect 117136 396772 117188 396778
rect 115768 393286 115888 393314
rect 115756 243024 115808 243030
rect 115756 242966 115808 242972
rect 114468 242072 114520 242078
rect 114468 242014 114520 242020
rect 114480 229094 114508 242014
rect 115768 229094 115796 242966
rect 114112 229066 114508 229094
rect 115032 229066 115796 229094
rect 114112 226658 114140 229066
rect 115032 226658 115060 229066
rect 115860 226658 115888 393286
rect 117056 242894 117084 396743
rect 117136 396714 117188 396720
rect 118620 395622 118648 397287
rect 119894 396808 119950 396817
rect 119894 396743 119950 396752
rect 118608 395616 118660 395622
rect 118608 395558 118660 395564
rect 119908 249354 119936 396743
rect 119896 249348 119948 249354
rect 119896 249290 119948 249296
rect 117136 244724 117188 244730
rect 117136 244666 117188 244672
rect 117044 242888 117096 242894
rect 117044 242830 117096 242836
rect 117148 229094 117176 244666
rect 118608 243092 118660 243098
rect 118608 243034 118660 243040
rect 118516 242004 118568 242010
rect 118516 241946 118568 241952
rect 118528 229094 118556 241946
rect 116872 229066 117176 229094
rect 117976 229066 118556 229094
rect 116872 226658 116900 229066
rect 117976 226658 118004 229066
rect 118620 226658 118648 243034
rect 120000 234614 120028 399774
rect 122932 399560 122984 399566
rect 122932 399502 122984 399508
rect 122748 398132 122800 398138
rect 122748 398074 122800 398080
rect 120078 396808 120134 396817
rect 120078 396743 120134 396752
rect 120092 246022 120120 396743
rect 120724 247648 120776 247654
rect 120724 247590 120776 247596
rect 120080 246016 120132 246022
rect 120080 245958 120132 245964
rect 119816 234586 120028 234614
rect 119816 226658 119844 234586
rect 120736 226658 120764 247590
rect 121274 237960 121330 237969
rect 121274 237895 121330 237904
rect 109894 226630 110276 226658
rect 110814 226630 111196 226658
rect 111826 226630 112300 226658
rect 112746 226630 113128 226658
rect 113666 226630 114140 226658
rect 114678 226630 115060 226658
rect 115598 226630 115888 226658
rect 116518 226630 116900 226658
rect 117530 226630 118004 226658
rect 118450 226630 118648 226658
rect 119370 226630 119844 226658
rect 120382 226630 120764 226658
rect 121288 226644 121316 237895
rect 122760 234614 122788 398074
rect 122944 248414 122972 399502
rect 169668 398200 169720 398206
rect 146022 398168 146078 398177
rect 169668 398142 169720 398148
rect 146022 398103 146078 398112
rect 143540 397520 143592 397526
rect 143540 397462 143592 397468
rect 123482 397352 123538 397361
rect 123482 397287 123538 397296
rect 125966 397352 126022 397361
rect 125966 397287 126022 397296
rect 136270 397352 136326 397361
rect 136270 397287 136326 397296
rect 138386 397352 138442 397361
rect 138386 397287 138442 397296
rect 123496 395418 123524 397287
rect 125980 395418 126008 397287
rect 134524 397180 134576 397186
rect 134524 397122 134576 397128
rect 129738 396808 129794 396817
rect 129738 396743 129794 396752
rect 133786 396808 133842 396817
rect 133786 396743 133842 396752
rect 129646 396128 129702 396137
rect 129646 396063 129702 396072
rect 123484 395412 123536 395418
rect 123484 395354 123536 395360
rect 125968 395412 126020 395418
rect 125968 395354 126020 395360
rect 122944 248386 123800 248414
rect 122576 234586 122788 234614
rect 122576 226658 122604 234586
rect 123206 228440 123262 228449
rect 123206 228375 123262 228384
rect 122222 226630 122604 226658
rect 123220 226644 123248 228375
rect 123772 226658 123800 248386
rect 126980 246220 127032 246226
rect 126980 246162 127032 246168
rect 125600 243160 125652 243166
rect 125600 243102 125652 243108
rect 125046 232520 125102 232529
rect 125046 232455 125102 232464
rect 123772 226630 124154 226658
rect 125060 226644 125088 232455
rect 125612 226658 125640 243102
rect 126992 230353 127020 246162
rect 127072 245540 127124 245546
rect 127072 245482 127124 245488
rect 127084 234614 127112 245482
rect 128544 244248 128596 244254
rect 128544 244190 128596 244196
rect 127084 234586 127204 234614
rect 126978 230344 127034 230353
rect 126978 230279 127034 230288
rect 127176 226658 127204 234586
rect 127530 230344 127586 230353
rect 127530 230279 127586 230288
rect 125612 226630 126086 226658
rect 127006 226630 127204 226658
rect 127544 226658 127572 230279
rect 128556 226658 128584 244190
rect 129660 242146 129688 396063
rect 129752 248402 129780 396743
rect 129740 248396 129792 248402
rect 129740 248338 129792 248344
rect 133800 246294 133828 396743
rect 132500 246288 132552 246294
rect 132500 246230 132552 246236
rect 133788 246288 133840 246294
rect 133788 246230 133840 246236
rect 129740 246152 129792 246158
rect 129740 246094 129792 246100
rect 129648 242140 129700 242146
rect 129648 242082 129700 242088
rect 129752 234025 129780 246094
rect 129832 245608 129884 245614
rect 129832 245550 129884 245556
rect 129738 234016 129794 234025
rect 129738 233951 129794 233960
rect 127544 226630 127926 226658
rect 128556 226630 128938 226658
rect 129844 226644 129872 245550
rect 131304 242548 131356 242554
rect 131304 242490 131356 242496
rect 130382 234016 130438 234025
rect 130382 233951 130438 233960
rect 130396 226658 130424 233951
rect 131316 226658 131344 242490
rect 132512 234025 132540 246230
rect 134536 245546 134564 397122
rect 136284 395486 136312 397287
rect 137284 397248 137336 397254
rect 137284 397190 137336 397196
rect 136272 395480 136324 395486
rect 136272 395422 136324 395428
rect 137296 246226 137324 397190
rect 138400 395554 138428 397287
rect 142804 397044 142856 397050
rect 142804 396986 142856 396992
rect 140778 396808 140834 396817
rect 140778 396743 140834 396752
rect 138388 395548 138440 395554
rect 138388 395490 138440 395496
rect 137284 246220 137336 246226
rect 137284 246162 137336 246168
rect 140792 246090 140820 396743
rect 142816 267734 142844 396986
rect 142816 267706 142936 267734
rect 142804 256760 142856 256766
rect 142804 256702 142856 256708
rect 142816 251802 142844 256702
rect 141424 251796 141476 251802
rect 141424 251738 141476 251744
rect 142804 251796 142856 251802
rect 142804 251738 142856 251744
rect 140872 247036 140924 247042
rect 140872 246978 140924 246984
rect 140780 246084 140832 246090
rect 140780 246026 140832 246032
rect 138572 245608 138624 245614
rect 138572 245550 138624 245556
rect 134524 245540 134576 245546
rect 134524 245482 134576 245488
rect 138112 245336 138164 245342
rect 138112 245278 138164 245284
rect 132592 244860 132644 244866
rect 132592 244802 132644 244808
rect 132498 234016 132554 234025
rect 132498 233951 132554 233960
rect 132604 226658 132632 244802
rect 135260 244792 135312 244798
rect 135260 244734 135312 244740
rect 134248 243500 134300 243506
rect 134248 243442 134300 243448
rect 133142 234016 133198 234025
rect 133142 233951 133198 233960
rect 133156 226658 133184 233951
rect 134260 226658 134288 243442
rect 135272 226658 135300 244734
rect 138020 244588 138072 244594
rect 138020 244530 138072 244536
rect 137008 244180 137060 244186
rect 137008 244122 137060 244128
rect 135904 243500 135956 243506
rect 135904 243442 135956 243448
rect 135352 243228 135404 243234
rect 135352 243170 135404 243176
rect 135364 229094 135392 243170
rect 135916 237969 135944 243442
rect 135902 237960 135958 237969
rect 135902 237895 135958 237904
rect 135364 229066 136128 229094
rect 136100 226658 136128 229066
rect 137020 226658 137048 244122
rect 138032 227497 138060 244530
rect 138018 227488 138074 227497
rect 138018 227423 138074 227432
rect 138124 226658 138152 245278
rect 138584 243506 138612 245550
rect 139952 244112 140004 244118
rect 139952 244054 140004 244060
rect 138572 243500 138624 243506
rect 138572 243442 138624 243448
rect 138938 227488 138994 227497
rect 138938 227423 138994 227432
rect 138952 226658 138980 227423
rect 139964 226658 139992 244054
rect 140884 226658 140912 246978
rect 141436 245682 141464 251738
rect 142908 249626 142936 267706
rect 142896 249620 142948 249626
rect 142896 249562 142948 249568
rect 143552 248414 143580 397462
rect 144826 396808 144882 396817
rect 144826 396743 144882 396752
rect 144184 262948 144236 262954
rect 144184 262890 144236 262896
rect 144196 256766 144224 262890
rect 144184 256760 144236 256766
rect 144184 256702 144236 256708
rect 143552 248386 143672 248414
rect 142160 247988 142212 247994
rect 142160 247930 142212 247936
rect 141424 245676 141476 245682
rect 141424 245618 141476 245624
rect 130396 226630 130778 226658
rect 131316 226630 131790 226658
rect 132604 226630 132710 226658
rect 133156 226630 133630 226658
rect 134260 226630 134642 226658
rect 135272 226630 135562 226658
rect 136100 226630 136482 226658
rect 137020 226630 137494 226658
rect 138124 226630 138414 226658
rect 138952 226630 139334 226658
rect 139964 226630 140346 226658
rect 140884 226630 141266 226658
rect 142172 226644 142200 247930
rect 142712 245404 142764 245410
rect 142712 245346 142764 245352
rect 142724 226658 142752 245346
rect 143644 226658 143672 248386
rect 144840 241942 144868 396743
rect 146036 395758 146064 398103
rect 156418 397352 156474 397361
rect 156418 397287 156474 397296
rect 163870 397352 163926 397361
rect 163870 397287 163926 397296
rect 147678 396808 147734 396817
rect 147678 396743 147734 396752
rect 151726 396808 151782 396817
rect 151726 396743 151782 396752
rect 154486 396808 154542 396817
rect 154486 396743 154542 396752
rect 146024 395752 146076 395758
rect 146024 395694 146076 395700
rect 144920 371272 144972 371278
rect 144920 371214 144972 371220
rect 144828 241936 144880 241942
rect 144828 241878 144880 241884
rect 144932 227497 144960 371214
rect 147692 358086 147720 396743
rect 147680 358080 147732 358086
rect 147680 358022 147732 358028
rect 147680 357468 147732 357474
rect 147680 357410 147732 357416
rect 146300 345092 146352 345098
rect 146300 345034 146352 345040
rect 145564 266416 145616 266422
rect 145564 266358 145616 266364
rect 145576 262954 145604 266358
rect 145564 262948 145616 262954
rect 145564 262890 145616 262896
rect 146312 248414 146340 345034
rect 146944 271244 146996 271250
rect 146944 271186 146996 271192
rect 146956 266422 146984 271186
rect 146944 266416 146996 266422
rect 146944 266358 146996 266364
rect 146312 248386 146616 248414
rect 145012 244656 145064 244662
rect 145012 244598 145064 244604
rect 144918 227488 144974 227497
rect 144918 227423 144974 227432
rect 142724 226630 143198 226658
rect 143644 226630 144118 226658
rect 145024 226644 145052 244598
rect 145746 227488 145802 227497
rect 145746 227423 145802 227432
rect 145760 226658 145788 227423
rect 146588 226658 146616 248386
rect 147692 226658 147720 357410
rect 147772 318844 147824 318850
rect 147772 318786 147824 318792
rect 147784 248414 147812 318786
rect 151084 306400 151136 306406
rect 151084 306342 151136 306348
rect 150440 305040 150492 305046
rect 150440 304982 150492 304988
rect 149704 299464 149756 299470
rect 149704 299406 149756 299412
rect 149060 292596 149112 292602
rect 149060 292538 149112 292544
rect 148324 282940 148376 282946
rect 148324 282882 148376 282888
rect 148336 271250 148364 282882
rect 148324 271244 148376 271250
rect 148324 271186 148376 271192
rect 149072 248414 149100 292538
rect 149716 282946 149744 299406
rect 149704 282940 149756 282946
rect 149704 282882 149756 282888
rect 147784 248386 148456 248414
rect 149072 248386 149376 248414
rect 148428 226658 148456 248386
rect 149348 226658 149376 248386
rect 150452 226658 150480 304982
rect 151096 299470 151124 306342
rect 151084 299464 151136 299470
rect 151084 299406 151136 299412
rect 151740 267034 151768 396743
rect 154500 367810 154528 396743
rect 156432 395894 156460 397287
rect 158626 396808 158682 396817
rect 158626 396743 158682 396752
rect 161386 396808 161442 396817
rect 161386 396743 161442 396752
rect 156420 395888 156472 395894
rect 156420 395830 156472 395836
rect 154488 367804 154540 367810
rect 154488 367746 154540 367752
rect 156604 346384 156656 346390
rect 156604 346326 156656 346332
rect 156616 311982 156644 346326
rect 154580 311976 154632 311982
rect 154580 311918 154632 311924
rect 156604 311976 156656 311982
rect 156604 311918 156656 311924
rect 154592 310570 154620 311918
rect 154500 310542 154620 310570
rect 154500 306406 154528 310542
rect 154488 306400 154540 306406
rect 154488 306342 154540 306348
rect 151728 267028 151780 267034
rect 151728 266970 151780 266976
rect 150532 266484 150584 266490
rect 150532 266426 150584 266432
rect 150544 248414 150572 266426
rect 153200 253972 153252 253978
rect 153200 253914 153252 253920
rect 150544 248386 151400 248414
rect 151372 226658 151400 248386
rect 152278 233880 152334 233889
rect 152278 233815 152334 233824
rect 152292 226658 152320 233815
rect 153212 226658 153240 253914
rect 158640 244254 158668 396743
rect 160100 359508 160152 359514
rect 160100 359450 160152 359456
rect 160112 357474 160140 359450
rect 159364 357468 159416 357474
rect 159364 357410 159416 357416
rect 160100 357468 160152 357474
rect 160100 357410 160152 357416
rect 159376 346390 159404 357410
rect 159364 346384 159416 346390
rect 159364 346326 159416 346332
rect 161400 247042 161428 396743
rect 163884 395962 163912 397287
rect 165618 396808 165674 396817
rect 165618 396743 165674 396752
rect 163872 395956 163924 395962
rect 163872 395898 163924 395904
rect 164884 372564 164936 372570
rect 164884 372506 164936 372512
rect 164896 359514 164924 372506
rect 164884 359508 164936 359514
rect 164884 359450 164936 359456
rect 161388 247036 161440 247042
rect 161388 246978 161440 246984
rect 158628 244248 158680 244254
rect 158628 244190 158680 244196
rect 165632 243302 165660 396743
rect 165620 243296 165672 243302
rect 165620 243238 165672 243244
rect 167366 234832 167422 234841
rect 167366 234767 167422 234776
rect 157982 232384 158038 232393
rect 157982 232319 158038 232328
rect 157430 229528 157486 229537
rect 157430 229463 157486 229472
rect 154578 229392 154634 229401
rect 154578 229327 154634 229336
rect 145760 226630 146050 226658
rect 146588 226630 146970 226658
rect 147692 226630 147890 226658
rect 148428 226630 148902 226658
rect 149348 226630 149822 226658
rect 150452 226630 150742 226658
rect 151372 226630 151754 226658
rect 152292 226630 152674 226658
rect 153212 226630 153594 226658
rect 154592 226644 154620 229327
rect 156602 227896 156658 227905
rect 156602 227831 156658 227840
rect 156616 226953 156644 227831
rect 156602 226944 156658 226953
rect 156602 226879 156658 226888
rect 156418 226808 156474 226817
rect 156418 226743 156474 226752
rect 155130 226672 155186 226681
rect 155186 226630 155526 226658
rect 156432 226644 156460 226743
rect 157444 226644 157472 229463
rect 157996 226658 158024 232319
rect 160742 232248 160798 232257
rect 160742 232183 160798 232192
rect 160282 230888 160338 230897
rect 160282 230823 160338 230832
rect 159270 228576 159326 228585
rect 159270 228511 159326 228520
rect 157996 226630 158378 226658
rect 159284 226644 159312 228511
rect 160296 226644 160324 230823
rect 160756 226658 160784 232183
rect 165986 231024 166042 231033
rect 165986 230959 166042 230968
rect 163134 229664 163190 229673
rect 163134 229599 163190 229608
rect 162122 228032 162178 228041
rect 162122 227967 162178 227976
rect 160756 226630 161230 226658
rect 162136 226644 162164 227967
rect 163148 226644 163176 229599
rect 164054 228304 164110 228313
rect 164054 228239 164110 228248
rect 164068 226644 164096 228239
rect 164974 228168 165030 228177
rect 164974 228103 165030 228112
rect 164988 226644 165016 228103
rect 166000 226644 166028 230959
rect 166906 227896 166962 227905
rect 166906 227831 166962 227840
rect 166920 226644 166948 227831
rect 167380 226658 167408 234767
rect 169680 229094 169708 398142
rect 170404 397112 170456 397118
rect 170404 397054 170456 397060
rect 169760 242684 169812 242690
rect 169760 242626 169812 242632
rect 169312 229066 169708 229094
rect 169312 226658 169340 229066
rect 167380 226630 167854 226658
rect 168866 226630 169340 226658
rect 169772 226644 169800 242626
rect 170416 242554 170444 397054
rect 173808 397044 173860 397050
rect 173808 396986 173860 396992
rect 171140 375148 171192 375154
rect 171140 375090 171192 375096
rect 171152 372638 171180 375090
rect 171140 372632 171192 372638
rect 171140 372574 171192 372580
rect 171232 248124 171284 248130
rect 171232 248066 171284 248072
rect 170404 242548 170456 242554
rect 170404 242490 170456 242496
rect 170678 228304 170734 228313
rect 170678 228239 170734 228248
rect 170692 226644 170720 228239
rect 171244 226658 171272 248066
rect 173716 244384 173768 244390
rect 173716 244326 173768 244332
rect 172886 226672 172942 226681
rect 171244 226630 171718 226658
rect 172638 226630 172886 226658
rect 155130 226607 155186 226616
rect 173728 226658 173756 244326
rect 173820 226681 173848 396986
rect 175280 377052 175332 377058
rect 175280 376994 175332 377000
rect 175292 375154 175320 376994
rect 175280 375148 175332 375154
rect 175280 375090 175332 375096
rect 176016 248328 176068 248334
rect 176016 248270 176068 248276
rect 174542 228440 174598 228449
rect 174542 228375 174598 228384
rect 173558 226630 173756 226658
rect 173806 226672 173862 226681
rect 172886 226607 172942 226616
rect 174556 226644 174584 228375
rect 175830 227488 175886 227497
rect 175830 227423 175886 227432
rect 175844 226658 175872 227423
rect 175490 226630 175872 226658
rect 176028 226658 176056 248270
rect 176580 227497 176608 399978
rect 184204 399968 184256 399974
rect 184204 399910 184256 399916
rect 180708 399560 180760 399566
rect 180708 399502 180760 399508
rect 177948 398268 178000 398274
rect 177948 398210 178000 398216
rect 177304 397180 177356 397186
rect 177304 397122 177356 397128
rect 177316 244390 177344 397122
rect 177396 388544 177448 388550
rect 177396 388486 177448 388492
rect 177408 377058 177436 388486
rect 177396 377052 177448 377058
rect 177396 376994 177448 377000
rect 177304 244384 177356 244390
rect 177304 244326 177356 244332
rect 177960 229094 177988 398210
rect 179328 395820 179380 395826
rect 179328 395762 179380 395768
rect 179340 229094 179368 395762
rect 180524 393372 180576 393378
rect 180524 393314 180576 393320
rect 180536 388550 180564 393314
rect 180524 388544 180576 388550
rect 180524 388486 180576 388492
rect 177776 229066 177988 229094
rect 178696 229066 179368 229094
rect 176566 227488 176622 227497
rect 176566 227423 176622 227432
rect 177776 226658 177804 229066
rect 178696 226658 178724 229066
rect 179234 228576 179290 228585
rect 179234 228511 179290 228520
rect 176028 226630 176410 226658
rect 177422 226630 177804 226658
rect 178342 226630 178724 226658
rect 179248 226644 179276 228511
rect 180720 226658 180748 399502
rect 182178 396808 182234 396817
rect 182178 396743 182234 396752
rect 183466 396808 183522 396817
rect 183466 396743 183522 396752
rect 180892 249552 180944 249558
rect 180892 249494 180944 249500
rect 180904 226681 180932 249494
rect 182192 241482 182220 396743
rect 183284 395548 183336 395554
rect 183284 395490 183336 395496
rect 183296 393378 183324 395490
rect 183284 393372 183336 393378
rect 183284 393314 183336 393320
rect 183480 245614 183508 396743
rect 183468 245608 183520 245614
rect 183468 245550 183520 245556
rect 183560 242480 183612 242486
rect 183560 242422 183612 242428
rect 182008 241454 182220 241482
rect 182008 241398 182036 241454
rect 181996 241392 182048 241398
rect 181996 241334 182048 241340
rect 182088 241392 182140 241398
rect 182088 241334 182140 241340
rect 182100 229094 182128 241334
rect 181640 229066 182128 229094
rect 180274 226630 180748 226658
rect 180890 226672 180946 226681
rect 173806 226607 173862 226616
rect 181640 226658 181668 229066
rect 183098 227896 183154 227905
rect 183098 227831 183154 227840
rect 181194 226630 181668 226658
rect 181810 226672 181866 226681
rect 180890 226607 180946 226616
rect 181866 226630 182114 226658
rect 183112 226644 183140 227831
rect 183572 226658 183600 242422
rect 184216 227905 184244 399910
rect 185584 398336 185636 398342
rect 185584 398278 185636 398284
rect 184296 397112 184348 397118
rect 184296 397054 184348 397060
rect 184308 241398 184336 397054
rect 185596 395554 185624 398278
rect 185584 395548 185636 395554
rect 185584 395490 185636 395496
rect 186228 245336 186280 245342
rect 186228 245278 186280 245284
rect 184296 241392 184348 241398
rect 184296 241334 184348 241340
rect 184938 228712 184994 228721
rect 184938 228647 184994 228656
rect 184202 227896 184258 227905
rect 184202 227831 184258 227840
rect 183572 226630 184046 226658
rect 184952 226644 184980 228647
rect 186240 226658 186268 245278
rect 187620 229094 187648 399978
rect 187792 396976 187844 396982
rect 187792 396918 187844 396924
rect 187344 229066 187648 229094
rect 187344 226658 187372 229066
rect 185978 226630 186268 226658
rect 186898 226630 187372 226658
rect 187804 226644 187832 396918
rect 191748 395684 191800 395690
rect 191748 395626 191800 395632
rect 188988 247988 189040 247994
rect 188988 247930 189040 247936
rect 189000 226658 189028 247930
rect 190368 241392 190420 241398
rect 190368 241334 190420 241340
rect 190380 229094 190408 241334
rect 191760 229094 191788 395626
rect 195888 395548 195940 395554
rect 195888 395490 195940 395496
rect 193220 248260 193272 248266
rect 193220 248202 193272 248208
rect 193128 248124 193180 248130
rect 193128 248066 193180 248072
rect 193140 229094 193168 248066
rect 190104 229066 190408 229094
rect 191024 229066 191788 229094
rect 193048 229066 193168 229094
rect 190104 226658 190132 229066
rect 191024 226658 191052 229066
rect 191654 227896 191710 227905
rect 191654 227831 191710 227840
rect 188830 226630 189028 226658
rect 189750 226630 190132 226658
rect 190670 226630 191052 226658
rect 191668 226644 191696 227831
rect 193048 226658 193076 229066
rect 192602 226630 193076 226658
rect 193232 226658 193260 248202
rect 194048 242548 194100 242554
rect 194048 242490 194100 242496
rect 194060 226658 194088 242490
rect 195900 229094 195928 395490
rect 195980 249484 196032 249490
rect 195980 249426 196032 249432
rect 195808 229066 195928 229094
rect 195808 226658 195836 229066
rect 193232 226630 193522 226658
rect 194060 226630 194534 226658
rect 195454 226630 195836 226658
rect 195992 226658 196020 249426
rect 196544 247654 196572 486118
rect 196716 483880 196768 483886
rect 196636 483828 196716 483834
rect 196636 483822 196768 483828
rect 196636 483806 196756 483822
rect 196636 398138 196664 483806
rect 196820 483698 196848 488506
rect 196728 483670 196848 483698
rect 196624 398132 196676 398138
rect 196624 398074 196676 398080
rect 196624 396976 196676 396982
rect 196624 396918 196676 396924
rect 196532 247648 196584 247654
rect 196532 247590 196584 247596
rect 196636 241398 196664 396918
rect 196624 241392 196676 241398
rect 196624 241334 196676 241340
rect 196728 228449 196756 483670
rect 197004 478874 197032 489886
rect 196820 478846 197032 478874
rect 196820 398342 196848 478846
rect 196808 398336 196860 398342
rect 196808 398278 196860 398284
rect 197372 228585 197400 504630
rect 197358 228576 197414 228585
rect 197358 228511 197414 228520
rect 196714 228440 196770 228449
rect 196714 228375 196770 228384
rect 197464 227905 197492 504834
rect 197542 413672 197598 413681
rect 197542 413607 197598 413616
rect 197556 400110 197584 413607
rect 197544 400104 197596 400110
rect 197544 400046 197596 400052
rect 197544 395616 197596 395622
rect 197544 395558 197596 395564
rect 197450 227896 197506 227905
rect 197450 227831 197506 227840
rect 197556 226658 197584 395558
rect 198016 243030 198044 700470
rect 200212 503532 200264 503538
rect 200212 503474 200264 503480
rect 200764 503532 200816 503538
rect 200764 503474 200816 503480
rect 198738 479224 198794 479233
rect 198738 479159 198794 479168
rect 198004 243024 198056 243030
rect 198004 242966 198056 242972
rect 198648 241392 198700 241398
rect 198648 241334 198700 241340
rect 198660 226658 198688 241334
rect 198752 241194 198780 479159
rect 198830 419384 198886 419393
rect 198830 419319 198886 419328
rect 198844 400042 198872 419319
rect 198922 417752 198978 417761
rect 198922 417687 198978 417696
rect 198832 400036 198884 400042
rect 198832 399978 198884 399984
rect 198936 399702 198964 417687
rect 199474 416392 199530 416401
rect 199474 416327 199530 416336
rect 199382 414896 199438 414905
rect 199382 414831 199438 414840
rect 198924 399696 198976 399702
rect 198924 399638 198976 399644
rect 198832 248192 198884 248198
rect 198832 248134 198884 248140
rect 198740 241188 198792 241194
rect 198740 241130 198792 241136
rect 195992 226630 196374 226658
rect 197386 226630 197584 226658
rect 198306 226630 198688 226658
rect 198844 226658 198872 248134
rect 199396 244866 199424 414831
rect 199488 399702 199516 416327
rect 199476 399696 199528 399702
rect 199476 399638 199528 399644
rect 199384 244860 199436 244866
rect 199384 244802 199436 244808
rect 198844 226630 199226 226658
rect 200224 226644 200252 503474
rect 200776 228721 200804 503474
rect 201512 243098 201540 702986
rect 204904 700732 204956 700738
rect 204904 700674 204956 700680
rect 201592 503600 201644 503606
rect 201592 503542 201644 503548
rect 201500 243092 201552 243098
rect 201500 243034 201552 243040
rect 201408 241188 201460 241194
rect 201408 241130 201460 241136
rect 200762 228712 200818 228721
rect 200762 228647 200818 228656
rect 201420 226658 201448 241130
rect 201158 226630 201448 226658
rect 201604 226658 201632 503542
rect 204168 243500 204220 243506
rect 204168 243442 204220 243448
rect 204076 242548 204128 242554
rect 204076 242490 204128 242496
rect 204088 234614 204116 242490
rect 203996 234586 204116 234614
rect 203430 230344 203486 230353
rect 203430 230279 203486 230288
rect 203444 226658 203472 230279
rect 201604 226630 202078 226658
rect 203090 226630 203472 226658
rect 203996 226644 204024 234586
rect 204180 230353 204208 243442
rect 204916 242010 204944 700674
rect 206376 700664 206428 700670
rect 206376 700606 206428 700612
rect 206284 563100 206336 563106
rect 206284 563042 206336 563048
rect 204996 510672 205048 510678
rect 204996 510614 205048 510620
rect 205008 242758 205036 510614
rect 205548 244180 205600 244186
rect 205548 244122 205600 244128
rect 204996 242752 205048 242758
rect 204996 242694 205048 242700
rect 204904 242004 204956 242010
rect 204904 241946 204956 241952
rect 205560 234614 205588 244122
rect 206296 243370 206324 563042
rect 206388 399906 206416 700606
rect 213276 700596 213328 700602
rect 213276 700538 213328 700544
rect 209044 700392 209096 700398
rect 209044 700334 209096 700340
rect 206468 504212 206520 504218
rect 206468 504154 206520 504160
rect 206376 399900 206428 399906
rect 206376 399842 206428 399848
rect 206284 243364 206336 243370
rect 206284 243306 206336 243312
rect 205376 234586 205588 234614
rect 204166 230344 204222 230353
rect 204166 230279 204222 230288
rect 205376 226658 205404 234586
rect 206480 228313 206508 504154
rect 207020 249416 207072 249422
rect 207020 249358 207072 249364
rect 207032 248414 207060 249358
rect 207032 248386 207336 248414
rect 206928 245404 206980 245410
rect 206928 245346 206980 245352
rect 206836 242684 206888 242690
rect 206836 242626 206888 242632
rect 206848 234614 206876 242626
rect 206572 234586 206876 234614
rect 206466 228304 206522 228313
rect 206466 228239 206522 228248
rect 206572 226794 206600 234586
rect 206296 226766 206600 226794
rect 206296 226658 206324 226766
rect 206940 226658 206968 245346
rect 204930 226630 205404 226658
rect 205942 226630 206324 226658
rect 206862 226630 206968 226658
rect 207308 226658 207336 248386
rect 208492 245540 208544 245546
rect 208492 245482 208544 245488
rect 208504 226658 208532 245482
rect 209056 242078 209084 700334
rect 209136 616888 209188 616894
rect 209136 616830 209188 616836
rect 209148 243438 209176 616830
rect 212448 504484 212500 504490
rect 212448 504426 212500 504432
rect 210516 430636 210568 430642
rect 210516 430578 210568 430584
rect 210424 407924 210476 407930
rect 210424 407866 210476 407872
rect 210436 398818 210464 407866
rect 210424 398812 210476 398818
rect 210424 398754 210476 398760
rect 209780 395752 209832 395758
rect 209780 395694 209832 395700
rect 209792 248414 209820 395694
rect 209792 248386 210280 248414
rect 209688 244112 209740 244118
rect 209688 244054 209740 244060
rect 209136 243432 209188 243438
rect 209136 243374 209188 243380
rect 209044 242072 209096 242078
rect 209044 242014 209096 242020
rect 207308 226630 207782 226658
rect 208504 226630 208794 226658
rect 209700 226644 209728 244054
rect 210252 226658 210280 248386
rect 210528 240990 210556 430578
rect 210608 429208 210660 429214
rect 210608 429150 210660 429156
rect 210620 398274 210648 429150
rect 210700 407176 210752 407182
rect 210700 407118 210752 407124
rect 210608 398268 210660 398274
rect 210608 398210 210660 398216
rect 210712 398206 210740 407118
rect 210700 398200 210752 398206
rect 210700 398142 210752 398148
rect 210516 240984 210568 240990
rect 210516 240926 210568 240932
rect 212460 234614 212488 504426
rect 213184 503396 213236 503402
rect 213184 503338 213236 503344
rect 213196 502382 213224 503338
rect 213184 502376 213236 502382
rect 213184 502318 213236 502324
rect 213196 407930 213224 502318
rect 213184 407924 213236 407930
rect 213184 407866 213236 407872
rect 212540 267028 212592 267034
rect 212540 266970 212592 266976
rect 212000 234586 212488 234614
rect 212000 226658 212028 234586
rect 212552 230353 212580 266970
rect 212632 246220 212684 246226
rect 212632 246162 212684 246168
rect 212644 234614 212672 246162
rect 213288 244730 213316 700538
rect 215944 700460 215996 700466
rect 215944 700402 215996 700408
rect 214564 700324 214616 700330
rect 214564 700266 214616 700272
rect 213368 670744 213420 670750
rect 213368 670686 213420 670692
rect 213276 244724 213328 244730
rect 213276 244666 213328 244672
rect 213380 242622 213408 670686
rect 214576 242826 214604 700266
rect 214656 699712 214708 699718
rect 214656 699654 214708 699660
rect 214668 399838 214696 699654
rect 215760 504824 215812 504830
rect 215760 504766 215812 504772
rect 215300 504756 215352 504762
rect 215300 504698 215352 504704
rect 214656 399832 214708 399838
rect 214656 399774 214708 399780
rect 214564 242820 214616 242826
rect 214564 242762 214616 242768
rect 213368 242616 213420 242622
rect 213368 242558 213420 242564
rect 215208 240644 215260 240650
rect 215208 240586 215260 240592
rect 215220 234614 215248 240586
rect 212644 234586 212764 234614
rect 212538 230344 212594 230353
rect 212538 230279 212594 230288
rect 212736 226658 212764 234586
rect 214944 234586 215248 234614
rect 213090 230344 213146 230353
rect 213090 230279 213146 230288
rect 210252 226630 210634 226658
rect 211646 226630 212028 226658
rect 212566 226630 212764 226658
rect 213104 226658 213132 230279
rect 214944 226658 214972 234586
rect 215312 232937 215340 504698
rect 215576 504552 215628 504558
rect 215576 504494 215628 504500
rect 215484 504416 215536 504422
rect 215484 504358 215536 504364
rect 215392 395888 215444 395894
rect 215392 395830 215444 395836
rect 215298 232928 215354 232937
rect 215298 232863 215354 232872
rect 215404 229094 215432 395830
rect 215496 232529 215524 504358
rect 215588 235249 215616 504494
rect 215668 504280 215720 504286
rect 215668 504222 215720 504228
rect 215574 235240 215630 235249
rect 215574 235175 215630 235184
rect 215680 233073 215708 504222
rect 215666 233064 215722 233073
rect 215666 232999 215722 233008
rect 215772 232665 215800 504766
rect 215852 504348 215904 504354
rect 215852 504290 215904 504296
rect 215864 232801 215892 504290
rect 215956 399770 215984 700402
rect 218992 699718 219020 703520
rect 235184 700738 235212 703520
rect 235172 700732 235224 700738
rect 235172 700674 235224 700680
rect 267660 700670 267688 703520
rect 267648 700664 267700 700670
rect 267648 700606 267700 700612
rect 283852 700602 283880 703520
rect 283840 700596 283892 700602
rect 283840 700538 283892 700544
rect 300136 700534 300164 703520
rect 300124 700528 300176 700534
rect 300124 700470 300176 700476
rect 332520 700466 332548 703520
rect 332508 700460 332560 700466
rect 332508 700402 332560 700408
rect 348804 700398 348832 703520
rect 348792 700392 348844 700398
rect 348792 700334 348844 700340
rect 364996 699718 365024 703520
rect 397472 700602 397500 703520
rect 377404 700596 377456 700602
rect 377404 700538 377456 700544
rect 397460 700596 397512 700602
rect 397460 700538 397512 700544
rect 376024 700528 376076 700534
rect 376024 700470 376076 700476
rect 374644 700392 374696 700398
rect 374644 700334 374696 700340
rect 218980 699712 219032 699718
rect 218980 699654 219032 699660
rect 360844 699712 360896 699718
rect 360844 699654 360896 699660
rect 364984 699712 365036 699718
rect 364984 699654 365036 699660
rect 218888 505776 218940 505782
rect 218888 505718 218940 505724
rect 218704 505708 218756 505714
rect 218704 505650 218756 505656
rect 216312 505640 216364 505646
rect 216312 505582 216364 505588
rect 216128 505572 216180 505578
rect 216128 505514 216180 505520
rect 216036 503736 216088 503742
rect 216036 503678 216088 503684
rect 215944 399764 215996 399770
rect 215944 399706 215996 399712
rect 215850 232792 215906 232801
rect 215850 232727 215906 232736
rect 215758 232656 215814 232665
rect 215758 232591 215814 232600
rect 215482 232520 215538 232529
rect 215482 232455 215538 232464
rect 215404 229066 215984 229094
rect 215758 227488 215814 227497
rect 215758 227423 215814 227432
rect 215772 226658 215800 227423
rect 213104 226630 213486 226658
rect 214498 226630 214972 226658
rect 215418 226630 215800 226658
rect 215956 226658 215984 229066
rect 216048 226953 216076 503678
rect 216140 230081 216168 505514
rect 216220 504280 216272 504286
rect 216220 504222 216272 504228
rect 216126 230072 216182 230081
rect 216126 230007 216182 230016
rect 216232 228721 216260 504222
rect 216324 229809 216352 505582
rect 216496 505504 216548 505510
rect 216496 505446 216548 505452
rect 216404 504348 216456 504354
rect 216404 504290 216456 504296
rect 216310 229800 216366 229809
rect 216310 229735 216366 229744
rect 216416 228857 216444 504290
rect 216508 229945 216536 505446
rect 217784 505232 217836 505238
rect 217784 505174 217836 505180
rect 216588 504416 216640 504422
rect 216588 504358 216640 504364
rect 216494 229936 216550 229945
rect 216494 229871 216550 229880
rect 216402 228848 216458 228857
rect 216402 228783 216458 228792
rect 216218 228712 216274 228721
rect 216218 228647 216274 228656
rect 216600 227497 216628 504358
rect 217690 435976 217746 435985
rect 217690 435911 217746 435920
rect 217598 433800 217654 433809
rect 217598 433735 217654 433744
rect 217414 432848 217470 432857
rect 217414 432783 217470 432792
rect 216678 431080 216734 431089
rect 216678 431015 216734 431024
rect 216692 430642 216720 431015
rect 216680 430636 216732 430642
rect 216680 430578 216732 430584
rect 216678 429992 216734 430001
rect 216678 429927 216734 429936
rect 216692 429214 216720 429927
rect 216680 429208 216732 429214
rect 216680 429150 216732 429156
rect 217230 410000 217286 410009
rect 217230 409935 217286 409944
rect 216678 408232 216734 408241
rect 216678 408167 216734 408176
rect 216692 407930 216720 408167
rect 216770 408096 216826 408105
rect 216770 408031 216826 408040
rect 216680 407924 216732 407930
rect 216680 407866 216732 407872
rect 216784 407182 216812 408031
rect 216772 407176 216824 407182
rect 216772 407118 216824 407124
rect 217244 240174 217272 409935
rect 217428 399974 217456 432783
rect 217416 399968 217468 399974
rect 217416 399910 217468 399916
rect 217612 399906 217640 433735
rect 217600 399900 217652 399906
rect 217600 399842 217652 399848
rect 217704 399838 217732 435911
rect 217692 399832 217744 399838
rect 217692 399774 217744 399780
rect 217796 398138 217824 505174
rect 218612 505164 218664 505170
rect 218612 505106 218664 505112
rect 218428 504824 218480 504830
rect 218428 504766 218480 504772
rect 218336 504688 218388 504694
rect 218336 504630 218388 504636
rect 218244 503736 218296 503742
rect 218244 503678 218296 503684
rect 218152 503532 218204 503538
rect 218152 503474 218204 503480
rect 218060 503464 218112 503470
rect 218060 503406 218112 503412
rect 217966 436928 218022 436937
rect 217966 436863 218022 436872
rect 217874 428224 217930 428233
rect 217874 428159 217930 428168
rect 217888 399770 217916 428159
rect 217876 399764 217928 399770
rect 217876 399706 217928 399712
rect 217784 398132 217836 398138
rect 217784 398074 217836 398080
rect 217232 240168 217284 240174
rect 217232 240110 217284 240116
rect 217322 230888 217378 230897
rect 217322 230823 217378 230832
rect 216586 227488 216642 227497
rect 216586 227423 216642 227432
rect 216034 226944 216090 226953
rect 216034 226879 216090 226888
rect 215956 226630 216338 226658
rect 217336 226644 217364 230823
rect 217980 228313 218008 436863
rect 218072 398206 218100 503406
rect 218164 398750 218192 503474
rect 218152 398744 218204 398750
rect 218152 398686 218204 398692
rect 218256 398274 218284 503678
rect 218348 398342 218376 504630
rect 218336 398336 218388 398342
rect 218336 398278 218388 398284
rect 218244 398268 218296 398274
rect 218244 398210 218296 398216
rect 218060 398200 218112 398206
rect 218060 398142 218112 398148
rect 218440 398002 218468 504766
rect 218520 504552 218572 504558
rect 218520 504494 218572 504500
rect 218532 398818 218560 504494
rect 218520 398812 218572 398818
rect 218520 398754 218572 398760
rect 218428 397996 218480 398002
rect 218428 397938 218480 397944
rect 218624 397866 218652 505106
rect 218612 397860 218664 397866
rect 218612 397802 218664 397808
rect 218152 244248 218204 244254
rect 218152 244190 218204 244196
rect 217966 228304 218022 228313
rect 217966 228239 218022 228248
rect 218164 226658 218192 244190
rect 218716 227361 218744 505650
rect 218796 505436 218848 505442
rect 218796 505378 218848 505384
rect 218808 230217 218836 505378
rect 218794 230208 218850 230217
rect 218794 230143 218850 230152
rect 218900 227497 218928 505718
rect 219808 505504 219860 505510
rect 219808 505446 219860 505452
rect 260840 505504 260892 505510
rect 260840 505446 260892 505452
rect 219164 505436 219216 505442
rect 219164 505378 219216 505384
rect 219072 505300 219124 505306
rect 219072 505242 219124 505248
rect 218980 504960 219032 504966
rect 218980 504902 219032 504908
rect 218992 233209 219020 504902
rect 218978 233200 219034 233209
rect 218978 233135 219034 233144
rect 218886 227488 218942 227497
rect 218886 227423 218942 227432
rect 218702 227352 218758 227361
rect 218702 227287 218758 227296
rect 219084 227089 219112 505242
rect 219176 398614 219204 505378
rect 219256 505368 219308 505374
rect 219256 505310 219308 505316
rect 219348 505368 219400 505374
rect 219348 505310 219400 505316
rect 219164 398608 219216 398614
rect 219164 398550 219216 398556
rect 219268 227225 219296 505310
rect 219360 398546 219388 505310
rect 219716 505300 219768 505306
rect 219716 505242 219768 505248
rect 219624 504960 219676 504966
rect 219624 504902 219676 504908
rect 219440 504892 219492 504898
rect 219440 504834 219492 504840
rect 219452 403102 219480 504834
rect 219532 504756 219584 504762
rect 219532 504698 219584 504704
rect 219440 403096 219492 403102
rect 219440 403038 219492 403044
rect 219544 402966 219572 504698
rect 219636 412690 219664 504902
rect 219624 412684 219676 412690
rect 219624 412626 219676 412632
rect 219624 412548 219676 412554
rect 219624 412490 219676 412496
rect 219636 405890 219664 412490
rect 219624 405884 219676 405890
rect 219624 405826 219676 405832
rect 219728 405770 219756 505242
rect 219820 486470 219848 505446
rect 219992 505096 220044 505102
rect 219992 505038 220044 505044
rect 219900 504620 219952 504626
rect 219900 504562 219952 504568
rect 219912 495434 219940 504562
rect 220004 499574 220032 505038
rect 252558 504112 252614 504121
rect 252558 504047 252614 504056
rect 220728 503668 220780 503674
rect 220728 503610 220780 503616
rect 245844 503668 245896 503674
rect 245844 503610 245896 503616
rect 220004 499546 220124 499574
rect 219912 495406 220032 495434
rect 220004 492674 220032 495406
rect 219912 492646 220032 492674
rect 219912 491294 219940 492646
rect 220096 491294 220124 499546
rect 220740 495434 220768 503610
rect 245856 503577 245884 503610
rect 245842 503568 245898 503577
rect 245842 503503 245898 503512
rect 252572 502334 252600 504047
rect 260852 503577 260880 505446
rect 288440 505436 288492 505442
rect 288440 505378 288492 505384
rect 273260 504960 273312 504966
rect 273260 504902 273312 504908
rect 270500 504144 270552 504150
rect 270500 504086 270552 504092
rect 265716 504076 265768 504082
rect 265716 504018 265768 504024
rect 263600 503600 263652 503606
rect 260838 503568 260894 503577
rect 265728 503577 265756 504018
rect 267740 504008 267792 504014
rect 267740 503950 267792 503956
rect 267752 503577 267780 503950
rect 270512 503577 270540 504086
rect 273272 503577 273300 504902
rect 277308 504892 277360 504898
rect 277308 504834 277360 504840
rect 277320 503577 277348 504834
rect 277400 504824 277452 504830
rect 277400 504766 277452 504772
rect 277412 503713 277440 504766
rect 280160 504756 280212 504762
rect 280160 504698 280212 504704
rect 277398 503704 277454 503713
rect 277398 503639 277454 503648
rect 280172 503577 280200 504698
rect 282920 504688 282972 504694
rect 282920 504630 282972 504636
rect 263600 503542 263652 503548
rect 265714 503568 265770 503577
rect 260838 503503 260894 503512
rect 252572 502306 253520 502334
rect 220188 495406 220768 495434
rect 220188 492674 220216 495406
rect 253492 494054 253520 502306
rect 263612 499574 263640 503542
rect 265714 503503 265770 503512
rect 267738 503568 267794 503577
rect 267738 503503 267794 503512
rect 270498 503568 270554 503577
rect 270498 503503 270554 503512
rect 273258 503568 273314 503577
rect 273258 503503 273314 503512
rect 277306 503568 277362 503577
rect 277306 503503 277362 503512
rect 280158 503568 280214 503577
rect 280158 503503 280214 503512
rect 282932 499574 282960 504630
rect 288452 503713 288480 505378
rect 298100 505368 298152 505374
rect 298100 505310 298152 505316
rect 295340 504552 295392 504558
rect 295340 504494 295392 504500
rect 292580 503736 292632 503742
rect 288438 503704 288494 503713
rect 292580 503678 292632 503684
rect 288438 503639 288494 503648
rect 292592 503577 292620 503678
rect 295352 503577 295380 504494
rect 285678 503568 285734 503577
rect 285678 503503 285680 503512
rect 285732 503503 285734 503512
rect 286874 503568 286930 503577
rect 286874 503503 286930 503512
rect 292578 503568 292634 503577
rect 292578 503503 292634 503512
rect 295338 503568 295394 503577
rect 295338 503503 295394 503512
rect 285680 503474 285732 503480
rect 286888 503470 286916 503503
rect 286876 503464 286928 503470
rect 286876 503406 286928 503412
rect 263612 499546 263732 499574
rect 282932 499546 284432 499574
rect 253308 494026 253520 494054
rect 220188 492646 220308 492674
rect 219912 491266 220032 491294
rect 220096 491266 220216 491294
rect 220004 486554 220032 491266
rect 220004 486526 220124 486554
rect 219808 486464 219860 486470
rect 219808 486406 219860 486412
rect 219806 486024 219862 486033
rect 220096 486010 220124 486526
rect 219862 485982 220124 486010
rect 219806 485959 219862 485968
rect 220188 483834 220216 491266
rect 219820 483806 220216 483834
rect 219820 483410 219848 483806
rect 220280 483698 220308 492646
rect 253308 487665 253336 494026
rect 263704 487665 263732 499546
rect 284404 487665 284432 499546
rect 298112 492697 298140 505310
rect 300860 505300 300912 505306
rect 300860 505242 300912 505248
rect 300872 492697 300900 505242
rect 316040 505232 316092 505238
rect 316040 505174 316092 505180
rect 307760 504484 307812 504490
rect 307760 504426 307812 504432
rect 302240 503940 302292 503946
rect 302240 503882 302292 503888
rect 302252 492697 302280 503882
rect 305000 503872 305052 503878
rect 305000 503814 305052 503820
rect 305012 492697 305040 503814
rect 307772 492697 307800 504426
rect 313280 504416 313332 504422
rect 313280 504358 313332 504364
rect 310520 503804 310572 503810
rect 310520 503746 310572 503752
rect 310532 492697 310560 503746
rect 313292 492697 313320 504358
rect 316052 492697 316080 505174
rect 325700 505164 325752 505170
rect 325700 505106 325752 505112
rect 317420 505028 317472 505034
rect 317420 504970 317472 504976
rect 317432 492697 317460 504970
rect 320180 504348 320232 504354
rect 320180 504290 320232 504296
rect 320192 492697 320220 504290
rect 322940 504280 322992 504286
rect 322940 504222 322992 504228
rect 322952 503577 322980 504222
rect 322938 503568 322994 503577
rect 322938 503503 322994 503512
rect 325712 498194 325740 505106
rect 339500 504212 339552 504218
rect 339500 504154 339552 504160
rect 339408 503532 339460 503538
rect 339408 503474 339460 503480
rect 325620 498166 325740 498194
rect 325620 495434 325648 498166
rect 325620 495406 326660 495434
rect 298098 492688 298154 492697
rect 298098 492623 298154 492632
rect 300858 492688 300914 492697
rect 300858 492623 300914 492632
rect 302238 492688 302294 492697
rect 302238 492623 302294 492632
rect 304998 492688 305054 492697
rect 304998 492623 305054 492632
rect 307758 492688 307814 492697
rect 307758 492623 307814 492632
rect 310518 492688 310574 492697
rect 310518 492623 310574 492632
rect 313278 492688 313334 492697
rect 313278 492623 313334 492632
rect 316038 492688 316094 492697
rect 316038 492623 316094 492632
rect 317418 492688 317474 492697
rect 317418 492623 317474 492632
rect 320178 492688 320234 492697
rect 320178 492623 320234 492632
rect 298112 492563 298140 492623
rect 300872 492563 300900 492623
rect 302252 492563 302280 492623
rect 305012 492563 305040 492623
rect 307772 492563 307800 492623
rect 310532 492563 310560 492623
rect 313292 492563 313320 492623
rect 316052 492563 316080 492623
rect 317432 492563 317460 492623
rect 320192 492563 320220 492623
rect 326632 488345 326660 495406
rect 339420 492697 339448 503474
rect 339512 492697 339540 504154
rect 356520 503532 356572 503538
rect 356520 503474 356572 503480
rect 350540 503464 350592 503470
rect 350540 503406 350592 503412
rect 350552 499574 350580 503406
rect 356532 499574 356560 503474
rect 350552 499546 351868 499574
rect 356532 499546 356744 499574
rect 339406 492688 339462 492697
rect 339406 492623 339462 492632
rect 339498 492688 339554 492697
rect 339498 492623 339554 492632
rect 339420 492563 339448 492623
rect 339512 492563 339540 492623
rect 326618 488336 326674 488345
rect 326618 488271 326674 488280
rect 253294 487656 253350 487665
rect 253294 487591 253350 487600
rect 263690 487656 263746 487665
rect 263690 487591 263746 487600
rect 284390 487656 284446 487665
rect 284390 487591 284446 487600
rect 351840 485874 351868 499546
rect 356716 492674 356744 499546
rect 356716 492646 356928 492674
rect 351840 485846 356468 485874
rect 356440 485774 356468 485846
rect 356440 485746 356652 485774
rect 356624 485466 356652 485746
rect 356794 485480 356850 485489
rect 356624 485438 356794 485466
rect 356794 485415 356850 485424
rect 220096 483670 220308 483698
rect 220096 483562 220124 483670
rect 219912 483534 220124 483562
rect 219808 483404 219860 483410
rect 219808 483346 219860 483352
rect 219808 483268 219860 483274
rect 219912 483256 219940 483534
rect 219860 483228 219940 483256
rect 219808 483210 219860 483216
rect 356900 483014 356928 492646
rect 356716 482986 356928 483014
rect 219808 481432 219860 481438
rect 219860 481380 220032 481386
rect 219808 481374 220032 481380
rect 219820 481358 220032 481374
rect 219806 480992 219862 481001
rect 219806 480927 219862 480936
rect 219820 480842 219848 480927
rect 219820 480814 219940 480842
rect 219808 480752 219860 480758
rect 219808 480694 219860 480700
rect 219820 470694 219848 480694
rect 219808 470688 219860 470694
rect 219808 470630 219860 470636
rect 219808 470552 219860 470558
rect 219808 470494 219860 470500
rect 219820 451382 219848 470494
rect 219808 451376 219860 451382
rect 219808 451318 219860 451324
rect 219808 451240 219860 451246
rect 219808 451182 219860 451188
rect 219820 432070 219848 451182
rect 219808 432064 219860 432070
rect 219808 432006 219860 432012
rect 219808 431928 219860 431934
rect 219808 431870 219860 431876
rect 219820 422414 219848 431870
rect 219808 422408 219860 422414
rect 219808 422350 219860 422356
rect 219808 422272 219860 422278
rect 219808 422214 219860 422220
rect 219820 412758 219848 422214
rect 219808 412752 219860 412758
rect 219808 412694 219860 412700
rect 219808 412646 219860 412652
rect 219808 412588 219860 412594
rect 219636 405742 219756 405770
rect 219532 402960 219584 402966
rect 219532 402902 219584 402908
rect 219440 402892 219492 402898
rect 219440 402834 219492 402840
rect 219348 398540 219400 398546
rect 219348 398482 219400 398488
rect 219452 398070 219480 402834
rect 219532 402824 219584 402830
rect 219532 402766 219584 402772
rect 219544 398818 219572 402766
rect 219532 398812 219584 398818
rect 219532 398754 219584 398760
rect 219636 398410 219664 405742
rect 219716 405680 219768 405686
rect 219716 405622 219768 405628
rect 219728 398478 219756 405622
rect 219820 398682 219848 412588
rect 219808 398676 219860 398682
rect 219808 398618 219860 398624
rect 219716 398472 219768 398478
rect 219716 398414 219768 398420
rect 219624 398404 219676 398410
rect 219624 398346 219676 398352
rect 219440 398064 219492 398070
rect 219440 398006 219492 398012
rect 219348 242480 219400 242486
rect 219348 242422 219400 242428
rect 219254 227216 219310 227225
rect 219254 227151 219310 227160
rect 219070 227080 219126 227089
rect 219070 227015 219126 227024
rect 219360 226658 219388 242422
rect 219912 230489 219940 480814
rect 219898 230480 219954 230489
rect 219898 230415 219954 230424
rect 220004 226817 220032 481358
rect 356716 470594 356744 482986
rect 357438 479224 357494 479233
rect 357438 479159 357494 479168
rect 356532 470566 356744 470594
rect 226340 399900 226392 399906
rect 226340 399842 226392 399848
rect 224500 398812 224552 398818
rect 224500 398754 224552 398760
rect 222108 396500 222160 396506
rect 222108 396442 222160 396448
rect 220084 396432 220136 396438
rect 220084 396374 220136 396380
rect 220096 230897 220124 396374
rect 220082 230888 220138 230897
rect 220082 230823 220138 230832
rect 222120 229094 222148 396442
rect 222844 396364 222896 396370
rect 222844 396306 222896 396312
rect 222200 395956 222252 395962
rect 222200 395898 222252 395904
rect 222212 248414 222240 395898
rect 222212 248386 222608 248414
rect 221568 229066 222148 229094
rect 220174 228848 220230 228857
rect 220174 228783 220230 228792
rect 219990 226808 220046 226817
rect 219990 226743 220046 226752
rect 218164 226630 218270 226658
rect 219190 226630 219388 226658
rect 220188 226644 220216 228783
rect 221568 226658 221596 229066
rect 222014 228712 222070 228721
rect 222014 228647 222070 228656
rect 221122 226630 221596 226658
rect 222028 226644 222056 228647
rect 222580 226658 222608 248386
rect 222856 227905 222884 396306
rect 223672 249348 223724 249354
rect 223672 249290 223724 249296
rect 222842 227896 222898 227905
rect 222842 227831 222898 227840
rect 222580 226630 223054 226658
rect 181810 226607 181866 226616
rect 223684 226001 223712 249290
rect 224222 226672 224278 226681
rect 223974 226630 224222 226658
rect 224222 226607 224278 226616
rect 61750 225992 61806 226001
rect 61750 225927 61806 225936
rect 78862 225992 78918 226001
rect 78862 225927 78918 225936
rect 223670 225992 223726 226001
rect 223670 225927 223726 225936
rect 59726 72040 59782 72049
rect 59726 71975 59782 71984
rect 59174 61296 59230 61305
rect 59174 61231 59230 61240
rect 59820 60308 59872 60314
rect 59820 60250 59872 60256
rect 59832 60058 59860 60250
rect 221738 60208 221794 60217
rect 221582 60166 221738 60194
rect 221738 60143 221794 60152
rect 222934 60072 222990 60081
rect 59832 60044 60122 60058
rect 59832 60030 60136 60044
rect 58714 57896 58770 57905
rect 58348 57860 58400 57866
rect 58714 57831 58770 57840
rect 58348 57802 58400 57808
rect 57244 56704 57296 56710
rect 57244 56646 57296 56652
rect 56140 55956 56192 55962
rect 56140 55898 56192 55904
rect 55772 33108 55824 33114
rect 55772 33050 55824 33056
rect 55680 20664 55732 20670
rect 55680 20606 55732 20612
rect 57256 6914 57284 56646
rect 60108 55894 60136 60030
rect 60384 56370 60412 60044
rect 60372 56364 60424 56370
rect 60372 56306 60424 56312
rect 60660 56030 60688 60044
rect 60936 57254 60964 60044
rect 61028 60030 61226 60058
rect 60924 57248 60976 57254
rect 60924 57190 60976 57196
rect 60648 56024 60700 56030
rect 60648 55966 60700 55972
rect 60096 55888 60148 55894
rect 60096 55830 60148 55836
rect 59268 55548 59320 55554
rect 59268 55490 59320 55496
rect 54956 6886 55168 6914
rect 57164 6886 57284 6914
rect 54956 480 54984 6886
rect 56048 3188 56100 3194
rect 56048 3130 56100 3136
rect 56060 480 56088 3130
rect 57164 3058 57192 6886
rect 59280 3534 59308 55490
rect 60832 4004 60884 4010
rect 60832 3946 60884 3952
rect 58440 3528 58492 3534
rect 58440 3470 58492 3476
rect 59268 3528 59320 3534
rect 59268 3470 59320 3476
rect 57152 3052 57204 3058
rect 57152 2994 57204 3000
rect 57244 3052 57296 3058
rect 57244 2994 57296 3000
rect 57256 480 57284 2994
rect 58452 480 58480 3470
rect 59636 2984 59688 2990
rect 59636 2926 59688 2932
rect 59648 480 59676 2926
rect 60844 480 60872 3946
rect 61028 3398 61056 60030
rect 61580 57390 61608 60044
rect 61568 57384 61620 57390
rect 61568 57326 61620 57332
rect 61856 56098 61884 60044
rect 61844 56092 61896 56098
rect 61844 56034 61896 56040
rect 62028 4820 62080 4826
rect 62028 4762 62080 4768
rect 61016 3392 61068 3398
rect 61016 3334 61068 3340
rect 62040 480 62068 4762
rect 62132 3602 62160 60044
rect 62408 57322 62436 60044
rect 62500 60030 62790 60058
rect 62396 57316 62448 57322
rect 62396 57258 62448 57264
rect 62500 3670 62528 60030
rect 62764 57384 62816 57390
rect 62764 57326 62816 57332
rect 62488 3664 62540 3670
rect 62488 3606 62540 3612
rect 62120 3596 62172 3602
rect 62120 3538 62172 3544
rect 62776 3126 62804 57326
rect 62948 56772 63000 56778
rect 62948 56714 63000 56720
rect 62856 56636 62908 56642
rect 62856 56578 62908 56584
rect 62868 3262 62896 56578
rect 62960 3738 62988 56714
rect 63052 56574 63080 60044
rect 63328 57526 63356 60044
rect 63512 60030 63618 60058
rect 63696 60030 63986 60058
rect 64064 60030 64262 60058
rect 63316 57520 63368 57526
rect 63316 57462 63368 57468
rect 63512 57458 63540 60030
rect 63696 57712 63724 60030
rect 63604 57684 63724 57712
rect 63604 57594 63632 57684
rect 63592 57588 63644 57594
rect 63592 57530 63644 57536
rect 63500 57452 63552 57458
rect 63500 57394 63552 57400
rect 63684 57316 63736 57322
rect 63684 57258 63736 57264
rect 63040 56568 63092 56574
rect 63040 56510 63092 56516
rect 63696 3942 63724 57258
rect 64064 56166 64092 60030
rect 64524 58002 64552 60044
rect 64616 60030 64814 60058
rect 65076 60030 65182 60058
rect 64512 57996 64564 58002
rect 64512 57938 64564 57944
rect 64144 57520 64196 57526
rect 64144 57462 64196 57468
rect 64052 56160 64104 56166
rect 64052 56102 64104 56108
rect 64156 4146 64184 57462
rect 64420 57452 64472 57458
rect 64420 57394 64472 57400
rect 64236 57248 64288 57254
rect 64236 57190 64288 57196
rect 64144 4140 64196 4146
rect 64144 4082 64196 4088
rect 64248 4026 64276 57190
rect 64328 56704 64380 56710
rect 64328 56646 64380 56652
rect 64156 3998 64276 4026
rect 64340 4010 64368 56646
rect 64328 4004 64380 4010
rect 63684 3936 63736 3942
rect 63684 3878 63736 3884
rect 63776 3936 63828 3942
rect 63776 3878 63828 3884
rect 62948 3732 63000 3738
rect 62948 3674 63000 3680
rect 63224 3528 63276 3534
rect 63224 3470 63276 3476
rect 62856 3256 62908 3262
rect 62856 3198 62908 3204
rect 62764 3120 62816 3126
rect 62764 3062 62816 3068
rect 63236 480 63264 3470
rect 63788 2922 63816 3878
rect 64156 3602 64184 3998
rect 64328 3946 64380 3952
rect 64328 3868 64380 3874
rect 64328 3810 64380 3816
rect 64144 3596 64196 3602
rect 64144 3538 64196 3544
rect 63776 2916 63828 2922
rect 63776 2858 63828 2864
rect 64340 480 64368 3810
rect 64432 3330 64460 57394
rect 64616 57322 64644 60030
rect 64604 57316 64656 57322
rect 64604 57258 64656 57264
rect 64788 56772 64840 56778
rect 64788 56714 64840 56720
rect 64800 56658 64828 56714
rect 64616 56630 64828 56658
rect 64616 56574 64644 56630
rect 64604 56568 64656 56574
rect 64604 56510 64656 56516
rect 64420 3324 64472 3330
rect 64420 3266 64472 3272
rect 65076 2854 65104 60030
rect 65444 56234 65472 60044
rect 65616 57588 65668 57594
rect 65616 57530 65668 57536
rect 65524 57384 65576 57390
rect 65524 57326 65576 57332
rect 65432 56228 65484 56234
rect 65432 56170 65484 56176
rect 65536 4146 65564 57326
rect 65524 4140 65576 4146
rect 65524 4082 65576 4088
rect 65524 3392 65576 3398
rect 65524 3334 65576 3340
rect 65064 2848 65116 2854
rect 65064 2790 65116 2796
rect 65536 480 65564 3334
rect 65628 3058 65656 57530
rect 65720 56642 65748 60044
rect 65996 57730 66024 60044
rect 66364 57798 66392 60044
rect 66352 57792 66404 57798
rect 66352 57734 66404 57740
rect 66640 57730 66668 60044
rect 66916 57934 66944 60044
rect 67008 60030 67206 60058
rect 66904 57928 66956 57934
rect 66904 57870 66956 57876
rect 65984 57724 66036 57730
rect 65984 57666 66036 57672
rect 66076 57724 66128 57730
rect 66076 57666 66128 57672
rect 66628 57724 66680 57730
rect 66628 57666 66680 57672
rect 65708 56636 65760 56642
rect 65708 56578 65760 56584
rect 65984 56636 66036 56642
rect 65984 56578 66036 56584
rect 65996 56370 66024 56578
rect 65984 56364 66036 56370
rect 65984 56306 66036 56312
rect 66088 56302 66116 57666
rect 67008 57610 67036 60030
rect 67088 57792 67140 57798
rect 67088 57734 67140 57740
rect 66456 57582 67036 57610
rect 66076 56296 66128 56302
rect 66076 56238 66128 56244
rect 66456 3466 66484 57582
rect 66904 57520 66956 57526
rect 66904 57462 66956 57468
rect 66916 3806 66944 57462
rect 66996 57044 67048 57050
rect 66996 56986 67048 56992
rect 67008 3874 67036 56986
rect 67100 4078 67128 57734
rect 67468 56642 67496 60044
rect 67548 57588 67600 57594
rect 67548 57530 67600 57536
rect 67456 56636 67508 56642
rect 67456 56578 67508 56584
rect 67088 4072 67140 4078
rect 67088 4014 67140 4020
rect 66996 3868 67048 3874
rect 66996 3810 67048 3816
rect 66904 3800 66956 3806
rect 66904 3742 66956 3748
rect 67560 3466 67588 57530
rect 67836 57458 67864 60044
rect 67824 57452 67876 57458
rect 67824 57394 67876 57400
rect 68112 57186 68140 60044
rect 68204 60030 68402 60058
rect 68100 57180 68152 57186
rect 68100 57122 68152 57128
rect 68204 56506 68232 60030
rect 68284 57928 68336 57934
rect 68284 57870 68336 57876
rect 68192 56500 68244 56506
rect 68192 56442 68244 56448
rect 66444 3460 66496 3466
rect 66444 3402 66496 3408
rect 66720 3460 66772 3466
rect 66720 3402 66772 3408
rect 67548 3460 67600 3466
rect 67548 3402 67600 3408
rect 67916 3460 67968 3466
rect 67916 3402 67968 3408
rect 65616 3052 65668 3058
rect 65616 2994 65668 3000
rect 66732 480 66760 3402
rect 67928 480 67956 3402
rect 68296 3194 68324 57870
rect 68664 57118 68692 60044
rect 69032 57526 69060 60044
rect 69216 60030 69322 60058
rect 69020 57520 69072 57526
rect 69020 57462 69072 57468
rect 68652 57112 68704 57118
rect 68652 57054 68704 57060
rect 68928 57112 68980 57118
rect 68928 57054 68980 57060
rect 68376 56772 68428 56778
rect 68376 56714 68428 56720
rect 68284 3188 68336 3194
rect 68284 3130 68336 3136
rect 68388 2990 68416 56714
rect 68940 3466 68968 57054
rect 69216 54534 69244 60030
rect 69584 57662 69612 60044
rect 69572 57656 69624 57662
rect 69572 57598 69624 57604
rect 69860 56982 69888 60044
rect 69952 60030 70242 60058
rect 69848 56976 69900 56982
rect 69848 56918 69900 56924
rect 69952 55826 69980 60030
rect 70308 57724 70360 57730
rect 70308 57666 70360 57672
rect 70216 57656 70268 57662
rect 70216 57598 70268 57604
rect 69940 55820 69992 55826
rect 69940 55762 69992 55768
rect 69204 54528 69256 54534
rect 69204 54470 69256 54476
rect 70228 3466 70256 57598
rect 68928 3460 68980 3466
rect 68928 3402 68980 3408
rect 69112 3460 69164 3466
rect 69112 3402 69164 3408
rect 70216 3460 70268 3466
rect 70216 3402 70268 3408
rect 68376 2984 68428 2990
rect 68376 2926 68428 2932
rect 69124 480 69152 3402
rect 70320 480 70348 57666
rect 70504 57254 70532 60044
rect 70780 57798 70808 60044
rect 70768 57792 70820 57798
rect 70768 57734 70820 57740
rect 71056 57458 71084 60044
rect 71148 60030 71438 60058
rect 71516 60030 71714 60058
rect 71044 57452 71096 57458
rect 71044 57394 71096 57400
rect 70492 57248 70544 57254
rect 70492 57190 70544 57196
rect 70400 56840 70452 56846
rect 70400 56782 70452 56788
rect 70412 55554 70440 56782
rect 71148 56760 71176 60030
rect 70964 56732 71176 56760
rect 70964 56642 70992 56732
rect 71516 56710 71544 60030
rect 71688 57248 71740 57254
rect 71688 57190 71740 57196
rect 71504 56704 71556 56710
rect 71504 56646 71556 56652
rect 70952 56636 71004 56642
rect 70952 56578 71004 56584
rect 71044 56636 71096 56642
rect 71044 56578 71096 56584
rect 70400 55548 70452 55554
rect 70400 55490 70452 55496
rect 71056 4826 71084 56578
rect 71700 6914 71728 57190
rect 71976 55758 72004 60044
rect 72252 57526 72280 60044
rect 72240 57520 72292 57526
rect 72240 57462 72292 57468
rect 72620 57186 72648 60044
rect 72608 57180 72660 57186
rect 72608 57122 72660 57128
rect 71964 55752 72016 55758
rect 71964 55694 72016 55700
rect 72896 55690 72924 60044
rect 73068 57452 73120 57458
rect 73068 57394 73120 57400
rect 72884 55684 72936 55690
rect 72884 55626 72936 55632
rect 71516 6886 71728 6914
rect 71044 4820 71096 4826
rect 71044 4762 71096 4768
rect 71516 480 71544 6886
rect 73080 3466 73108 57394
rect 73172 57322 73200 60044
rect 73160 57316 73212 57322
rect 73160 57258 73212 57264
rect 73448 56982 73476 60044
rect 73436 56976 73488 56982
rect 73436 56918 73488 56924
rect 73816 55622 73844 60044
rect 74092 57934 74120 60044
rect 74080 57928 74132 57934
rect 74080 57870 74132 57876
rect 74368 57798 74396 60044
rect 74552 60030 74658 60058
rect 74356 57792 74408 57798
rect 74356 57734 74408 57740
rect 74552 56846 74580 60030
rect 74724 57588 74776 57594
rect 74724 57530 74776 57536
rect 74540 56840 74592 56846
rect 74540 56782 74592 56788
rect 73804 55616 73856 55622
rect 73804 55558 73856 55564
rect 74736 3534 74764 57530
rect 74920 56778 74948 60044
rect 75012 60030 75302 60058
rect 75012 57390 75040 60030
rect 75184 57452 75236 57458
rect 75184 57394 75236 57400
rect 75000 57384 75052 57390
rect 75000 57326 75052 57332
rect 74908 56772 74960 56778
rect 74908 56714 74960 56720
rect 74724 3528 74776 3534
rect 74724 3470 74776 3476
rect 75000 3528 75052 3534
rect 75000 3470 75052 3476
rect 72608 3460 72660 3466
rect 72608 3402 72660 3408
rect 73068 3460 73120 3466
rect 73068 3402 73120 3408
rect 73804 3460 73856 3466
rect 73804 3402 73856 3408
rect 72620 480 72648 3402
rect 73816 480 73844 3402
rect 75012 480 75040 3470
rect 75196 3466 75224 57394
rect 75564 56642 75592 60044
rect 75656 60030 75854 60058
rect 75656 57594 75684 60030
rect 75644 57588 75696 57594
rect 75644 57530 75696 57536
rect 75828 57180 75880 57186
rect 75828 57122 75880 57128
rect 75552 56636 75604 56642
rect 75552 56578 75604 56584
rect 75840 3534 75868 57122
rect 76116 57050 76144 60044
rect 76208 60030 76498 60058
rect 76104 57044 76156 57050
rect 76104 56986 76156 56992
rect 76208 6914 76236 60030
rect 76760 57526 76788 60044
rect 76748 57520 76800 57526
rect 76748 57462 76800 57468
rect 77036 57118 77064 60044
rect 77312 57662 77340 60044
rect 77680 57730 77708 60044
rect 77668 57724 77720 57730
rect 77668 57666 77720 57672
rect 77300 57656 77352 57662
rect 77300 57598 77352 57604
rect 77208 57588 77260 57594
rect 77208 57530 77260 57536
rect 77024 57112 77076 57118
rect 77024 57054 77076 57060
rect 76116 6886 76236 6914
rect 75828 3528 75880 3534
rect 75828 3470 75880 3476
rect 75184 3460 75236 3466
rect 75184 3402 75236 3408
rect 76116 3398 76144 6886
rect 77220 3534 77248 57530
rect 77956 57254 77984 60044
rect 78232 57390 78260 60044
rect 78508 57458 78536 60044
rect 78772 57656 78824 57662
rect 78772 57598 78824 57604
rect 78496 57452 78548 57458
rect 78496 57394 78548 57400
rect 78220 57384 78272 57390
rect 78220 57326 78272 57332
rect 77944 57248 77996 57254
rect 77944 57190 77996 57196
rect 78784 6914 78812 57598
rect 78876 57186 78904 60044
rect 79152 57594 79180 60044
rect 79244 60030 79442 60058
rect 79520 60030 79718 60058
rect 80086 60030 80284 60058
rect 79140 57588 79192 57594
rect 79140 57530 79192 57536
rect 78864 57180 78916 57186
rect 78864 57122 78916 57128
rect 79244 45554 79272 60030
rect 79520 57662 79548 60030
rect 79508 57656 79560 57662
rect 79508 57598 79560 57604
rect 80256 57118 80284 60030
rect 80244 57112 80296 57118
rect 80244 57054 80296 57060
rect 80348 55706 80376 60044
rect 80428 57112 80480 57118
rect 80428 57054 80480 57060
rect 80256 55678 80376 55706
rect 80256 48314 80284 55678
rect 80256 48286 80376 48314
rect 78692 6886 78812 6914
rect 78968 45526 79272 45554
rect 76196 3528 76248 3534
rect 76196 3470 76248 3476
rect 77208 3528 77260 3534
rect 78692 3482 78720 6886
rect 77208 3470 77260 3476
rect 76104 3392 76156 3398
rect 76104 3334 76156 3340
rect 76208 480 76236 3470
rect 77392 3460 77444 3466
rect 77392 3402 77444 3408
rect 78600 3454 78720 3482
rect 78968 3466 78996 45526
rect 80348 3534 80376 48286
rect 80336 3528 80388 3534
rect 80336 3470 80388 3476
rect 80440 3466 80468 57054
rect 80624 56642 80652 60044
rect 80900 56846 80928 60044
rect 81190 60030 81388 60058
rect 80888 56840 80940 56846
rect 80888 56782 80940 56788
rect 80612 56636 80664 56642
rect 80612 56578 80664 56584
rect 81256 56636 81308 56642
rect 81256 56578 81308 56584
rect 81268 3534 81296 56578
rect 81360 3602 81388 60030
rect 81544 56642 81572 60044
rect 81820 56710 81848 60044
rect 82096 56778 82124 60044
rect 82386 60030 82676 60058
rect 82084 56772 82136 56778
rect 82084 56714 82136 56720
rect 81808 56704 81860 56710
rect 81808 56646 81860 56652
rect 81532 56636 81584 56642
rect 81532 56578 81584 56584
rect 82544 56636 82596 56642
rect 82544 56578 82596 56584
rect 82556 3874 82584 56578
rect 82544 3868 82596 3874
rect 82544 3810 82596 3816
rect 81348 3596 81400 3602
rect 81348 3538 81400 3544
rect 80888 3528 80940 3534
rect 80888 3470 80940 3476
rect 81256 3528 81308 3534
rect 81256 3470 81308 3476
rect 82084 3528 82136 3534
rect 82084 3470 82136 3476
rect 78956 3460 79008 3466
rect 77404 480 77432 3402
rect 78600 480 78628 3454
rect 78956 3402 79008 3408
rect 79692 3460 79744 3466
rect 79692 3402 79744 3408
rect 80428 3460 80480 3466
rect 80428 3402 80480 3408
rect 79704 480 79732 3402
rect 80900 480 80928 3470
rect 82096 480 82124 3470
rect 82648 3466 82676 60030
rect 82740 56982 82768 60044
rect 82728 56976 82780 56982
rect 82728 56918 82780 56924
rect 83016 56710 83044 60044
rect 83188 56840 83240 56846
rect 83188 56782 83240 56788
rect 82728 56704 82780 56710
rect 82728 56646 82780 56652
rect 83004 56704 83056 56710
rect 83004 56646 83056 56652
rect 82636 3460 82688 3466
rect 82636 3402 82688 3408
rect 82740 2922 82768 56646
rect 83200 16574 83228 56782
rect 83292 56642 83320 60044
rect 83568 57118 83596 60044
rect 83950 60030 84148 60058
rect 83556 57112 83608 57118
rect 83556 57054 83608 57060
rect 83464 56772 83516 56778
rect 83464 56714 83516 56720
rect 83280 56636 83332 56642
rect 83280 56578 83332 56584
rect 83200 16546 83320 16574
rect 82728 2916 82780 2922
rect 82728 2858 82780 2864
rect 83292 480 83320 16546
rect 83476 3602 83504 56714
rect 84016 56704 84068 56710
rect 84016 56646 84068 56652
rect 83924 56636 83976 56642
rect 83924 56578 83976 56584
rect 83464 3596 83516 3602
rect 83464 3538 83516 3544
rect 83936 2854 83964 56578
rect 84028 3670 84056 56646
rect 84016 3664 84068 3670
rect 84016 3606 84068 3612
rect 84120 3058 84148 60030
rect 84212 56778 84240 60044
rect 84488 56914 84516 60044
rect 84476 56908 84528 56914
rect 84476 56850 84528 56856
rect 84764 56846 84792 60044
rect 85146 60030 85344 60058
rect 84752 56840 84804 56846
rect 84752 56782 84804 56788
rect 84200 56772 84252 56778
rect 84200 56714 84252 56720
rect 85316 51074 85344 60030
rect 85408 57186 85436 60044
rect 85396 57180 85448 57186
rect 85396 57122 85448 57128
rect 85684 56642 85712 60044
rect 85960 56710 85988 60044
rect 86342 60030 86540 60058
rect 86618 60030 86724 60058
rect 86224 56772 86276 56778
rect 86224 56714 86276 56720
rect 85948 56704 86000 56710
rect 85948 56646 86000 56652
rect 85672 56636 85724 56642
rect 85672 56578 85724 56584
rect 85316 51046 85528 51074
rect 85500 3534 85528 51046
rect 85672 3868 85724 3874
rect 85672 3810 85724 3816
rect 84476 3528 84528 3534
rect 84476 3470 84528 3476
rect 85488 3528 85540 3534
rect 85488 3470 85540 3476
rect 84108 3052 84160 3058
rect 84108 2994 84160 3000
rect 83924 2848 83976 2854
rect 83924 2790 83976 2796
rect 84488 480 84516 3470
rect 85684 480 85712 3810
rect 86236 2990 86264 56714
rect 86512 51074 86540 60030
rect 86512 51046 86632 51074
rect 86604 22778 86632 51046
rect 86592 22772 86644 22778
rect 86592 22714 86644 22720
rect 86696 3330 86724 60030
rect 86880 57322 86908 60044
rect 87156 57866 87184 60044
rect 87144 57860 87196 57866
rect 87144 57802 87196 57808
rect 86868 57316 86920 57322
rect 86868 57258 86920 57264
rect 86868 56704 86920 56710
rect 86868 56646 86920 56652
rect 86776 56636 86828 56642
rect 86776 56578 86828 56584
rect 86684 3324 86736 3330
rect 86684 3266 86736 3272
rect 86788 3262 86816 56578
rect 86776 3256 86828 3262
rect 86776 3198 86828 3204
rect 86880 3126 86908 56646
rect 87524 56642 87552 60044
rect 87800 56982 87828 60044
rect 88090 60030 88196 60058
rect 87696 56976 87748 56982
rect 87696 56918 87748 56924
rect 87788 56976 87840 56982
rect 87788 56918 87840 56924
rect 87604 56840 87656 56846
rect 87604 56782 87656 56788
rect 87512 56636 87564 56642
rect 87512 56578 87564 56584
rect 87616 3194 87644 56782
rect 87708 4214 87736 56918
rect 88168 10334 88196 60030
rect 88352 56710 88380 60044
rect 88628 57458 88656 60044
rect 88616 57452 88668 57458
rect 88616 57394 88668 57400
rect 88892 56908 88944 56914
rect 88892 56850 88944 56856
rect 88340 56704 88392 56710
rect 88340 56646 88392 56652
rect 88248 56636 88300 56642
rect 88248 56578 88300 56584
rect 88156 10328 88208 10334
rect 88156 10270 88208 10276
rect 87696 4208 87748 4214
rect 87696 4150 87748 4156
rect 87972 3596 88024 3602
rect 87972 3538 88024 3544
rect 87604 3188 87656 3194
rect 87604 3130 87656 3136
rect 86868 3120 86920 3126
rect 86868 3062 86920 3068
rect 86224 2984 86276 2990
rect 86224 2926 86276 2932
rect 86868 2916 86920 2922
rect 86868 2858 86920 2864
rect 86880 480 86908 2858
rect 87984 480 88012 3538
rect 88260 3398 88288 56578
rect 88904 51074 88932 56850
rect 88996 56642 89024 60044
rect 89286 60030 89392 60058
rect 89562 60030 89668 60058
rect 88984 56636 89036 56642
rect 88984 56578 89036 56584
rect 88904 51046 89024 51074
rect 88996 18630 89024 51046
rect 88984 18624 89036 18630
rect 88984 18566 89036 18572
rect 89364 3534 89392 60030
rect 89444 56704 89496 56710
rect 89444 56646 89496 56652
rect 89456 4146 89484 56646
rect 89536 56636 89588 56642
rect 89536 56578 89588 56584
rect 89444 4140 89496 4146
rect 89444 4082 89496 4088
rect 89548 4078 89576 56578
rect 89536 4072 89588 4078
rect 89536 4014 89588 4020
rect 89640 3942 89668 60030
rect 89824 57322 89852 60044
rect 90192 57526 90220 60044
rect 90482 60030 90680 60058
rect 90758 60030 90956 60058
rect 90548 57724 90600 57730
rect 90548 57666 90600 57672
rect 90180 57520 90232 57526
rect 90180 57462 90232 57468
rect 89812 57316 89864 57322
rect 89812 57258 89864 57264
rect 90560 55214 90588 57666
rect 90652 57610 90680 60030
rect 90928 57610 90956 60030
rect 91020 57730 91048 60044
rect 91008 57724 91060 57730
rect 91008 57666 91060 57672
rect 90652 57582 90864 57610
rect 90928 57582 91048 57610
rect 90732 57316 90784 57322
rect 90732 57258 90784 57264
rect 90560 55186 90680 55214
rect 90364 4208 90416 4214
rect 90364 4150 90416 4156
rect 89628 3936 89680 3942
rect 89628 3878 89680 3884
rect 89352 3528 89404 3534
rect 89352 3470 89404 3476
rect 89168 3460 89220 3466
rect 89168 3402 89220 3408
rect 88248 3392 88300 3398
rect 88248 3334 88300 3340
rect 89180 480 89208 3402
rect 90376 480 90404 4150
rect 90652 3602 90680 55186
rect 90744 3874 90772 57258
rect 90732 3868 90784 3874
rect 90732 3810 90784 3816
rect 90836 3806 90864 57582
rect 90916 57520 90968 57526
rect 90916 57462 90968 57468
rect 90928 4010 90956 57462
rect 90916 4004 90968 4010
rect 90916 3946 90968 3952
rect 90824 3800 90876 3806
rect 90824 3742 90876 3748
rect 91020 3738 91048 57582
rect 91388 57118 91416 60044
rect 91664 57730 91692 60044
rect 91954 60030 92152 60058
rect 91652 57724 91704 57730
rect 91652 57666 91704 57672
rect 91376 57112 91428 57118
rect 91376 57054 91428 57060
rect 92124 55214 92152 60030
rect 92216 57186 92244 60044
rect 92584 57594 92612 60044
rect 92860 57662 92888 60044
rect 92848 57656 92900 57662
rect 92848 57598 92900 57604
rect 92572 57588 92624 57594
rect 92572 57530 92624 57536
rect 92204 57180 92256 57186
rect 92204 57122 92256 57128
rect 92388 57112 92440 57118
rect 92388 57054 92440 57060
rect 92124 55186 92336 55214
rect 92308 4350 92336 55186
rect 92296 4344 92348 4350
rect 92296 4286 92348 4292
rect 91008 3732 91060 3738
rect 91008 3674 91060 3680
rect 92400 3670 92428 57054
rect 93136 56030 93164 60044
rect 93124 56024 93176 56030
rect 93124 55966 93176 55972
rect 93412 4690 93440 60044
rect 93504 60030 93794 60058
rect 93504 6186 93532 60030
rect 93584 57656 93636 57662
rect 93584 57598 93636 57604
rect 93596 6254 93624 57598
rect 94056 57594 94084 60044
rect 94332 57730 94360 60044
rect 94320 57724 94372 57730
rect 94320 57666 94372 57672
rect 93676 57588 93728 57594
rect 93676 57530 93728 57536
rect 94044 57588 94096 57594
rect 94044 57530 94096 57536
rect 93584 6248 93636 6254
rect 93584 6190 93636 6196
rect 93492 6180 93544 6186
rect 93492 6122 93544 6128
rect 93400 4684 93452 4690
rect 93400 4626 93452 4632
rect 93688 4282 93716 57530
rect 94228 57248 94280 57254
rect 94228 57190 94280 57196
rect 94240 6914 94268 57190
rect 94608 57050 94636 60044
rect 94898 60030 95004 60058
rect 94872 57588 94924 57594
rect 94872 57530 94924 57536
rect 94596 57044 94648 57050
rect 94596 56986 94648 56992
rect 94884 17270 94912 57530
rect 94872 17264 94924 17270
rect 94872 17206 94924 17212
rect 94976 15978 95004 60030
rect 95148 57724 95200 57730
rect 95148 57666 95200 57672
rect 95056 57044 95108 57050
rect 95056 56986 95108 56992
rect 94964 15972 95016 15978
rect 94964 15914 95016 15920
rect 95068 7886 95096 56986
rect 95056 7880 95108 7886
rect 95056 7822 95108 7828
rect 93964 6886 94268 6914
rect 93676 4276 93728 4282
rect 93676 4218 93728 4224
rect 91560 3664 91612 3670
rect 91560 3606 91612 3612
rect 92388 3664 92440 3670
rect 92388 3606 92440 3612
rect 90640 3596 90692 3602
rect 90640 3538 90692 3544
rect 91572 480 91600 3606
rect 92756 2848 92808 2854
rect 92756 2790 92808 2796
rect 92768 480 92796 2790
rect 93964 480 93992 6886
rect 95160 4418 95188 57666
rect 95252 57594 95280 60044
rect 95240 57588 95292 57594
rect 95240 57530 95292 57536
rect 95528 57526 95556 60044
rect 95804 57730 95832 60044
rect 96094 60030 96384 60058
rect 96462 60030 96568 60058
rect 95792 57724 95844 57730
rect 95792 57666 95844 57672
rect 96356 57610 96384 60030
rect 96540 57746 96568 60030
rect 96540 57718 96660 57746
rect 96356 57582 96476 57610
rect 95516 57520 95568 57526
rect 95516 57462 95568 57468
rect 96344 57520 96396 57526
rect 96344 57462 96396 57468
rect 96356 7818 96384 57462
rect 96344 7812 96396 7818
rect 96344 7754 96396 7760
rect 96448 4554 96476 57582
rect 96528 57588 96580 57594
rect 96528 57530 96580 57536
rect 96436 4548 96488 4554
rect 96436 4490 96488 4496
rect 96540 4486 96568 57530
rect 96632 57254 96660 57718
rect 96724 57594 96752 60044
rect 96712 57588 96764 57594
rect 96712 57530 96764 57536
rect 96620 57248 96672 57254
rect 96620 57190 96672 57196
rect 97000 56914 97028 60044
rect 97276 57526 97304 60044
rect 97540 57724 97592 57730
rect 97540 57666 97592 57672
rect 97264 57520 97316 57526
rect 97264 57462 97316 57468
rect 96988 56908 97040 56914
rect 96988 56850 97040 56856
rect 97552 51746 97580 57666
rect 97540 51740 97592 51746
rect 97540 51682 97592 51688
rect 97644 18630 97672 60044
rect 97828 60030 97934 60058
rect 97724 57588 97776 57594
rect 97724 57530 97776 57536
rect 96620 18624 96672 18630
rect 96620 18566 96672 18572
rect 97632 18624 97684 18630
rect 97632 18566 97684 18572
rect 96632 16574 96660 18566
rect 97736 17338 97764 57530
rect 97724 17332 97776 17338
rect 97724 17274 97776 17280
rect 96632 16546 97488 16574
rect 96528 4480 96580 4486
rect 96528 4422 96580 4428
rect 95148 4412 95200 4418
rect 95148 4354 95200 4360
rect 95148 3052 95200 3058
rect 95148 2994 95200 3000
rect 95160 480 95188 2994
rect 96252 2984 96304 2990
rect 96252 2926 96304 2932
rect 96264 480 96292 2926
rect 97460 480 97488 16546
rect 97828 4758 97856 60030
rect 98196 57594 98224 60044
rect 98486 60030 98776 60058
rect 98184 57588 98236 57594
rect 98184 57530 98236 57536
rect 98644 57316 98696 57322
rect 98644 57258 98696 57264
rect 97908 56908 97960 56914
rect 97908 56850 97960 56856
rect 97816 4752 97868 4758
rect 97816 4694 97868 4700
rect 97920 4622 97948 56850
rect 97908 4616 97960 4622
rect 97908 4558 97960 4564
rect 98656 4214 98684 57258
rect 98748 55214 98776 60030
rect 98840 57118 98868 60044
rect 99130 60030 99236 60058
rect 99104 57588 99156 57594
rect 99104 57530 99156 57536
rect 98828 57112 98880 57118
rect 98828 57054 98880 57060
rect 98748 55186 99052 55214
rect 99024 16046 99052 55186
rect 99012 16040 99064 16046
rect 99012 15982 99064 15988
rect 99116 7750 99144 57530
rect 99104 7744 99156 7750
rect 99104 7686 99156 7692
rect 99208 7682 99236 60030
rect 99288 57112 99340 57118
rect 99288 57054 99340 57060
rect 99196 7676 99248 7682
rect 99196 7618 99248 7624
rect 99300 5506 99328 57054
rect 99392 55894 99420 60044
rect 99668 57730 99696 60044
rect 99656 57724 99708 57730
rect 99656 57666 99708 57672
rect 100036 57594 100064 60044
rect 100326 60030 100432 60058
rect 100602 60030 100708 60058
rect 100024 57588 100076 57594
rect 100024 57530 100076 57536
rect 99380 55888 99432 55894
rect 99380 55830 99432 55836
rect 99288 5500 99340 5506
rect 99288 5442 99340 5448
rect 98644 4208 98696 4214
rect 98644 4150 98696 4156
rect 100404 3466 100432 60030
rect 100576 57724 100628 57730
rect 100576 57666 100628 57672
rect 100484 57588 100536 57594
rect 100484 57530 100536 57536
rect 100496 7614 100524 57530
rect 100484 7608 100536 7614
rect 100484 7550 100536 7556
rect 100588 5438 100616 57666
rect 100680 57322 100708 60030
rect 100864 57458 100892 60044
rect 101232 57730 101260 60044
rect 101508 57798 101536 60044
rect 101798 60030 101996 60058
rect 101496 57792 101548 57798
rect 101496 57734 101548 57740
rect 101220 57724 101272 57730
rect 101220 57666 101272 57672
rect 101864 57724 101916 57730
rect 101864 57666 101916 57672
rect 101772 57588 101824 57594
rect 101772 57530 101824 57536
rect 100852 57452 100904 57458
rect 100852 57394 100904 57400
rect 101404 57384 101456 57390
rect 101404 57326 101456 57332
rect 100668 57316 100720 57322
rect 100668 57258 100720 57264
rect 100576 5432 100628 5438
rect 100576 5374 100628 5380
rect 101036 4208 101088 4214
rect 101036 4150 101088 4156
rect 99840 3460 99892 3466
rect 99840 3402 99892 3408
rect 100392 3460 100444 3466
rect 100392 3402 100444 3408
rect 98644 3188 98696 3194
rect 98644 3130 98696 3136
rect 98656 480 98684 3130
rect 99852 480 99880 3402
rect 101048 480 101076 4150
rect 101416 3058 101444 57326
rect 101784 9518 101812 57530
rect 101876 9586 101904 57666
rect 101864 9580 101916 9586
rect 101864 9522 101916 9528
rect 101772 9512 101824 9518
rect 101772 9454 101824 9460
rect 101968 5302 101996 60030
rect 102060 57594 102088 60044
rect 102048 57588 102100 57594
rect 102048 57530 102100 57536
rect 102336 57526 102364 60044
rect 102704 57594 102732 60044
rect 102994 60030 103192 60058
rect 102692 57588 102744 57594
rect 102692 57530 102744 57536
rect 102324 57520 102376 57526
rect 102324 57462 102376 57468
rect 102048 57452 102100 57458
rect 102048 57394 102100 57400
rect 102060 5370 102088 57394
rect 102876 57044 102928 57050
rect 102876 56986 102928 56992
rect 102784 56976 102836 56982
rect 102784 56918 102836 56924
rect 102048 5364 102100 5370
rect 102048 5306 102100 5312
rect 101956 5296 102008 5302
rect 101956 5238 102008 5244
rect 102232 3256 102284 3262
rect 102232 3198 102284 3204
rect 101404 3052 101456 3058
rect 101404 2994 101456 3000
rect 102244 480 102272 3198
rect 102796 3194 102824 56918
rect 102888 3262 102916 56986
rect 103164 55214 103192 60030
rect 103256 57458 103284 60044
rect 103428 57588 103480 57594
rect 103428 57530 103480 57536
rect 103244 57452 103296 57458
rect 103244 57394 103296 57400
rect 103164 55186 103376 55214
rect 103348 9450 103376 55186
rect 103336 9444 103388 9450
rect 103336 9386 103388 9392
rect 103440 5234 103468 57530
rect 103532 57390 103560 60044
rect 103900 57594 103928 60044
rect 103888 57588 103940 57594
rect 103888 57530 103940 57536
rect 103520 57384 103572 57390
rect 103520 57326 103572 57332
rect 104176 56914 104204 60044
rect 104466 60030 104572 60058
rect 104164 56908 104216 56914
rect 104164 56850 104216 56856
rect 103520 22772 103572 22778
rect 103520 22714 103572 22720
rect 103532 6914 103560 22714
rect 104544 9246 104572 60030
rect 104636 60030 104742 60058
rect 104636 9314 104664 60030
rect 104716 57588 104768 57594
rect 104716 57530 104768 57536
rect 104728 9382 104756 57530
rect 104808 57384 104860 57390
rect 104808 57326 104860 57332
rect 104716 9376 104768 9382
rect 104716 9318 104768 9324
rect 104624 9308 104676 9314
rect 104624 9250 104676 9256
rect 104532 9240 104584 9246
rect 104532 9182 104584 9188
rect 103532 6886 104572 6914
rect 103428 5228 103480 5234
rect 103428 5170 103480 5176
rect 102876 3256 102928 3262
rect 102876 3198 102928 3204
rect 102784 3188 102836 3194
rect 102784 3130 102836 3136
rect 103336 3120 103388 3126
rect 103336 3062 103388 3068
rect 103348 480 103376 3062
rect 104544 480 104572 6886
rect 104820 5166 104848 57326
rect 105096 57050 105124 60044
rect 105372 57594 105400 60044
rect 105452 57860 105504 57866
rect 105452 57802 105504 57808
rect 105360 57588 105412 57594
rect 105360 57530 105412 57536
rect 105084 57044 105136 57050
rect 105084 56986 105136 56992
rect 105464 55214 105492 57802
rect 105544 57180 105596 57186
rect 105544 57122 105596 57128
rect 105556 56794 105584 57122
rect 105648 56982 105676 60044
rect 105938 60030 106044 60058
rect 105636 56976 105688 56982
rect 105636 56918 105688 56924
rect 105556 56766 105676 56794
rect 105464 55186 105584 55214
rect 104808 5160 104860 5166
rect 104808 5102 104860 5108
rect 105556 4214 105584 55186
rect 105648 6322 105676 56766
rect 106016 14482 106044 60030
rect 106292 57866 106320 60044
rect 106280 57860 106332 57866
rect 106280 57802 106332 57808
rect 106568 57594 106596 60044
rect 106188 57588 106240 57594
rect 106188 57530 106240 57536
rect 106556 57588 106608 57594
rect 106556 57530 106608 57536
rect 106096 56976 106148 56982
rect 106096 56918 106148 56924
rect 106004 14476 106056 14482
rect 106004 14418 106056 14424
rect 106108 9110 106136 56918
rect 106200 9178 106228 57530
rect 106844 57050 106872 60044
rect 107134 60030 107332 60058
rect 106832 57044 106884 57050
rect 106832 56986 106884 56992
rect 107304 11014 107332 60030
rect 107396 60030 107502 60058
rect 107292 11008 107344 11014
rect 107292 10950 107344 10956
rect 107396 10946 107424 60030
rect 107568 57860 107620 57866
rect 107568 57802 107620 57808
rect 107476 57588 107528 57594
rect 107476 57530 107528 57536
rect 107384 10940 107436 10946
rect 107384 10882 107436 10888
rect 106924 10328 106976 10334
rect 106924 10270 106976 10276
rect 106188 9172 106240 9178
rect 106188 9114 106240 9120
rect 106096 9104 106148 9110
rect 106096 9046 106148 9052
rect 105636 6316 105688 6322
rect 105636 6258 105688 6264
rect 105544 4208 105596 4214
rect 105544 4150 105596 4156
rect 106936 3330 106964 10270
rect 107488 8974 107516 57530
rect 107580 9042 107608 57802
rect 107764 57186 107792 60044
rect 107752 57180 107804 57186
rect 107752 57122 107804 57128
rect 108040 57118 108068 60044
rect 108330 60030 108528 60058
rect 108606 60030 108896 60058
rect 108500 57610 108528 60030
rect 108500 57582 108804 57610
rect 108580 57384 108632 57390
rect 108580 57326 108632 57332
rect 108028 57112 108080 57118
rect 108028 57054 108080 57060
rect 108592 10674 108620 57326
rect 108672 57112 108724 57118
rect 108672 57054 108724 57060
rect 108684 10878 108712 57054
rect 108672 10872 108724 10878
rect 108672 10814 108724 10820
rect 108776 10810 108804 57582
rect 108764 10804 108816 10810
rect 108764 10746 108816 10752
rect 108580 10668 108632 10674
rect 108580 10610 108632 10616
rect 107568 9036 107620 9042
rect 107568 8978 107620 8984
rect 107476 8968 107528 8974
rect 107476 8910 107528 8916
rect 108868 5030 108896 60030
rect 108960 57390 108988 60044
rect 109236 57390 109264 60044
rect 109512 57866 109540 60044
rect 109500 57860 109552 57866
rect 109500 57802 109552 57808
rect 109788 57594 109816 60044
rect 110064 60030 110170 60058
rect 109776 57588 109828 57594
rect 109776 57530 109828 57536
rect 108948 57384 109000 57390
rect 108948 57326 109000 57332
rect 109224 57384 109276 57390
rect 109224 57326 109276 57332
rect 108948 57180 109000 57186
rect 108948 57122 109000 57128
rect 108960 5098 108988 57122
rect 110064 10538 110092 60030
rect 110328 57860 110380 57866
rect 110328 57802 110380 57808
rect 110144 57588 110196 57594
rect 110144 57530 110196 57536
rect 110156 10606 110184 57530
rect 110236 57384 110288 57390
rect 110236 57326 110288 57332
rect 110248 10742 110276 57326
rect 110236 10736 110288 10742
rect 110236 10678 110288 10684
rect 110144 10600 110196 10606
rect 110144 10542 110196 10548
rect 110052 10532 110104 10538
rect 110052 10474 110104 10480
rect 108948 5092 109000 5098
rect 108948 5034 109000 5040
rect 108856 5024 108908 5030
rect 108856 4966 108908 4972
rect 110340 4962 110368 57802
rect 110432 57050 110460 60044
rect 110708 57390 110736 60044
rect 110998 60030 111288 60058
rect 111366 60030 111564 60058
rect 111642 60030 111748 60058
rect 111260 57610 111288 60030
rect 111536 57746 111564 60030
rect 111536 57718 111656 57746
rect 111260 57582 111564 57610
rect 110696 57384 110748 57390
rect 110696 57326 110748 57332
rect 111432 57384 111484 57390
rect 111432 57326 111484 57332
rect 111340 57180 111392 57186
rect 111340 57122 111392 57128
rect 110420 57044 110472 57050
rect 110420 56986 110472 56992
rect 111352 10334 111380 57122
rect 111444 10402 111472 57326
rect 111536 10470 111564 57582
rect 111524 10464 111576 10470
rect 111524 10406 111576 10412
rect 111432 10396 111484 10402
rect 111432 10338 111484 10344
rect 111340 10328 111392 10334
rect 111340 10270 111392 10276
rect 110328 4956 110380 4962
rect 110328 4898 110380 4904
rect 111628 4826 111656 57718
rect 111720 57186 111748 60030
rect 111904 57594 111932 60044
rect 111892 57588 111944 57594
rect 111892 57530 111944 57536
rect 111708 57180 111760 57186
rect 111708 57122 111760 57128
rect 111708 57044 111760 57050
rect 111708 56986 111760 56992
rect 111720 4894 111748 56986
rect 112180 55418 112208 60044
rect 112562 60030 112760 60058
rect 112838 60030 112944 60058
rect 112444 56024 112496 56030
rect 112444 55966 112496 55972
rect 112168 55412 112220 55418
rect 112168 55354 112220 55360
rect 111708 4888 111760 4894
rect 111708 4830 111760 4836
rect 111616 4820 111668 4826
rect 111616 4762 111668 4768
rect 108120 4208 108172 4214
rect 108120 4150 108172 4156
rect 105728 3324 105780 3330
rect 105728 3266 105780 3272
rect 106924 3324 106976 3330
rect 106924 3266 106976 3272
rect 105740 480 105768 3266
rect 106924 3052 106976 3058
rect 106924 2994 106976 3000
rect 106936 480 106964 2994
rect 108132 480 108160 4150
rect 112456 4146 112484 55966
rect 112732 55214 112760 60030
rect 112732 55186 112852 55214
rect 112824 9790 112852 55186
rect 112916 15366 112944 60030
rect 112996 57588 113048 57594
rect 112996 57530 113048 57536
rect 113008 15910 113036 57530
rect 113100 55554 113128 60044
rect 113376 57186 113404 60044
rect 113758 60030 113956 60058
rect 113364 57180 113416 57186
rect 113364 57122 113416 57128
rect 113088 55548 113140 55554
rect 113088 55490 113140 55496
rect 113928 55214 113956 60030
rect 114020 56778 114048 60044
rect 114310 60030 114416 60058
rect 114008 56772 114060 56778
rect 114008 56714 114060 56720
rect 113928 55186 114324 55214
rect 112996 15904 113048 15910
rect 112996 15846 113048 15852
rect 114296 15434 114324 55186
rect 114284 15428 114336 15434
rect 114284 15370 114336 15376
rect 112904 15360 112956 15366
rect 112904 15302 112956 15308
rect 114388 10130 114416 60030
rect 114468 57180 114520 57186
rect 114468 57122 114520 57128
rect 114376 10124 114428 10130
rect 114376 10066 114428 10072
rect 114480 9858 114508 57122
rect 114572 57118 114600 60044
rect 114560 57112 114612 57118
rect 114560 57054 114612 57060
rect 114940 55622 114968 60044
rect 115230 60030 115428 60058
rect 114928 55616 114980 55622
rect 114928 55558 114980 55564
rect 115400 55214 115428 60030
rect 115492 57186 115520 60044
rect 115584 60030 115782 60058
rect 115480 57180 115532 57186
rect 115480 57122 115532 57128
rect 115400 55186 115520 55214
rect 115204 15972 115256 15978
rect 115204 15914 115256 15920
rect 114468 9852 114520 9858
rect 114468 9794 114520 9800
rect 112812 9784 112864 9790
rect 112812 9726 112864 9732
rect 112444 4140 112496 4146
rect 112444 4082 112496 4088
rect 115216 4078 115244 15914
rect 115492 9926 115520 55186
rect 115584 18494 115612 60030
rect 116044 57186 116072 60044
rect 115756 57180 115808 57186
rect 115756 57122 115808 57128
rect 116032 57180 116084 57186
rect 116032 57122 116084 57128
rect 115664 57112 115716 57118
rect 115664 57054 115716 57060
rect 115572 18488 115624 18494
rect 115572 18430 115624 18436
rect 115676 15502 115704 57054
rect 115768 15570 115796 57122
rect 116412 56914 116440 60044
rect 116400 56908 116452 56914
rect 116400 56850 116452 56856
rect 116688 55690 116716 60044
rect 116860 57180 116912 57186
rect 116860 57122 116912 57128
rect 116676 55684 116728 55690
rect 116676 55626 116728 55632
rect 116584 16040 116636 16046
rect 116584 15982 116636 15988
rect 115756 15564 115808 15570
rect 115756 15506 115808 15512
rect 115664 15496 115716 15502
rect 115664 15438 115716 15444
rect 115480 9920 115532 9926
rect 115480 9862 115532 9868
rect 112812 4072 112864 4078
rect 112812 4014 112864 4020
rect 115204 4072 115256 4078
rect 115204 4014 115256 4020
rect 109316 3392 109368 3398
rect 109316 3334 109368 3340
rect 109328 480 109356 3334
rect 111616 3324 111668 3330
rect 111616 3266 111668 3272
rect 110512 3188 110564 3194
rect 110512 3130 110564 3136
rect 110524 480 110552 3130
rect 111628 480 111656 3266
rect 112824 480 112852 4014
rect 116596 3534 116624 15982
rect 116872 9994 116900 57122
rect 116964 57050 116992 60044
rect 117056 60030 117254 60058
rect 116952 57044 117004 57050
rect 116952 56986 117004 56992
rect 116952 56908 117004 56914
rect 116952 56850 117004 56856
rect 116964 15638 116992 56850
rect 117056 15706 117084 60030
rect 117136 57044 117188 57050
rect 117136 56986 117188 56992
rect 117044 15700 117096 15706
rect 117044 15642 117096 15648
rect 116952 15632 117004 15638
rect 116952 15574 117004 15580
rect 117148 10062 117176 56986
rect 117608 56982 117636 60044
rect 117700 60030 117898 60058
rect 118174 60030 118372 60058
rect 117596 56976 117648 56982
rect 117596 56918 117648 56924
rect 117700 52766 117728 60030
rect 118344 55214 118372 60030
rect 118436 56914 118464 60044
rect 118818 60030 118924 60058
rect 118424 56908 118476 56914
rect 118424 56850 118476 56856
rect 118344 55186 118648 55214
rect 117688 52760 117740 52766
rect 117688 52702 117740 52708
rect 118620 15774 118648 55186
rect 118896 52834 118924 60030
rect 119080 57118 119108 60044
rect 119370 60030 119568 60058
rect 119252 57180 119304 57186
rect 119252 57122 119304 57128
rect 119068 57112 119120 57118
rect 119068 57054 119120 57060
rect 118884 52828 118936 52834
rect 118884 52770 118936 52776
rect 119264 51542 119292 57122
rect 119540 55214 119568 60030
rect 119632 57186 119660 60044
rect 119816 60030 120014 60058
rect 119620 57180 119672 57186
rect 119620 57122 119672 57128
rect 119540 55186 119660 55214
rect 119252 51536 119304 51542
rect 119252 51478 119304 51484
rect 119344 17332 119396 17338
rect 119344 17274 119396 17280
rect 118608 15768 118660 15774
rect 118608 15710 118660 15716
rect 117136 10056 117188 10062
rect 117136 9998 117188 10004
rect 116860 9988 116912 9994
rect 116860 9930 116912 9936
rect 117596 3936 117648 3942
rect 117596 3878 117648 3884
rect 116400 3528 116452 3534
rect 116400 3470 116452 3476
rect 116584 3528 116636 3534
rect 116584 3470 116636 3476
rect 115204 3324 115256 3330
rect 115204 3266 115256 3272
rect 114008 3256 114060 3262
rect 114008 3198 114060 3204
rect 114020 480 114048 3198
rect 115216 480 115244 3266
rect 116412 480 116440 3470
rect 117608 480 117636 3878
rect 119356 3874 119384 17274
rect 119632 5642 119660 55186
rect 119816 16590 119844 60030
rect 119896 57112 119948 57118
rect 119896 57054 119948 57060
rect 119804 16584 119856 16590
rect 119804 16526 119856 16532
rect 119908 15842 119936 57054
rect 120276 57050 120304 60044
rect 120552 57118 120580 60044
rect 120842 60030 121132 60058
rect 121210 60030 121408 60058
rect 120540 57112 120592 57118
rect 120540 57054 120592 57060
rect 120264 57044 120316 57050
rect 120264 56986 120316 56992
rect 121104 55214 121132 60030
rect 121276 57044 121328 57050
rect 121276 56986 121328 56992
rect 121104 55186 121224 55214
rect 121196 16522 121224 55186
rect 121184 16516 121236 16522
rect 121184 16458 121236 16464
rect 119896 15836 119948 15842
rect 119896 15778 119948 15784
rect 121288 5710 121316 56986
rect 121380 5778 121408 60030
rect 121472 57050 121500 60044
rect 121748 57186 121776 60044
rect 121736 57180 121788 57186
rect 121736 57122 121788 57128
rect 121460 57044 121512 57050
rect 121460 56986 121512 56992
rect 122024 56846 122052 60044
rect 122314 60030 122512 60058
rect 122012 56840 122064 56846
rect 122012 56782 122064 56788
rect 122484 18562 122512 60030
rect 122564 57180 122616 57186
rect 122564 57122 122616 57128
rect 122472 18556 122524 18562
rect 122472 18498 122524 18504
rect 122104 17264 122156 17270
rect 122104 17206 122156 17212
rect 121368 5772 121420 5778
rect 121368 5714 121420 5720
rect 121276 5704 121328 5710
rect 121276 5646 121328 5652
rect 119620 5636 119672 5642
rect 119620 5578 119672 5584
rect 119896 4004 119948 4010
rect 119896 3946 119948 3952
rect 118792 3868 118844 3874
rect 118792 3810 118844 3816
rect 119344 3868 119396 3874
rect 119344 3810 119396 3816
rect 118804 480 118832 3810
rect 119908 480 119936 3946
rect 122116 3806 122144 17206
rect 122576 16454 122604 57122
rect 122564 16448 122616 16454
rect 122564 16390 122616 16396
rect 122668 16386 122696 60044
rect 122748 56840 122800 56846
rect 122748 56782 122800 56788
rect 122656 16380 122708 16386
rect 122656 16322 122708 16328
rect 122760 5846 122788 56782
rect 122944 56778 122972 60044
rect 122932 56772 122984 56778
rect 122932 56714 122984 56720
rect 123024 56704 123076 56710
rect 123024 56646 123076 56652
rect 123036 51610 123064 56646
rect 123220 52902 123248 60044
rect 123496 57662 123524 60044
rect 123772 60030 123878 60058
rect 123484 57656 123536 57662
rect 123484 57598 123536 57604
rect 123208 52896 123260 52902
rect 123208 52838 123260 52844
rect 123024 51604 123076 51610
rect 123024 51546 123076 51552
rect 123772 5982 123800 60030
rect 123944 57656 123996 57662
rect 123944 57598 123996 57604
rect 123956 16318 123984 57598
rect 124036 56772 124088 56778
rect 124036 56714 124088 56720
rect 123944 16312 123996 16318
rect 123944 16254 123996 16260
rect 123760 5976 123812 5982
rect 123760 5918 123812 5924
rect 124048 5914 124076 56714
rect 124140 56710 124168 60044
rect 124416 56778 124444 60044
rect 124706 60030 124996 60058
rect 124864 57792 124916 57798
rect 124864 57734 124916 57740
rect 124404 56772 124456 56778
rect 124404 56714 124456 56720
rect 124128 56704 124180 56710
rect 124128 56646 124180 56652
rect 124220 56704 124272 56710
rect 124220 56646 124272 56652
rect 124232 52970 124260 56646
rect 124220 52964 124272 52970
rect 124220 52906 124272 52912
rect 124036 5908 124088 5914
rect 124036 5850 124088 5856
rect 122748 5840 122800 5846
rect 122748 5782 122800 5788
rect 121092 3800 121144 3806
rect 121092 3742 121144 3748
rect 122104 3800 122156 3806
rect 122104 3742 122156 3748
rect 121104 480 121132 3742
rect 122288 3732 122340 3738
rect 122288 3674 122340 3680
rect 122300 480 122328 3674
rect 124680 3664 124732 3670
rect 124680 3606 124732 3612
rect 123484 3596 123536 3602
rect 123484 3538 123536 3544
rect 123496 480 123524 3538
rect 124692 480 124720 3606
rect 124876 3602 124904 57734
rect 124968 55214 124996 60030
rect 125060 56710 125088 60044
rect 125350 60030 125456 60058
rect 125324 56772 125376 56778
rect 125324 56714 125376 56720
rect 125048 56704 125100 56710
rect 125048 56646 125100 56652
rect 124968 55186 125272 55214
rect 125244 6050 125272 55186
rect 125336 17134 125364 56714
rect 125428 17202 125456 60030
rect 125612 57798 125640 60044
rect 125600 57792 125652 57798
rect 125600 57734 125652 57740
rect 125888 57730 125916 60044
rect 126270 60030 126468 60058
rect 125876 57724 125928 57730
rect 125876 57666 125928 57672
rect 126440 55214 126468 60030
rect 126532 57662 126560 60044
rect 126624 60030 126822 60058
rect 126520 57656 126572 57662
rect 126520 57598 126572 57604
rect 126440 55186 126560 55214
rect 126532 17950 126560 55186
rect 126520 17944 126572 17950
rect 126520 17886 126572 17892
rect 125416 17196 125468 17202
rect 125416 17138 125468 17144
rect 125324 17128 125376 17134
rect 125324 17070 125376 17076
rect 126624 11286 126652 60030
rect 126888 57792 126940 57798
rect 126888 57734 126940 57740
rect 126704 57724 126756 57730
rect 126704 57666 126756 57672
rect 126612 11280 126664 11286
rect 126612 11222 126664 11228
rect 126716 11218 126744 57666
rect 126796 57656 126848 57662
rect 126796 57598 126848 57604
rect 126704 11212 126756 11218
rect 126704 11154 126756 11160
rect 126808 6866 126836 57598
rect 126796 6860 126848 6866
rect 126796 6802 126848 6808
rect 126900 6118 126928 57734
rect 127084 57662 127112 60044
rect 127452 57798 127480 60044
rect 127440 57792 127492 57798
rect 127440 57734 127492 57740
rect 127728 57730 127756 60044
rect 127716 57724 127768 57730
rect 127716 57666 127768 57672
rect 127072 57656 127124 57662
rect 127072 57598 127124 57604
rect 127900 57656 127952 57662
rect 127900 57598 127952 57604
rect 127912 17882 127940 57598
rect 127900 17876 127952 17882
rect 127900 17818 127952 17824
rect 128004 17814 128032 60044
rect 128176 57792 128228 57798
rect 128176 57734 128228 57740
rect 128084 57724 128136 57730
rect 128084 57666 128136 57672
rect 127992 17808 128044 17814
rect 127992 17750 128044 17756
rect 128096 11354 128124 57666
rect 128084 11348 128136 11354
rect 128084 11290 128136 11296
rect 128188 6798 128216 57734
rect 128176 6792 128228 6798
rect 128176 6734 128228 6740
rect 128280 6730 128308 60044
rect 128648 57662 128676 60044
rect 128938 60030 129136 60058
rect 128636 57656 128688 57662
rect 128636 57598 128688 57604
rect 129004 56908 129056 56914
rect 129004 56850 129056 56856
rect 128268 6724 128320 6730
rect 128268 6666 128320 6672
rect 128176 6316 128228 6322
rect 128176 6258 128228 6264
rect 126888 6112 126940 6118
rect 126888 6054 126940 6060
rect 125232 6044 125284 6050
rect 125232 5986 125284 5992
rect 126980 4344 127032 4350
rect 126980 4286 127032 4292
rect 124864 3596 124916 3602
rect 124864 3538 124916 3544
rect 125876 3596 125928 3602
rect 125876 3538 125928 3544
rect 125888 480 125916 3538
rect 126992 480 127020 4286
rect 128188 480 128216 6258
rect 129016 3806 129044 56850
rect 129108 55214 129136 60030
rect 129200 56778 129228 60044
rect 129188 56772 129240 56778
rect 129188 56714 129240 56720
rect 129108 55186 129412 55214
rect 129384 17746 129412 55186
rect 129372 17740 129424 17746
rect 129372 17682 129424 17688
rect 129476 11490 129504 60044
rect 129766 60030 130056 60058
rect 129556 57656 129608 57662
rect 129556 57598 129608 57604
rect 129464 11484 129516 11490
rect 129464 11426 129516 11432
rect 129568 11422 129596 57598
rect 130028 56914 130056 60030
rect 130120 57730 130148 60044
rect 130108 57724 130160 57730
rect 130108 57666 130160 57672
rect 130396 57662 130424 60044
rect 130686 60030 130792 60058
rect 130962 60030 131068 60058
rect 130384 57656 130436 57662
rect 130384 57598 130436 57604
rect 130016 56908 130068 56914
rect 130016 56850 130068 56856
rect 129740 56840 129792 56846
rect 129740 56782 129792 56788
rect 129648 56772 129700 56778
rect 129648 56714 129700 56720
rect 129556 11416 129608 11422
rect 129556 11358 129608 11364
rect 129660 6662 129688 56714
rect 129752 55350 129780 56782
rect 129740 55344 129792 55350
rect 129740 55286 129792 55292
rect 130764 17678 130792 60030
rect 130936 57724 130988 57730
rect 130936 57666 130988 57672
rect 130844 57656 130896 57662
rect 130844 57598 130896 57604
rect 130752 17672 130804 17678
rect 130752 17614 130804 17620
rect 130856 11558 130884 57598
rect 130844 11552 130896 11558
rect 130844 11494 130896 11500
rect 129648 6656 129700 6662
rect 129648 6598 129700 6604
rect 130948 6594 130976 57666
rect 130936 6588 130988 6594
rect 130936 6530 130988 6536
rect 131040 6526 131068 60030
rect 131316 57730 131344 60044
rect 131592 57798 131620 60044
rect 131580 57792 131632 57798
rect 131580 57734 131632 57740
rect 131304 57724 131356 57730
rect 131304 57666 131356 57672
rect 131868 57662 131896 60044
rect 132158 60030 132356 60058
rect 132224 57724 132276 57730
rect 132224 57666 132276 57672
rect 131856 57656 131908 57662
rect 131856 57598 131908 57604
rect 132236 11626 132264 57666
rect 132328 11694 132356 60030
rect 132512 57730 132540 60044
rect 132500 57724 132552 57730
rect 132500 57666 132552 57672
rect 132788 57662 132816 60044
rect 133078 60030 133276 60058
rect 133144 57860 133196 57866
rect 133144 57802 133196 57808
rect 132408 57656 132460 57662
rect 132408 57598 132460 57604
rect 132776 57656 132828 57662
rect 132776 57598 132828 57604
rect 132316 11688 132368 11694
rect 132316 11630 132368 11636
rect 132224 11620 132276 11626
rect 132224 11562 132276 11568
rect 131028 6520 131080 6526
rect 131028 6462 131080 6468
rect 132420 6458 132448 57598
rect 132408 6452 132460 6458
rect 132408 6394 132460 6400
rect 130568 6248 130620 6254
rect 130568 6190 130620 6196
rect 129372 4276 129424 4282
rect 129372 4218 129424 4224
rect 129004 3800 129056 3806
rect 129004 3742 129056 3748
rect 129384 480 129412 4218
rect 130580 480 130608 6190
rect 133156 4690 133184 57802
rect 133248 55214 133276 60030
rect 133340 56642 133368 60044
rect 133722 60030 133828 60058
rect 133696 57656 133748 57662
rect 133696 57598 133748 57604
rect 133512 56976 133564 56982
rect 133512 56918 133564 56924
rect 133328 56636 133380 56642
rect 133328 56578 133380 56584
rect 133524 55486 133552 56918
rect 133512 55480 133564 55486
rect 133512 55422 133564 55428
rect 133248 55186 133644 55214
rect 133616 12442 133644 55186
rect 133604 12436 133656 12442
rect 133604 12378 133656 12384
rect 133708 6390 133736 57598
rect 133696 6384 133748 6390
rect 133696 6326 133748 6332
rect 133800 6322 133828 60030
rect 133984 56846 134012 60044
rect 134274 60030 134472 60058
rect 134064 57180 134116 57186
rect 134064 57122 134116 57128
rect 133972 56840 134024 56846
rect 133972 56782 134024 56788
rect 134076 54194 134104 57122
rect 134444 56710 134472 60030
rect 134536 57594 134564 60044
rect 134918 60030 135024 60058
rect 134524 57588 134576 57594
rect 134524 57530 134576 57536
rect 134248 56704 134300 56710
rect 134248 56646 134300 56652
rect 134432 56704 134484 56710
rect 134432 56646 134484 56652
rect 134260 55214 134288 56646
rect 134260 55186 134564 55214
rect 134064 54188 134116 54194
rect 134064 54130 134116 54136
rect 133788 6316 133840 6322
rect 133788 6258 133840 6264
rect 134156 6180 134208 6186
rect 134156 6122 134208 6128
rect 132960 4684 133012 4690
rect 132960 4626 133012 4632
rect 133144 4684 133196 4690
rect 133144 4626 133196 4632
rect 131764 4140 131816 4146
rect 131764 4082 131816 4088
rect 131776 480 131804 4082
rect 132972 480 133000 4626
rect 134168 480 134196 6122
rect 134536 3670 134564 55186
rect 134996 12306 135024 60030
rect 135180 57746 135208 60044
rect 135180 57718 135300 57746
rect 135272 57662 135300 57718
rect 135260 57656 135312 57662
rect 135260 57598 135312 57604
rect 135168 57588 135220 57594
rect 135168 57530 135220 57536
rect 135076 56840 135128 56846
rect 135076 56782 135128 56788
rect 135088 12374 135116 56782
rect 135076 12368 135128 12374
rect 135076 12310 135128 12316
rect 134984 12300 135036 12306
rect 134984 12242 135036 12248
rect 135180 6254 135208 57530
rect 135456 57526 135484 60044
rect 135732 57594 135760 60044
rect 136008 57798 136036 60044
rect 136390 60030 136588 60058
rect 135996 57792 136048 57798
rect 135996 57734 136048 57740
rect 136560 57610 136588 60030
rect 136652 57730 136680 60044
rect 136732 57860 136784 57866
rect 136732 57802 136784 57808
rect 136640 57724 136692 57730
rect 136640 57666 136692 57672
rect 135720 57588 135772 57594
rect 135720 57530 135772 57536
rect 136456 57588 136508 57594
rect 136560 57582 136680 57610
rect 136456 57530 136508 57536
rect 135444 57520 135496 57526
rect 135444 57462 135496 57468
rect 136468 12238 136496 57530
rect 136548 57520 136600 57526
rect 136548 57462 136600 57468
rect 136456 12232 136508 12238
rect 136456 12174 136508 12180
rect 135168 6248 135220 6254
rect 135168 6190 135220 6196
rect 136560 6186 136588 57462
rect 136652 54262 136680 57582
rect 136744 56642 136772 57802
rect 136928 57186 136956 60044
rect 136916 57180 136968 57186
rect 136916 57122 136968 57128
rect 136732 56636 136784 56642
rect 136732 56578 136784 56584
rect 137204 54330 137232 60044
rect 137586 60030 137784 60058
rect 137862 60030 137968 60058
rect 137284 57112 137336 57118
rect 137284 57054 137336 57060
rect 137192 54324 137244 54330
rect 137192 54266 137244 54272
rect 136640 54256 136692 54262
rect 136640 54198 136692 54204
rect 136548 6180 136600 6186
rect 136548 6122 136600 6128
rect 136456 4412 136508 4418
rect 136456 4354 136508 4360
rect 135260 3732 135312 3738
rect 135260 3674 135312 3680
rect 134524 3664 134576 3670
rect 134524 3606 134576 3612
rect 135272 480 135300 3674
rect 136468 480 136496 4354
rect 137296 3602 137324 57054
rect 137756 12102 137784 60030
rect 137836 57724 137888 57730
rect 137836 57666 137888 57672
rect 137848 12170 137876 57666
rect 137940 56914 137968 60030
rect 138124 57866 138152 60044
rect 138112 57860 138164 57866
rect 138112 57802 138164 57808
rect 137928 56908 137980 56914
rect 137928 56850 137980 56856
rect 138400 56642 138428 60044
rect 138768 57866 138796 60044
rect 138756 57860 138808 57866
rect 138756 57802 138808 57808
rect 137928 56636 137980 56642
rect 137928 56578 137980 56584
rect 138388 56636 138440 56642
rect 138388 56578 138440 56584
rect 137940 50250 137968 56578
rect 139044 54466 139072 60044
rect 139228 60030 139334 60058
rect 139124 56636 139176 56642
rect 139124 56578 139176 56584
rect 139032 54460 139084 54466
rect 139032 54402 139084 54408
rect 137928 50244 137980 50250
rect 137928 50186 137980 50192
rect 137836 12164 137888 12170
rect 137836 12106 137888 12112
rect 137744 12096 137796 12102
rect 137744 12038 137796 12044
rect 139136 12034 139164 56578
rect 139124 12028 139176 12034
rect 139124 11970 139176 11976
rect 139228 11966 139256 60030
rect 139596 56642 139624 60044
rect 139676 56772 139728 56778
rect 139676 56714 139728 56720
rect 139584 56636 139636 56642
rect 139584 56578 139636 56584
rect 139688 49570 139716 56714
rect 139964 55214 139992 60044
rect 140254 60030 140452 60058
rect 140320 57792 140372 57798
rect 140320 57734 140372 57740
rect 140044 56840 140096 56846
rect 140044 56782 140096 56788
rect 139952 55208 140004 55214
rect 139952 55150 140004 55156
rect 139676 49564 139728 49570
rect 139676 49506 139728 49512
rect 140056 16574 140084 56782
rect 140332 54398 140360 57734
rect 140320 54392 140372 54398
rect 140320 54334 140372 54340
rect 140424 51074 140452 60030
rect 140516 57798 140544 60044
rect 140504 57792 140556 57798
rect 140504 57734 140556 57740
rect 140792 55146 140820 60044
rect 141160 56642 141188 60044
rect 141332 57112 141384 57118
rect 141332 57054 141384 57060
rect 140872 56636 140924 56642
rect 140872 56578 140924 56584
rect 141148 56636 141200 56642
rect 141148 56578 141200 56584
rect 140780 55140 140832 55146
rect 140780 55082 140832 55088
rect 140424 51046 140728 51074
rect 140056 16546 140176 16574
rect 139216 11960 139268 11966
rect 139216 11902 139268 11908
rect 137652 7880 137704 7886
rect 137652 7822 137704 7828
rect 137284 3596 137336 3602
rect 137284 3538 137336 3544
rect 137664 480 137692 7822
rect 140148 4486 140176 16546
rect 140700 11898 140728 51046
rect 140884 49230 140912 56578
rect 141344 51074 141372 57054
rect 141436 56982 141464 60044
rect 141424 56976 141476 56982
rect 141424 56918 141476 56924
rect 141712 55078 141740 60044
rect 141804 60030 142002 60058
rect 141700 55072 141752 55078
rect 141700 55014 141752 55020
rect 141344 51046 141464 51074
rect 140872 49224 140924 49230
rect 140872 49166 140924 49172
rect 140688 11892 140740 11898
rect 140688 11834 140740 11840
rect 141240 7812 141292 7818
rect 141240 7754 141292 7760
rect 140044 4480 140096 4486
rect 140044 4422 140096 4428
rect 140136 4480 140188 4486
rect 140136 4422 140188 4428
rect 138848 4072 138900 4078
rect 138848 4014 138900 4020
rect 138860 480 138888 4014
rect 140056 480 140084 4422
rect 141252 480 141280 7754
rect 141436 4146 141464 51046
rect 141804 11762 141832 60030
rect 142356 57254 142384 60044
rect 142540 60030 142646 60058
rect 142922 60030 143120 60058
rect 142252 57248 142304 57254
rect 142252 57190 142304 57196
rect 142344 57248 142396 57254
rect 142344 57190 142396 57196
rect 141976 56636 142028 56642
rect 141976 56578 142028 56584
rect 141988 11830 142016 56578
rect 142160 51740 142212 51746
rect 142160 51682 142212 51688
rect 142172 16574 142200 51682
rect 142264 51474 142292 57190
rect 142540 55010 142568 60030
rect 142804 57588 142856 57594
rect 142804 57530 142856 57536
rect 142816 57474 142844 57530
rect 142620 57452 142672 57458
rect 142816 57446 143028 57474
rect 142620 57394 142672 57400
rect 142528 55004 142580 55010
rect 142528 54946 142580 54952
rect 142252 51468 142304 51474
rect 142252 51410 142304 51416
rect 142632 51074 142660 57394
rect 142712 57044 142764 57050
rect 142712 56986 142764 56992
rect 142724 56896 142752 56986
rect 142724 56868 142936 56896
rect 142632 51046 142844 51074
rect 142172 16546 142476 16574
rect 141976 11824 142028 11830
rect 141976 11766 142028 11772
rect 141792 11756 141844 11762
rect 141792 11698 141844 11704
rect 141424 4140 141476 4146
rect 141424 4082 141476 4088
rect 142448 480 142476 16546
rect 142816 3738 142844 51046
rect 142908 17066 142936 56868
rect 143000 17474 143028 57446
rect 143092 57118 143120 60030
rect 143184 57458 143212 60044
rect 143172 57452 143224 57458
rect 143172 57394 143224 57400
rect 143080 57112 143132 57118
rect 143080 57054 143132 57060
rect 143460 53038 143488 60044
rect 143828 56642 143856 60044
rect 144104 57322 144132 60044
rect 144394 60030 144592 60058
rect 144184 57384 144236 57390
rect 144184 57326 144236 57332
rect 144092 57316 144144 57322
rect 144092 57258 144144 57264
rect 143816 56636 143868 56642
rect 143816 56578 143868 56584
rect 143448 53032 143500 53038
rect 143448 52974 143500 52980
rect 142988 17468 143040 17474
rect 142988 17410 143040 17416
rect 142896 17060 142948 17066
rect 142896 17002 142948 17008
rect 143540 4548 143592 4554
rect 143540 4490 143592 4496
rect 142804 3732 142856 3738
rect 142804 3674 142856 3680
rect 143552 480 143580 4490
rect 144196 3942 144224 57326
rect 144368 57112 144420 57118
rect 144368 57054 144420 57060
rect 144380 51678 144408 57054
rect 144460 56636 144512 56642
rect 144460 56578 144512 56584
rect 144368 51672 144420 51678
rect 144368 51614 144420 51620
rect 144472 51074 144500 56578
rect 144564 52306 144592 60030
rect 144656 52426 144684 60044
rect 145024 57390 145052 60044
rect 145012 57384 145064 57390
rect 145012 57326 145064 57332
rect 145300 56642 145328 60044
rect 145288 56636 145340 56642
rect 145288 56578 145340 56584
rect 144644 52420 144696 52426
rect 144644 52362 144696 52368
rect 145576 52358 145604 60044
rect 145852 57730 145880 60044
rect 146128 60030 146234 60058
rect 145840 57724 145892 57730
rect 145840 57666 145892 57672
rect 145564 52352 145616 52358
rect 144564 52278 144868 52306
rect 145564 52294 145616 52300
rect 144472 51046 144776 51074
rect 144748 17338 144776 51046
rect 144736 17332 144788 17338
rect 144736 17274 144788 17280
rect 144840 7070 144868 52278
rect 146128 7206 146156 60030
rect 146208 56636 146260 56642
rect 146208 56578 146260 56584
rect 146116 7200 146168 7206
rect 146116 7142 146168 7148
rect 146220 7138 146248 56578
rect 146496 52290 146524 60044
rect 146772 57118 146800 60044
rect 147062 60030 147352 60058
rect 147220 57656 147272 57662
rect 147220 57598 147272 57604
rect 147036 57520 147088 57526
rect 147036 57462 147088 57468
rect 146760 57112 146812 57118
rect 146760 57054 146812 57060
rect 146944 56840 146996 56846
rect 146944 56782 146996 56788
rect 146484 52284 146536 52290
rect 146484 52226 146536 52232
rect 146956 17406 146984 56782
rect 147048 19310 147076 57462
rect 147232 51074 147260 57598
rect 147324 52034 147352 60030
rect 147416 52222 147444 60044
rect 147706 60030 147904 60058
rect 147876 56778 147904 60030
rect 147680 56772 147732 56778
rect 147680 56714 147732 56720
rect 147864 56772 147916 56778
rect 147864 56714 147916 56720
rect 147404 52216 147456 52222
rect 147404 52158 147456 52164
rect 147324 52006 147628 52034
rect 147232 51046 147444 51074
rect 147416 48958 147444 51046
rect 147404 48952 147456 48958
rect 147404 48894 147456 48900
rect 147036 19304 147088 19310
rect 147036 19246 147088 19252
rect 147128 18624 147180 18630
rect 147128 18566 147180 18572
rect 146944 17400 146996 17406
rect 146944 17342 146996 17348
rect 146208 7132 146260 7138
rect 146208 7074 146260 7080
rect 144828 7064 144880 7070
rect 144828 7006 144880 7012
rect 147036 4616 147088 4622
rect 147036 4558 147088 4564
rect 144736 4140 144788 4146
rect 144736 4082 144788 4088
rect 144184 3936 144236 3942
rect 144184 3878 144236 3884
rect 144748 480 144776 4082
rect 145932 3868 145984 3874
rect 145932 3810 145984 3816
rect 145944 480 145972 3810
rect 147048 2394 147076 4558
rect 147140 3466 147168 18566
rect 147600 7274 147628 52006
rect 147692 51074 147720 56714
rect 147968 56642 147996 60044
rect 147956 56636 148008 56642
rect 147956 56578 148008 56584
rect 148244 52154 148272 60044
rect 148612 57662 148640 60044
rect 148600 57656 148652 57662
rect 148600 57598 148652 57604
rect 148324 56704 148376 56710
rect 148324 56646 148376 56652
rect 148232 52148 148284 52154
rect 148232 52090 148284 52096
rect 147692 51046 147996 51074
rect 147968 49434 147996 51046
rect 147956 49428 148008 49434
rect 147956 49370 148008 49376
rect 147588 7268 147640 7274
rect 147588 7210 147640 7216
rect 148336 4622 148364 56646
rect 148888 7410 148916 60044
rect 148968 56636 149020 56642
rect 148968 56578 149020 56584
rect 148876 7404 148928 7410
rect 148876 7346 148928 7352
rect 148980 7342 149008 56578
rect 149164 53786 149192 60044
rect 149440 57866 149468 60044
rect 149730 60030 150020 60058
rect 149428 57860 149480 57866
rect 149428 57802 149480 57808
rect 149152 53780 149204 53786
rect 149152 53722 149204 53728
rect 149992 51074 150020 60030
rect 150084 52086 150112 60044
rect 150360 57526 150388 60044
rect 150348 57520 150400 57526
rect 150348 57462 150400 57468
rect 150532 56840 150584 56846
rect 150532 56782 150584 56788
rect 150072 52080 150124 52086
rect 150072 52022 150124 52028
rect 150544 51074 150572 56782
rect 150636 56642 150664 60044
rect 150926 60030 151216 60058
rect 150900 56976 150952 56982
rect 150900 56918 150952 56924
rect 150624 56636 150676 56642
rect 150624 56578 150676 56584
rect 149992 51046 150388 51074
rect 150544 51046 150664 51074
rect 150360 7478 150388 51046
rect 150636 49706 150664 51046
rect 150912 50318 150940 56918
rect 151188 51074 151216 60030
rect 151280 56982 151308 60044
rect 151570 60030 151676 60058
rect 151268 56976 151320 56982
rect 151268 56918 151320 56924
rect 151188 51046 151584 51074
rect 150900 50312 150952 50318
rect 150900 50254 150952 50260
rect 150624 49700 150676 49706
rect 150624 49642 150676 49648
rect 151556 12578 151584 51046
rect 151544 12572 151596 12578
rect 151544 12514 151596 12520
rect 151648 8294 151676 60030
rect 151832 56710 151860 60044
rect 152108 57050 152136 60044
rect 152096 57044 152148 57050
rect 152096 56986 152148 56992
rect 151912 56908 151964 56914
rect 151912 56850 151964 56856
rect 151820 56704 151872 56710
rect 151820 56646 151872 56652
rect 151728 56636 151780 56642
rect 151728 56578 151780 56584
rect 151636 8288 151688 8294
rect 151636 8230 151688 8236
rect 151740 7546 151768 56578
rect 151924 51074 151952 56850
rect 152476 56642 152504 60044
rect 152766 60030 152964 60058
rect 152464 56636 152516 56642
rect 152464 56578 152516 56584
rect 152464 55888 152516 55894
rect 152464 55830 152516 55836
rect 151832 51046 151952 51074
rect 151832 49638 151860 51046
rect 151820 49632 151872 49638
rect 151820 49574 151872 49580
rect 151820 7744 151872 7750
rect 151820 7686 151872 7692
rect 151728 7540 151780 7546
rect 151728 7482 151780 7488
rect 150348 7472 150400 7478
rect 150348 7414 150400 7420
rect 148968 7336 149020 7342
rect 148968 7278 149020 7284
rect 150624 4752 150676 4758
rect 150624 4694 150676 4700
rect 148324 4616 148376 4622
rect 148324 4558 148376 4564
rect 148324 3800 148376 3806
rect 148324 3742 148376 3748
rect 147128 3460 147180 3466
rect 147128 3402 147180 3408
rect 147048 2366 147168 2394
rect 147140 480 147168 2366
rect 148336 480 148364 3742
rect 149520 3460 149572 3466
rect 149520 3402 149572 3408
rect 149532 480 149560 3402
rect 150636 480 150664 4694
rect 151832 480 151860 7686
rect 152476 3466 152504 55830
rect 152936 12714 152964 60030
rect 153028 56846 153056 60044
rect 153016 56840 153068 56846
rect 153016 56782 153068 56788
rect 153304 56778 153332 60044
rect 153686 60030 153884 60058
rect 153856 56794 153884 60030
rect 153948 56914 153976 60044
rect 154238 60030 154436 60058
rect 153936 56908 153988 56914
rect 153936 56850 153988 56856
rect 153292 56772 153344 56778
rect 153856 56766 154344 56794
rect 153292 56714 153344 56720
rect 153016 56704 153068 56710
rect 153016 56646 153068 56652
rect 154212 56704 154264 56710
rect 154212 56646 154264 56652
rect 152924 12708 152976 12714
rect 152924 12650 152976 12656
rect 153028 12646 153056 56646
rect 153108 56636 153160 56642
rect 153108 56578 153160 56584
rect 153016 12640 153068 12646
rect 153016 12582 153068 12588
rect 153120 8226 153148 56578
rect 154224 12850 154252 56646
rect 154212 12844 154264 12850
rect 154212 12786 154264 12792
rect 154316 12782 154344 56766
rect 154304 12776 154356 12782
rect 154304 12718 154356 12724
rect 153108 8220 153160 8226
rect 153108 8162 153160 8168
rect 154408 8090 154436 60030
rect 154500 56710 154528 60044
rect 154488 56704 154540 56710
rect 154488 56646 154540 56652
rect 154488 56568 154540 56574
rect 154488 56510 154540 56516
rect 154500 8158 154528 56510
rect 154868 49162 154896 60044
rect 155158 60030 155356 60058
rect 155434 60030 155632 60058
rect 155710 60030 155908 60058
rect 155224 56840 155276 56846
rect 155224 56782 155276 56788
rect 154856 49156 154908 49162
rect 154856 49098 154908 49104
rect 155236 18698 155264 56782
rect 155328 51074 155356 60030
rect 155500 57384 155552 57390
rect 155500 57326 155552 57332
rect 155512 53990 155540 57326
rect 155604 55570 155632 60030
rect 155604 55542 155816 55570
rect 155500 53984 155552 53990
rect 155500 53926 155552 53932
rect 155328 51046 155632 51074
rect 155224 18692 155276 18698
rect 155224 18634 155276 18640
rect 154488 8152 154540 8158
rect 154488 8094 154540 8100
rect 154396 8084 154448 8090
rect 154396 8026 154448 8032
rect 155604 8022 155632 51046
rect 155788 12918 155816 55542
rect 155880 54126 155908 60030
rect 156064 57526 156092 60044
rect 156052 57520 156104 57526
rect 156052 57462 156104 57468
rect 156340 56642 156368 60044
rect 156616 56914 156644 60044
rect 156892 57458 156920 60044
rect 157076 60030 157182 60058
rect 156880 57452 156932 57458
rect 156880 57394 156932 57400
rect 156604 56908 156656 56914
rect 156604 56850 156656 56856
rect 156328 56636 156380 56642
rect 156328 56578 156380 56584
rect 156972 56636 157024 56642
rect 156972 56578 157024 56584
rect 155868 54120 155920 54126
rect 155868 54062 155920 54068
rect 155868 53984 155920 53990
rect 155868 53926 155920 53932
rect 155880 49502 155908 53926
rect 155868 49496 155920 49502
rect 155868 49438 155920 49444
rect 156984 12986 157012 56578
rect 157076 13054 157104 60030
rect 157536 57662 157564 60044
rect 157524 57656 157576 57662
rect 157524 57598 157576 57604
rect 157156 57520 157208 57526
rect 157156 57462 157208 57468
rect 157064 13048 157116 13054
rect 157064 12990 157116 12996
rect 156972 12980 157024 12986
rect 156972 12922 157024 12928
rect 155776 12912 155828 12918
rect 155776 12854 155828 12860
rect 155592 8016 155644 8022
rect 155592 7958 155644 7964
rect 157168 7954 157196 57462
rect 157248 57452 157300 57458
rect 157248 57394 157300 57400
rect 157156 7948 157208 7954
rect 157156 7890 157208 7896
rect 157260 7886 157288 57394
rect 157708 56908 157760 56914
rect 157708 56850 157760 56856
rect 157720 51074 157748 56850
rect 157812 56710 157840 60044
rect 157800 56704 157852 56710
rect 157800 56646 157852 56652
rect 158088 56642 158116 60044
rect 158378 60030 158484 60058
rect 158746 60030 158944 60058
rect 158076 56636 158128 56642
rect 158076 56578 158128 56584
rect 157720 51046 157840 51074
rect 157812 49094 157840 51046
rect 157800 49088 157852 49094
rect 157800 49030 157852 49036
rect 158456 48006 158484 60030
rect 158916 56710 158944 60030
rect 159008 56778 159036 60044
rect 159100 60030 159298 60058
rect 158996 56772 159048 56778
rect 158996 56714 159048 56720
rect 158628 56704 158680 56710
rect 158628 56646 158680 56652
rect 158904 56704 158956 56710
rect 158904 56646 158956 56652
rect 158536 56636 158588 56642
rect 158536 56578 158588 56584
rect 158444 48000 158496 48006
rect 158444 47942 158496 47948
rect 158548 13802 158576 56578
rect 158536 13796 158588 13802
rect 158536 13738 158588 13744
rect 157248 7880 157300 7886
rect 157248 7822 157300 7828
rect 158640 7818 158668 56646
rect 159100 51066 159128 60030
rect 159560 56642 159588 60044
rect 159744 60030 159942 60058
rect 160218 60030 160416 60058
rect 159640 56704 159692 56710
rect 159640 56646 159692 56652
rect 159548 56636 159600 56642
rect 159548 56578 159600 56584
rect 159088 51060 159140 51066
rect 159088 51002 159140 51008
rect 158628 7812 158680 7818
rect 158628 7754 158680 7760
rect 159652 7750 159680 56646
rect 159744 13666 159772 60030
rect 159824 56772 159876 56778
rect 159824 56714 159876 56720
rect 159836 13734 159864 56714
rect 159916 56636 159968 56642
rect 159916 56578 159968 56584
rect 159824 13728 159876 13734
rect 159824 13670 159876 13676
rect 159732 13660 159784 13666
rect 159732 13602 159784 13608
rect 159640 7744 159692 7750
rect 159640 7686 159692 7692
rect 159928 7682 159956 56578
rect 160388 49026 160416 60030
rect 160480 56710 160508 60044
rect 160468 56704 160520 56710
rect 160468 56646 160520 56652
rect 160756 56642 160784 60044
rect 160744 56636 160796 56642
rect 160744 56578 160796 56584
rect 160376 49020 160428 49026
rect 160376 48962 160428 48968
rect 161124 47870 161152 60044
rect 161216 60030 161414 60058
rect 161112 47864 161164 47870
rect 161112 47806 161164 47812
rect 161216 18630 161244 60030
rect 161572 57860 161624 57866
rect 161572 57802 161624 57808
rect 161388 56704 161440 56710
rect 161388 56646 161440 56652
rect 161296 56636 161348 56642
rect 161296 56578 161348 56584
rect 161204 18624 161256 18630
rect 161204 18566 161256 18572
rect 161308 13598 161336 56578
rect 161296 13592 161348 13598
rect 161296 13534 161348 13540
rect 155408 7676 155460 7682
rect 155408 7618 155460 7624
rect 159916 7676 159968 7682
rect 159916 7618 159968 7624
rect 154212 5500 154264 5506
rect 154212 5442 154264 5448
rect 153016 3528 153068 3534
rect 153016 3470 153068 3476
rect 152464 3460 152516 3466
rect 152464 3402 152516 3408
rect 153028 480 153056 3470
rect 154224 480 154252 5442
rect 155420 480 155448 7618
rect 161400 7614 161428 56646
rect 161584 49298 161612 57802
rect 161676 56642 161704 60044
rect 161952 57866 161980 60044
rect 161940 57860 161992 57866
rect 161940 57802 161992 57808
rect 162124 57724 162176 57730
rect 162124 57666 162176 57672
rect 161664 56636 161716 56642
rect 161664 56578 161716 56584
rect 161572 49292 161624 49298
rect 161572 49234 161624 49240
rect 162136 19106 162164 57666
rect 162320 54942 162348 60044
rect 162610 60030 162716 60058
rect 162584 56636 162636 56642
rect 162584 56578 162636 56584
rect 162308 54936 162360 54942
rect 162308 54878 162360 54884
rect 162124 19100 162176 19106
rect 162124 19042 162176 19048
rect 162596 13530 162624 56578
rect 162584 13524 162636 13530
rect 162584 13466 162636 13472
rect 162688 13462 162716 60030
rect 162872 56642 162900 60044
rect 162860 56636 162912 56642
rect 162860 56578 162912 56584
rect 163148 55758 163176 60044
rect 163438 60030 163728 60058
rect 163136 55752 163188 55758
rect 163136 55694 163188 55700
rect 163700 51074 163728 60030
rect 163792 57254 163820 60044
rect 164082 60030 164188 60058
rect 163780 57248 163832 57254
rect 163780 57190 163832 57196
rect 164056 56636 164108 56642
rect 164056 56578 164108 56584
rect 163700 51046 164004 51074
rect 162676 13456 162728 13462
rect 162676 13398 162728 13404
rect 163976 13394 164004 51046
rect 164068 47802 164096 56578
rect 164160 54874 164188 60030
rect 164344 56642 164372 60044
rect 164620 57798 164648 60044
rect 164608 57792 164660 57798
rect 164608 57734 164660 57740
rect 164332 56636 164384 56642
rect 164332 56578 164384 56584
rect 164148 54868 164200 54874
rect 164148 54810 164200 54816
rect 164988 54806 165016 60044
rect 165264 56642 165292 60044
rect 165356 60030 165554 60058
rect 165160 56636 165212 56642
rect 165160 56578 165212 56584
rect 165252 56636 165304 56642
rect 165252 56578 165304 56584
rect 164976 54800 165028 54806
rect 164976 54742 165028 54748
rect 165172 51074 165200 56578
rect 165172 51046 165292 51074
rect 164056 47796 164108 47802
rect 164056 47738 164108 47744
rect 163964 13388 164016 13394
rect 163964 13330 164016 13336
rect 165264 13326 165292 51046
rect 165356 47598 165384 60030
rect 165436 56636 165488 56642
rect 165436 56578 165488 56584
rect 165344 47592 165396 47598
rect 165344 47534 165396 47540
rect 165252 13320 165304 13326
rect 165252 13262 165304 13268
rect 165448 13258 165476 56578
rect 165816 53718 165844 60044
rect 166184 56642 166212 60044
rect 166460 57730 166488 60044
rect 166264 57724 166316 57730
rect 166264 57666 166316 57672
rect 166448 57724 166500 57730
rect 166448 57666 166500 57672
rect 166172 56636 166224 56642
rect 166172 56578 166224 56584
rect 165804 53712 165856 53718
rect 165804 53654 165856 53660
rect 166276 17610 166304 57666
rect 166356 56704 166408 56710
rect 166356 56646 166408 56652
rect 166368 18834 166396 56646
rect 166736 53650 166764 60044
rect 167012 57662 167040 60044
rect 167000 57656 167052 57662
rect 167000 57598 167052 57604
rect 167380 57594 167408 60044
rect 167368 57588 167420 57594
rect 167368 57530 167420 57536
rect 166908 56636 166960 56642
rect 166908 56578 166960 56584
rect 166724 53644 166776 53650
rect 166724 53586 166776 53592
rect 166356 18828 166408 18834
rect 166356 18770 166408 18776
rect 166264 17604 166316 17610
rect 166264 17546 166316 17552
rect 165436 13252 165488 13258
rect 165436 13194 165488 13200
rect 166920 13190 166948 56578
rect 167656 55826 167684 60044
rect 167748 60030 167946 60058
rect 168116 60030 168222 60058
rect 168392 60030 168590 60058
rect 168760 60030 168866 60058
rect 167644 55820 167696 55826
rect 167644 55762 167696 55768
rect 167748 54738 167776 60030
rect 167736 54732 167788 54738
rect 167736 54674 167788 54680
rect 166908 13184 166960 13190
rect 166908 13126 166960 13132
rect 163688 9580 163740 9586
rect 163688 9522 163740 9528
rect 158904 7608 158956 7614
rect 158904 7550 158956 7556
rect 161388 7608 161440 7614
rect 161388 7550 161440 7556
rect 157800 5432 157852 5438
rect 157800 5374 157852 5380
rect 156604 3460 156656 3466
rect 156604 3402 156656 3408
rect 156616 480 156644 3402
rect 157812 480 157840 5374
rect 158916 480 158944 7550
rect 162492 5364 162544 5370
rect 162492 5306 162544 5312
rect 161296 3936 161348 3942
rect 161296 3878 161348 3884
rect 160100 3392 160152 3398
rect 160100 3334 160152 3340
rect 160112 480 160140 3334
rect 161308 480 161336 3878
rect 162504 480 162532 5306
rect 163700 480 163728 9522
rect 167184 9512 167236 9518
rect 167184 9454 167236 9460
rect 166080 5296 166132 5302
rect 166080 5238 166132 5244
rect 164884 3664 164936 3670
rect 164884 3606 164936 3612
rect 164896 480 164924 3606
rect 166092 480 166120 5238
rect 167196 480 167224 9454
rect 168116 4010 168144 60030
rect 168196 57656 168248 57662
rect 168196 57598 168248 57604
rect 168208 13122 168236 57598
rect 168392 53514 168420 60030
rect 168380 53508 168432 53514
rect 168380 53450 168432 53456
rect 168760 52018 168788 60030
rect 169128 57118 169156 60044
rect 169418 60030 169708 60058
rect 169786 60030 169984 60058
rect 169116 57112 169168 57118
rect 169116 57054 169168 57060
rect 169024 56840 169076 56846
rect 169024 56782 169076 56788
rect 168748 52012 168800 52018
rect 168748 51954 168800 51960
rect 169036 18970 169064 56782
rect 169116 56636 169168 56642
rect 169116 56578 169168 56584
rect 169128 19038 169156 56578
rect 169116 19032 169168 19038
rect 169116 18974 169168 18980
rect 169024 18964 169076 18970
rect 169024 18906 169076 18912
rect 168196 13116 168248 13122
rect 168196 13058 168248 13064
rect 169680 8430 169708 60030
rect 169956 51950 169984 60030
rect 170048 56982 170076 60044
rect 170324 57866 170352 60044
rect 170416 60030 170614 60058
rect 170312 57860 170364 57866
rect 170312 57802 170364 57808
rect 170416 57644 170444 60030
rect 170876 57798 170904 60044
rect 170956 57860 171008 57866
rect 170956 57802 171008 57808
rect 170864 57792 170916 57798
rect 170864 57734 170916 57740
rect 170324 57616 170444 57644
rect 170036 56976 170088 56982
rect 170036 56918 170088 56924
rect 169944 51944 169996 51950
rect 169944 51886 169996 51892
rect 170324 50998 170352 57616
rect 170496 56772 170548 56778
rect 170496 56714 170548 56720
rect 170404 56704 170456 56710
rect 170404 56646 170456 56652
rect 170312 50992 170364 50998
rect 170312 50934 170364 50940
rect 170416 17542 170444 56646
rect 170508 18902 170536 56714
rect 170968 55214 170996 57802
rect 171244 57322 171272 60044
rect 171232 57316 171284 57322
rect 171232 57258 171284 57264
rect 171324 57248 171376 57254
rect 171324 57190 171376 57196
rect 170968 55186 171088 55214
rect 170496 18896 170548 18902
rect 170496 18838 170548 18844
rect 170404 17536 170456 17542
rect 170404 17478 170456 17484
rect 170772 9444 170824 9450
rect 170772 9386 170824 9392
rect 169668 8424 169720 8430
rect 169668 8366 169720 8372
rect 169576 5228 169628 5234
rect 169576 5170 169628 5176
rect 168104 4004 168156 4010
rect 168104 3946 168156 3952
rect 168380 3596 168432 3602
rect 168380 3538 168432 3544
rect 168392 480 168420 3538
rect 169588 480 169616 5170
rect 170784 480 170812 9386
rect 171060 8498 171088 55186
rect 171336 53378 171364 57190
rect 171520 56574 171548 60044
rect 171810 60030 172008 60058
rect 172086 60030 172376 60058
rect 171508 56568 171560 56574
rect 171508 56510 171560 56516
rect 171980 55214 172008 60030
rect 172244 57316 172296 57322
rect 172244 57258 172296 57264
rect 171980 55186 172192 55214
rect 171324 53372 171376 53378
rect 171324 53314 171376 53320
rect 171048 8492 171100 8498
rect 171048 8434 171100 8440
rect 172164 3874 172192 55186
rect 172256 8566 172284 57258
rect 172348 8634 172376 60030
rect 172440 57254 172468 60044
rect 172428 57248 172480 57254
rect 172428 57190 172480 57196
rect 172716 57050 172744 60044
rect 172520 57044 172572 57050
rect 172520 56986 172572 56992
rect 172704 57044 172756 57050
rect 172704 56986 172756 56992
rect 172532 49366 172560 56986
rect 172992 56710 173020 60044
rect 173084 60030 173282 60058
rect 172980 56704 173032 56710
rect 172980 56646 173032 56652
rect 173084 50930 173112 60030
rect 173636 57186 173664 60044
rect 173912 57254 173940 60044
rect 174096 60030 174202 60058
rect 174478 60030 174676 60058
rect 173992 57316 174044 57322
rect 173992 57258 174044 57264
rect 173900 57248 173952 57254
rect 173900 57190 173952 57196
rect 173164 57180 173216 57186
rect 173164 57122 173216 57128
rect 173624 57180 173676 57186
rect 173624 57122 173676 57128
rect 173072 50924 173124 50930
rect 173072 50866 173124 50872
rect 172520 49360 172572 49366
rect 172520 49302 172572 49308
rect 173176 18766 173204 57122
rect 173256 56840 173308 56846
rect 173256 56782 173308 56788
rect 173268 19174 173296 56782
rect 173808 56704 173860 56710
rect 173808 56646 173860 56652
rect 173256 19168 173308 19174
rect 173256 19110 173308 19116
rect 173164 18760 173216 18766
rect 173164 18702 173216 18708
rect 173820 8702 173848 56646
rect 174004 50862 174032 57258
rect 174096 51882 174124 60030
rect 174648 56982 174676 60030
rect 174544 56976 174596 56982
rect 174544 56918 174596 56924
rect 174636 56976 174688 56982
rect 174636 56918 174688 56924
rect 174084 51876 174136 51882
rect 174084 51818 174136 51824
rect 173992 50856 174044 50862
rect 173992 50798 174044 50804
rect 174268 9376 174320 9382
rect 174268 9318 174320 9324
rect 173808 8696 173860 8702
rect 173808 8638 173860 8644
rect 172336 8628 172388 8634
rect 172336 8570 172388 8576
rect 172244 8560 172296 8566
rect 172244 8502 172296 8508
rect 173164 5160 173216 5166
rect 173164 5102 173216 5108
rect 172152 3868 172204 3874
rect 172152 3810 172204 3816
rect 171968 3732 172020 3738
rect 171968 3674 172020 3680
rect 171980 480 172008 3674
rect 173176 480 173204 5102
rect 174280 480 174308 9318
rect 174556 3942 174584 56918
rect 174832 56846 174860 60044
rect 174924 60030 175122 60058
rect 174924 57322 174952 60030
rect 175384 57322 175412 60044
rect 174912 57316 174964 57322
rect 174912 57258 174964 57264
rect 175372 57316 175424 57322
rect 175372 57258 175424 57264
rect 175096 57248 175148 57254
rect 175096 57190 175148 57196
rect 174820 56840 174872 56846
rect 174820 56782 174872 56788
rect 175108 8770 175136 57190
rect 175188 56840 175240 56846
rect 175188 56782 175240 56788
rect 175200 8838 175228 56782
rect 175660 56778 175688 60044
rect 176042 60030 176240 60058
rect 175924 57180 175976 57186
rect 175924 57122 175976 57128
rect 175648 56772 175700 56778
rect 175648 56714 175700 56720
rect 175188 8832 175240 8838
rect 175188 8774 175240 8780
rect 175096 8764 175148 8770
rect 175096 8706 175148 8712
rect 175464 4616 175516 4622
rect 175464 4558 175516 4564
rect 174544 3936 174596 3942
rect 174544 3878 174596 3884
rect 175476 480 175504 4558
rect 175936 3806 175964 57122
rect 176212 55214 176240 60030
rect 176304 57186 176332 60044
rect 176396 60030 176594 60058
rect 176292 57180 176344 57186
rect 176292 57122 176344 57128
rect 176212 55186 176332 55214
rect 176304 13938 176332 55186
rect 176292 13932 176344 13938
rect 176292 13874 176344 13880
rect 176396 9654 176424 60030
rect 176856 57322 176884 60044
rect 176568 57316 176620 57322
rect 176568 57258 176620 57264
rect 176844 57316 176896 57322
rect 176844 57258 176896 57264
rect 176476 56772 176528 56778
rect 176476 56714 176528 56720
rect 176384 9648 176436 9654
rect 176384 9590 176436 9596
rect 176488 8906 176516 56714
rect 176476 8900 176528 8906
rect 176476 8842 176528 8848
rect 175924 3800 175976 3806
rect 175924 3742 175976 3748
rect 176580 3738 176608 57258
rect 177132 57186 177160 60044
rect 177500 57254 177528 60044
rect 177672 57316 177724 57322
rect 177672 57258 177724 57264
rect 177488 57248 177540 57254
rect 177488 57190 177540 57196
rect 177120 57180 177172 57186
rect 177120 57122 177172 57128
rect 177684 14006 177712 57258
rect 177776 14074 177804 60044
rect 177856 57248 177908 57254
rect 177856 57190 177908 57196
rect 177764 14068 177816 14074
rect 177764 14010 177816 14016
rect 177672 14000 177724 14006
rect 177672 13942 177724 13948
rect 177868 9586 177896 57190
rect 177948 57180 178000 57186
rect 177948 57122 178000 57128
rect 177856 9580 177908 9586
rect 177856 9522 177908 9528
rect 177856 9308 177908 9314
rect 177856 9250 177908 9256
rect 176660 9240 176712 9246
rect 176660 9182 176712 9188
rect 176568 3732 176620 3738
rect 176568 3674 176620 3680
rect 176672 480 176700 9182
rect 177868 480 177896 9250
rect 177960 3670 177988 57122
rect 178052 57050 178080 60044
rect 178328 57254 178356 60044
rect 178710 60030 178908 60058
rect 178316 57248 178368 57254
rect 178316 57190 178368 57196
rect 178040 57044 178092 57050
rect 178040 56986 178092 56992
rect 178880 55214 178908 60030
rect 178972 57322 179000 60044
rect 179156 60030 179262 60058
rect 179538 60030 179828 60058
rect 178960 57316 179012 57322
rect 178960 57258 179012 57264
rect 178880 55186 179092 55214
rect 179064 14142 179092 55186
rect 179052 14136 179104 14142
rect 179052 14078 179104 14084
rect 179156 9450 179184 60030
rect 179328 57316 179380 57322
rect 179328 57258 179380 57264
rect 179236 57248 179288 57254
rect 179236 57190 179288 57196
rect 179248 9518 179276 57190
rect 179236 9512 179288 9518
rect 179236 9454 179288 9460
rect 179144 9444 179196 9450
rect 179144 9386 179196 9392
rect 179052 4480 179104 4486
rect 179052 4422 179104 4428
rect 177948 3664 178000 3670
rect 177948 3606 178000 3612
rect 179064 480 179092 4422
rect 179340 3602 179368 57258
rect 179800 56710 179828 60030
rect 179892 57254 179920 60044
rect 179880 57248 179932 57254
rect 179880 57190 179932 57196
rect 180168 56846 180196 60044
rect 180458 60030 180564 60058
rect 180156 56840 180208 56846
rect 180156 56782 180208 56788
rect 179788 56704 179840 56710
rect 179788 56646 179840 56652
rect 179512 56636 179564 56642
rect 179512 56578 179564 56584
rect 179524 47938 179552 56578
rect 179512 47932 179564 47938
rect 179512 47874 179564 47880
rect 180536 14278 180564 60030
rect 180720 57254 180748 60044
rect 180708 57248 180760 57254
rect 180708 57190 180760 57196
rect 180708 56840 180760 56846
rect 180708 56782 180760 56788
rect 180616 56704 180668 56710
rect 180616 56646 180668 56652
rect 180524 14272 180576 14278
rect 180524 14214 180576 14220
rect 180628 14210 180656 56646
rect 180616 14204 180668 14210
rect 180616 14146 180668 14152
rect 180720 9382 180748 56782
rect 181088 56506 181116 60044
rect 181378 60030 181576 60058
rect 181654 60030 181852 60058
rect 181930 60030 182128 60058
rect 181076 56500 181128 56506
rect 181076 56442 181128 56448
rect 181548 55214 181576 60030
rect 181824 57610 181852 60030
rect 181824 57582 182036 57610
rect 181548 55186 181944 55214
rect 180708 9376 180760 9382
rect 180708 9318 180760 9324
rect 181916 9314 181944 55186
rect 182008 14346 182036 57582
rect 182100 56098 182128 60030
rect 182284 56914 182312 60044
rect 182560 57390 182588 60044
rect 182548 57384 182600 57390
rect 182548 57326 182600 57332
rect 182272 56908 182324 56914
rect 182272 56850 182324 56856
rect 182836 56370 182864 60044
rect 182824 56364 182876 56370
rect 182824 56306 182876 56312
rect 182088 56092 182140 56098
rect 182088 56034 182140 56040
rect 182548 14476 182600 14482
rect 182548 14418 182600 14424
rect 181996 14340 182048 14346
rect 181996 14282 182048 14288
rect 181904 9308 181956 9314
rect 181904 9250 181956 9256
rect 180248 9172 180300 9178
rect 180248 9114 180300 9120
rect 179328 3596 179380 3602
rect 179328 3538 179380 3544
rect 180260 480 180288 9114
rect 181444 9104 181496 9110
rect 181444 9046 181496 9052
rect 181456 480 181484 9046
rect 182560 480 182588 14418
rect 183112 9178 183140 60044
rect 183204 60030 183494 60058
rect 183204 15162 183232 60030
rect 183284 57384 183336 57390
rect 183284 57326 183336 57332
rect 183192 15156 183244 15162
rect 183192 15098 183244 15104
rect 183296 14414 183324 57326
rect 183376 56908 183428 56914
rect 183376 56850 183428 56856
rect 183284 14408 183336 14414
rect 183284 14350 183336 14356
rect 183388 9246 183416 56850
rect 183756 56438 183784 60044
rect 184032 57390 184060 60044
rect 184322 60030 184520 60058
rect 184598 60030 184888 60058
rect 184492 57610 184520 60030
rect 184492 57582 184796 57610
rect 184020 57384 184072 57390
rect 184020 57326 184072 57332
rect 184664 57384 184716 57390
rect 184664 57326 184716 57332
rect 184204 56840 184256 56846
rect 184204 56782 184256 56788
rect 183744 56432 183796 56438
rect 183744 56374 183796 56380
rect 184216 20126 184244 56782
rect 184204 20120 184256 20126
rect 184204 20062 184256 20068
rect 183376 9240 183428 9246
rect 183376 9182 183428 9188
rect 183100 9172 183152 9178
rect 183100 9114 183152 9120
rect 184676 9110 184704 57326
rect 184768 15094 184796 57582
rect 184860 56302 184888 60030
rect 184952 57390 184980 60044
rect 184940 57384 184992 57390
rect 184940 57326 184992 57332
rect 185228 56642 185256 60044
rect 185216 56636 185268 56642
rect 185216 56578 185268 56584
rect 184848 56296 184900 56302
rect 184848 56238 184900 56244
rect 185504 56234 185532 60044
rect 185780 56982 185808 60044
rect 186056 60030 186162 60058
rect 186438 60030 186636 60058
rect 185860 57384 185912 57390
rect 185860 57326 185912 57332
rect 185768 56976 185820 56982
rect 185768 56918 185820 56924
rect 185492 56228 185544 56234
rect 185492 56170 185544 56176
rect 184756 15088 184808 15094
rect 184756 15030 184808 15036
rect 184664 9104 184716 9110
rect 184664 9046 184716 9052
rect 185872 9042 185900 57326
rect 185952 56636 186004 56642
rect 185952 56578 186004 56584
rect 185964 15026 185992 56578
rect 185952 15020 186004 15026
rect 185952 14962 186004 14968
rect 186056 14958 186084 60030
rect 186504 57384 186556 57390
rect 186504 57326 186556 57332
rect 186136 56976 186188 56982
rect 186136 56918 186188 56924
rect 186320 56976 186372 56982
rect 186320 56918 186372 56924
rect 186044 14952 186096 14958
rect 186044 14894 186096 14900
rect 183744 9036 183796 9042
rect 183744 8978 183796 8984
rect 185860 9036 185912 9042
rect 185860 8978 185912 8984
rect 183756 480 183784 8978
rect 186148 8974 186176 56918
rect 186332 53310 186360 56918
rect 186516 53446 186544 57326
rect 186608 56030 186636 60030
rect 186700 56982 186728 60044
rect 186990 60030 187280 60058
rect 186688 56976 186740 56982
rect 186688 56918 186740 56924
rect 186964 56704 187016 56710
rect 186964 56646 187016 56652
rect 186596 56024 186648 56030
rect 186596 55966 186648 55972
rect 186504 53440 186556 53446
rect 186504 53382 186556 53388
rect 186320 53304 186372 53310
rect 186320 53246 186372 53252
rect 186976 20262 187004 56646
rect 187252 55214 187280 60030
rect 187344 56166 187372 60044
rect 187620 57390 187648 60044
rect 187608 57384 187660 57390
rect 187608 57326 187660 57332
rect 187792 57384 187844 57390
rect 187792 57326 187844 57332
rect 187332 56160 187384 56166
rect 187332 56102 187384 56108
rect 187252 55186 187372 55214
rect 186964 20256 187016 20262
rect 186964 20198 187016 20204
rect 187344 14890 187372 55186
rect 187804 53582 187832 57326
rect 187896 56982 187924 60044
rect 187988 60030 188186 60058
rect 187884 56976 187936 56982
rect 187884 56918 187936 56924
rect 187988 54602 188016 60030
rect 188540 57390 188568 60044
rect 188724 60030 188830 60058
rect 188528 57384 188580 57390
rect 188528 57326 188580 57332
rect 188344 56772 188396 56778
rect 188344 56714 188396 56720
rect 187976 54596 188028 54602
rect 187976 54538 188028 54544
rect 187792 53576 187844 53582
rect 187792 53518 187844 53524
rect 188356 47734 188384 56714
rect 188344 47728 188396 47734
rect 188344 47670 188396 47676
rect 187332 14884 187384 14890
rect 187332 14826 187384 14832
rect 188724 14754 188752 60030
rect 189092 57390 189120 60044
rect 189080 57384 189132 57390
rect 189080 57326 189132 57332
rect 188896 56976 188948 56982
rect 188896 56918 188948 56924
rect 188908 14822 188936 56918
rect 189368 55894 189396 60044
rect 189750 60030 189948 60058
rect 190026 60030 190224 60058
rect 190302 60030 190408 60058
rect 189920 57610 189948 60030
rect 190196 57746 190224 60030
rect 190196 57718 190316 57746
rect 189920 57582 190224 57610
rect 190092 57384 190144 57390
rect 190092 57326 190144 57332
rect 189540 56840 189592 56846
rect 189540 56782 189592 56788
rect 189356 55888 189408 55894
rect 189356 55830 189408 55836
rect 189552 54670 189580 56782
rect 189540 54664 189592 54670
rect 189540 54606 189592 54612
rect 188896 14816 188948 14822
rect 188896 14758 188948 14764
rect 188712 14748 188764 14754
rect 188712 14690 188764 14696
rect 187332 11008 187384 11014
rect 187332 10950 187384 10956
rect 184940 8968 184992 8974
rect 184940 8910 184992 8916
rect 186136 8968 186188 8974
rect 186136 8910 186188 8916
rect 184952 480 184980 8910
rect 186136 4684 186188 4690
rect 186136 4626 186188 4632
rect 186148 480 186176 4626
rect 187344 480 187372 10950
rect 188528 10940 188580 10946
rect 188528 10882 188580 10888
rect 188540 480 188568 10882
rect 189724 5092 189776 5098
rect 189724 5034 189776 5040
rect 189736 480 189764 5034
rect 190104 4282 190132 57326
rect 190196 14686 190224 57582
rect 190184 14680 190236 14686
rect 190184 14622 190236 14628
rect 190288 4350 190316 57718
rect 190380 56846 190408 60030
rect 190564 57390 190592 60044
rect 190552 57384 190604 57390
rect 190552 57326 190604 57332
rect 190840 56846 190868 60044
rect 190932 60030 191222 60058
rect 190368 56840 190420 56846
rect 190368 56782 190420 56788
rect 190828 56840 190880 56846
rect 190828 56782 190880 56788
rect 190932 53174 190960 60030
rect 191380 56840 191432 56846
rect 191380 56782 191432 56788
rect 190920 53168 190972 53174
rect 190920 53110 190972 53116
rect 190828 10872 190880 10878
rect 190828 10814 190880 10820
rect 190276 4344 190328 4350
rect 190276 4286 190328 4292
rect 190092 4276 190144 4282
rect 190092 4218 190144 4224
rect 190840 480 190868 10814
rect 191392 4418 191420 56782
rect 191484 14550 191512 60044
rect 191668 60030 191774 60058
rect 191944 60030 192050 60058
rect 191564 57384 191616 57390
rect 191564 57326 191616 57332
rect 191576 14618 191604 57326
rect 191564 14612 191616 14618
rect 191564 14554 191616 14560
rect 191472 14544 191524 14550
rect 191472 14486 191524 14492
rect 191668 4486 191696 60030
rect 191944 53242 191972 60030
rect 192404 57390 192432 60044
rect 192694 60030 192892 60058
rect 192392 57384 192444 57390
rect 192392 57326 192444 57332
rect 192116 56908 192168 56914
rect 192116 56850 192168 56856
rect 191932 53236 191984 53242
rect 191932 53178 191984 53184
rect 192128 53106 192156 56850
rect 192116 53100 192168 53106
rect 192116 53042 192168 53048
rect 192024 10804 192076 10810
rect 192024 10746 192076 10752
rect 191656 4480 191708 4486
rect 191656 4422 191708 4428
rect 191380 4412 191432 4418
rect 191380 4354 191432 4360
rect 192036 480 192064 10746
rect 192864 4554 192892 60030
rect 192956 56914 192984 60044
rect 193232 57390 193260 60044
rect 193324 60030 193614 60058
rect 193692 60030 193890 60058
rect 193036 57384 193088 57390
rect 193036 57326 193088 57332
rect 193220 57384 193272 57390
rect 193220 57326 193272 57332
rect 192944 56908 192996 56914
rect 192944 56850 192996 56856
rect 193048 14482 193076 57326
rect 193324 56846 193352 60030
rect 193692 57610 193720 60030
rect 193416 57582 193720 57610
rect 193312 56840 193364 56846
rect 193312 56782 193364 56788
rect 193416 54534 193444 57582
rect 193680 57384 193732 57390
rect 193680 57326 193732 57332
rect 193496 56908 193548 56914
rect 193496 56850 193548 56856
rect 193404 54528 193456 54534
rect 193404 54470 193456 54476
rect 193508 50794 193536 56850
rect 193692 51814 193720 57326
rect 194152 56914 194180 60044
rect 194244 60030 194442 60058
rect 194140 56908 194192 56914
rect 194140 56850 194192 56856
rect 193680 51808 193732 51814
rect 193680 51750 193732 51756
rect 193496 50788 193548 50794
rect 193496 50730 193548 50736
rect 194244 45554 194272 60030
rect 194796 56914 194824 60044
rect 194888 60030 195086 60058
rect 194784 56908 194836 56914
rect 194784 56850 194836 56856
rect 194416 56840 194468 56846
rect 194416 56782 194468 56788
rect 194152 45526 194272 45554
rect 193036 14476 193088 14482
rect 193036 14418 193088 14424
rect 193220 10668 193272 10674
rect 193220 10610 193272 10616
rect 192852 4548 192904 4554
rect 192852 4490 192904 4496
rect 193232 3534 193260 10610
rect 194152 5030 194180 45526
rect 194428 16574 194456 56782
rect 194888 50590 194916 60030
rect 195348 57390 195376 60044
rect 195638 60030 195836 60058
rect 196006 60030 196204 60058
rect 195336 57384 195388 57390
rect 195336 57326 195388 57332
rect 195704 56908 195756 56914
rect 195704 56850 195756 56856
rect 194876 50584 194928 50590
rect 194876 50526 194928 50532
rect 194428 16546 194548 16574
rect 193312 5024 193364 5030
rect 193312 4966 193364 4972
rect 194140 5024 194192 5030
rect 194140 4966 194192 4972
rect 193220 3528 193272 3534
rect 193220 3470 193272 3476
rect 193324 2530 193352 4966
rect 194520 4622 194548 16546
rect 195612 10736 195664 10742
rect 195612 10678 195664 10684
rect 194508 4616 194560 4622
rect 194508 4558 194560 4564
rect 194416 3528 194468 3534
rect 194416 3470 194468 3476
rect 193232 2502 193352 2530
rect 193232 480 193260 2502
rect 194428 480 194456 3470
rect 195624 480 195652 10678
rect 195716 10198 195744 56850
rect 195808 10266 195836 60030
rect 195888 57384 195940 57390
rect 195888 57326 195940 57332
rect 195796 10260 195848 10266
rect 195796 10202 195848 10208
rect 195704 10192 195756 10198
rect 195704 10134 195756 10140
rect 195900 4690 195928 57326
rect 196176 50522 196204 60030
rect 196268 56914 196296 60044
rect 196544 57390 196572 60044
rect 196636 60030 196834 60058
rect 196532 57384 196584 57390
rect 196532 57326 196584 57332
rect 196256 56908 196308 56914
rect 196256 56850 196308 56856
rect 196164 50516 196216 50522
rect 196164 50458 196216 50464
rect 196636 50454 196664 60030
rect 197084 57384 197136 57390
rect 197084 57326 197136 57332
rect 196900 56908 196952 56914
rect 196900 56850 196952 56856
rect 196624 50448 196676 50454
rect 196624 50390 196676 50396
rect 196912 5506 196940 56850
rect 197096 11014 197124 57326
rect 197084 11008 197136 11014
rect 197084 10950 197136 10956
rect 196900 5500 196952 5506
rect 196900 5442 196952 5448
rect 197188 5438 197216 60044
rect 197464 57390 197492 60044
rect 197452 57384 197504 57390
rect 197452 57326 197504 57332
rect 197636 56908 197688 56914
rect 197636 56850 197688 56856
rect 197648 50726 197676 56850
rect 197636 50720 197688 50726
rect 197636 50662 197688 50668
rect 197740 50386 197768 60044
rect 198030 60030 198228 60058
rect 198306 60030 198596 60058
rect 198200 55214 198228 60030
rect 198464 57384 198516 57390
rect 198464 57326 198516 57332
rect 198200 55186 198320 55214
rect 197728 50380 197780 50386
rect 197728 50322 197780 50328
rect 197912 10600 197964 10606
rect 197912 10542 197964 10548
rect 197176 5432 197228 5438
rect 197176 5374 197228 5380
rect 196808 4956 196860 4962
rect 196808 4898 196860 4904
rect 195888 4684 195940 4690
rect 195888 4626 195940 4632
rect 196820 480 196848 4898
rect 197924 480 197952 10542
rect 198292 5370 198320 55186
rect 198476 10946 198504 57326
rect 198464 10940 198516 10946
rect 198464 10882 198516 10888
rect 198568 10878 198596 60030
rect 198660 56914 198688 60044
rect 198936 56914 198964 60044
rect 199212 57390 199240 60044
rect 199304 60030 199502 60058
rect 199870 60030 200068 60058
rect 199200 57384 199252 57390
rect 199200 57326 199252 57332
rect 198648 56908 198700 56914
rect 198648 56850 198700 56856
rect 198924 56908 198976 56914
rect 198924 56850 198976 56856
rect 199304 50658 199332 60030
rect 199844 57384 199896 57390
rect 199844 57326 199896 57332
rect 199292 50652 199344 50658
rect 199292 50594 199344 50600
rect 198556 10872 198608 10878
rect 198556 10814 198608 10820
rect 199856 10810 199884 57326
rect 199936 56908 199988 56914
rect 199936 56850 199988 56856
rect 199844 10804 199896 10810
rect 199844 10746 199896 10752
rect 199108 10532 199160 10538
rect 199108 10474 199160 10480
rect 198280 5364 198332 5370
rect 198280 5306 198332 5312
rect 199120 480 199148 10474
rect 199948 5302 199976 56850
rect 199936 5296 199988 5302
rect 199936 5238 199988 5244
rect 200040 5234 200068 60030
rect 200132 57390 200160 60044
rect 200120 57384 200172 57390
rect 200120 57326 200172 57332
rect 200408 51746 200436 60044
rect 200698 60030 200988 60058
rect 200960 55214 200988 60030
rect 201052 57526 201080 60044
rect 201144 60030 201342 60058
rect 201040 57520 201092 57526
rect 201040 57462 201092 57468
rect 200960 55186 201080 55214
rect 200396 51740 200448 51746
rect 200396 51682 200448 51688
rect 200028 5228 200080 5234
rect 200028 5170 200080 5176
rect 201052 4894 201080 55186
rect 201144 16250 201172 60030
rect 201316 57520 201368 57526
rect 201316 57462 201368 57468
rect 201224 57384 201276 57390
rect 201224 57326 201276 57332
rect 201132 16244 201184 16250
rect 201132 16186 201184 16192
rect 201236 10742 201264 57326
rect 201224 10736 201276 10742
rect 201224 10678 201276 10684
rect 201328 10674 201356 57462
rect 201604 57390 201632 60044
rect 201880 57866 201908 60044
rect 202262 60030 202460 60058
rect 202538 60030 202736 60058
rect 201868 57860 201920 57866
rect 201868 57802 201920 57808
rect 201592 57384 201644 57390
rect 201592 57326 201644 57332
rect 202432 16182 202460 60030
rect 202604 57860 202656 57866
rect 202604 57802 202656 57808
rect 202512 57520 202564 57526
rect 202512 57462 202564 57468
rect 202420 16176 202472 16182
rect 202420 16118 202472 16124
rect 201316 10668 201368 10674
rect 201316 10610 201368 10616
rect 202524 10606 202552 57462
rect 202616 10606 202644 57802
rect 202512 10600 202564 10606
rect 202512 10542 202564 10548
rect 202604 10600 202656 10606
rect 202604 10542 202656 10548
rect 202512 10464 202564 10470
rect 202512 10406 202564 10412
rect 201500 10396 201552 10402
rect 201500 10338 201552 10344
rect 201040 4888 201092 4894
rect 201040 4830 201092 4836
rect 200304 4752 200356 4758
rect 200304 4694 200356 4700
rect 200316 480 200344 4694
rect 201512 480 201540 10338
rect 202524 3482 202552 10406
rect 202708 6914 202736 60030
rect 202800 57526 202828 60044
rect 203076 57526 203104 60044
rect 202788 57520 202840 57526
rect 202788 57462 202840 57468
rect 203064 57520 203116 57526
rect 203064 57462 203116 57468
rect 203444 57390 203472 60044
rect 203720 57866 203748 60044
rect 203708 57860 203760 57866
rect 203708 57802 203760 57808
rect 203892 57520 203944 57526
rect 203892 57462 203944 57468
rect 202788 57384 202840 57390
rect 202788 57326 202840 57332
rect 203432 57384 203484 57390
rect 203432 57326 203484 57332
rect 202616 6886 202736 6914
rect 202616 5166 202644 6886
rect 202604 5160 202656 5166
rect 202604 5102 202656 5108
rect 202800 5098 202828 57326
rect 203904 16114 203932 57462
rect 203892 16108 203944 16114
rect 203892 16050 203944 16056
rect 203996 16046 204024 60044
rect 204076 57860 204128 57866
rect 204076 57802 204128 57808
rect 203984 16040 204036 16046
rect 203984 15982 204036 15988
rect 204088 10470 204116 57802
rect 204272 57390 204300 60044
rect 204548 57866 204576 60044
rect 204930 60030 205128 60058
rect 204536 57860 204588 57866
rect 204536 57802 204588 57808
rect 204168 57384 204220 57390
rect 204168 57326 204220 57332
rect 204260 57384 204312 57390
rect 204260 57326 204312 57332
rect 204076 10464 204128 10470
rect 204076 10406 204128 10412
rect 202788 5092 202840 5098
rect 202788 5034 202840 5040
rect 204180 4962 204208 57326
rect 205100 55214 205128 60030
rect 205192 57526 205220 60044
rect 205284 60030 205482 60058
rect 205180 57520 205232 57526
rect 205180 57462 205232 57468
rect 205100 55186 205220 55214
rect 205192 15978 205220 55186
rect 205180 15972 205232 15978
rect 205180 15914 205232 15920
rect 205284 10334 205312 60030
rect 205364 57860 205416 57866
rect 205364 57802 205416 57808
rect 205376 10402 205404 57802
rect 205744 57526 205772 60044
rect 206112 57866 206140 60044
rect 206100 57860 206152 57866
rect 206100 57802 206152 57808
rect 205456 57520 205508 57526
rect 205456 57462 205508 57468
rect 205732 57520 205784 57526
rect 205732 57462 205784 57468
rect 205364 10396 205416 10402
rect 205364 10338 205416 10344
rect 205088 10328 205140 10334
rect 205088 10270 205140 10276
rect 205272 10328 205324 10334
rect 205272 10270 205324 10276
rect 204168 4956 204220 4962
rect 204168 4898 204220 4904
rect 203892 4820 203944 4826
rect 203892 4762 203944 4768
rect 202524 3454 202736 3482
rect 202708 480 202736 3454
rect 203904 480 203932 4762
rect 205100 480 205128 10270
rect 205468 4826 205496 57462
rect 206388 57390 206416 60044
rect 206678 60030 206876 60058
rect 206744 57520 206796 57526
rect 206744 57462 206796 57468
rect 205548 57384 205600 57390
rect 205548 57326 205600 57332
rect 206376 57384 206428 57390
rect 206376 57326 206428 57332
rect 205560 4894 205588 57326
rect 206756 15910 206784 57462
rect 206192 15904 206244 15910
rect 206192 15846 206244 15852
rect 206744 15904 206796 15910
rect 206744 15846 206796 15852
rect 205548 4888 205600 4894
rect 205548 4830 205600 4836
rect 205456 4820 205508 4826
rect 205456 4762 205508 4768
rect 206204 480 206232 15846
rect 206848 3466 206876 60030
rect 206940 58018 206968 60044
rect 206940 57990 207060 58018
rect 206928 57860 206980 57866
rect 206928 57802 206980 57808
rect 206940 3534 206968 57802
rect 207032 56914 207060 57990
rect 207308 57361 207336 60044
rect 207294 57352 207350 57361
rect 207294 57287 207350 57296
rect 207020 56908 207072 56914
rect 207020 56850 207072 56856
rect 207584 56778 207612 60044
rect 207860 58818 207888 60044
rect 207848 58812 207900 58818
rect 207848 58754 207900 58760
rect 208136 58546 208164 60044
rect 208124 58540 208176 58546
rect 208124 58482 208176 58488
rect 208504 56953 208532 60044
rect 208780 57225 208808 60044
rect 209056 58614 209084 60044
rect 209044 58608 209096 58614
rect 209044 58550 209096 58556
rect 209332 57934 209360 60044
rect 209700 59838 209728 60044
rect 209688 59832 209740 59838
rect 209688 59774 209740 59780
rect 209320 57928 209372 57934
rect 209320 57870 209372 57876
rect 208766 57216 208822 57225
rect 208766 57151 208822 57160
rect 208490 56944 208546 56953
rect 208490 56879 208546 56888
rect 209136 56840 209188 56846
rect 209136 56782 209188 56788
rect 207572 56772 207624 56778
rect 207572 56714 207624 56720
rect 209044 56704 209096 56710
rect 209044 56646 209096 56652
rect 207020 55412 207072 55418
rect 207020 55354 207072 55360
rect 207032 16574 207060 55354
rect 209056 17270 209084 56646
rect 209148 19242 209176 56782
rect 209976 56710 210004 60044
rect 210252 59265 210280 60044
rect 210238 59256 210294 59265
rect 210238 59191 210294 59200
rect 210528 58478 210556 60044
rect 210516 58472 210568 58478
rect 210516 58414 210568 58420
rect 210424 56976 210476 56982
rect 210424 56918 210476 56924
rect 209964 56704 210016 56710
rect 209964 56646 210016 56652
rect 209780 55548 209832 55554
rect 209780 55490 209832 55496
rect 209136 19236 209188 19242
rect 209136 19178 209188 19184
rect 209044 17264 209096 17270
rect 209044 17206 209096 17212
rect 207032 16546 207428 16574
rect 206928 3528 206980 3534
rect 206928 3470 206980 3476
rect 206836 3460 206888 3466
rect 206836 3402 206888 3408
rect 207400 480 207428 16546
rect 208584 9784 208636 9790
rect 208584 9726 208636 9732
rect 208596 480 208624 9726
rect 209792 4078 209820 55490
rect 210436 47666 210464 56918
rect 210896 56846 210924 60044
rect 211172 57497 211200 60044
rect 211448 58682 211476 60044
rect 211724 58886 211752 60044
rect 212000 59362 212028 60044
rect 212368 59401 212396 60044
rect 212644 59770 212672 60044
rect 212632 59764 212684 59770
rect 212632 59706 212684 59712
rect 212354 59392 212410 59401
rect 211988 59356 212040 59362
rect 212354 59327 212410 59336
rect 211988 59298 212040 59304
rect 211712 58880 211764 58886
rect 211712 58822 211764 58828
rect 211436 58676 211488 58682
rect 211436 58618 211488 58624
rect 211158 57488 211214 57497
rect 211158 57423 211214 57432
rect 210884 56840 210936 56846
rect 210884 56782 210936 56788
rect 212920 56642 212948 60044
rect 213196 59226 213224 60044
rect 213184 59220 213236 59226
rect 213184 59162 213236 59168
rect 213564 58342 213592 60044
rect 213552 58336 213604 58342
rect 213552 58278 213604 58284
rect 213184 57724 213236 57730
rect 213184 57666 213236 57672
rect 212908 56636 212960 56642
rect 212908 56578 212960 56584
rect 210424 47660 210476 47666
rect 210424 47602 210476 47608
rect 213196 19990 213224 57666
rect 213276 57656 213328 57662
rect 213276 57598 213328 57604
rect 213288 20194 213316 57598
rect 213840 57089 213868 60044
rect 214116 58954 214144 60044
rect 214104 58948 214156 58954
rect 214104 58890 214156 58896
rect 214392 58274 214420 60044
rect 214380 58268 214432 58274
rect 214380 58210 214432 58216
rect 214760 57905 214788 60044
rect 214746 57896 214802 57905
rect 214746 57831 214802 57840
rect 214564 57792 214616 57798
rect 214564 57734 214616 57740
rect 213826 57080 213882 57089
rect 213826 57015 213882 57024
rect 213920 55344 213972 55350
rect 213920 55286 213972 55292
rect 213276 20188 213328 20194
rect 213276 20130 213328 20136
rect 213184 19984 213236 19990
rect 213184 19926 213236 19932
rect 213932 16574 213960 55286
rect 214576 21418 214604 57734
rect 215036 56982 215064 60044
rect 215312 57662 215340 60044
rect 215588 58206 215616 60044
rect 215956 59362 215984 60044
rect 215944 59356 215996 59362
rect 215944 59298 215996 59304
rect 215576 58200 215628 58206
rect 215576 58142 215628 58148
rect 216232 58070 216260 60044
rect 216220 58064 216272 58070
rect 216220 58006 216272 58012
rect 216508 57769 216536 60044
rect 216784 58138 216812 60044
rect 217152 59294 217180 60044
rect 217140 59288 217192 59294
rect 217140 59230 217192 59236
rect 216772 58132 216824 58138
rect 216772 58074 216824 58080
rect 216494 57760 216550 57769
rect 217428 57730 217456 60044
rect 217704 58750 217732 60044
rect 217692 58744 217744 58750
rect 217692 58686 217744 58692
rect 216494 57695 216550 57704
rect 217416 57724 217468 57730
rect 217416 57666 217468 57672
rect 215300 57656 215352 57662
rect 215300 57598 215352 57604
rect 217980 57526 218008 60044
rect 218256 57905 218284 60044
rect 218624 59158 218652 60044
rect 218612 59152 218664 59158
rect 218612 59094 218664 59100
rect 218242 57896 218298 57905
rect 218242 57831 218298 57840
rect 218900 57594 218928 60044
rect 219176 59702 219204 60044
rect 219466 60030 219756 60058
rect 219164 59696 219216 59702
rect 219164 59638 219216 59644
rect 219728 57905 219756 60030
rect 219820 59022 219848 60044
rect 219808 59016 219860 59022
rect 219808 58958 219860 58964
rect 220096 57934 220124 60044
rect 220084 57928 220136 57934
rect 219530 57896 219586 57905
rect 219530 57831 219586 57840
rect 219714 57896 219770 57905
rect 220084 57870 220136 57876
rect 220372 57866 220400 60044
rect 219714 57831 219770 57840
rect 220360 57860 220412 57866
rect 219544 57633 219572 57831
rect 220360 57802 220412 57808
rect 220648 57798 220676 60044
rect 221016 59634 221044 60044
rect 221004 59628 221056 59634
rect 221004 59570 221056 59576
rect 221292 59226 221320 60044
rect 221844 59498 221872 60044
rect 221832 59492 221884 59498
rect 221832 59434 221884 59440
rect 221280 59220 221332 59226
rect 221280 59162 221332 59168
rect 222212 59090 222240 60044
rect 222488 59566 222516 60044
rect 222778 60030 222934 60058
rect 223054 60030 223344 60058
rect 222934 60007 222990 60016
rect 223316 59945 223344 60030
rect 223302 59936 223358 59945
rect 223302 59871 223358 59880
rect 222476 59560 222528 59566
rect 222476 59502 222528 59508
rect 222200 59084 222252 59090
rect 222200 59026 222252 59032
rect 220636 57792 220688 57798
rect 220636 57734 220688 57740
rect 219530 57624 219586 57633
rect 218888 57588 218940 57594
rect 219530 57559 219586 57568
rect 218888 57530 218940 57536
rect 215944 57520 215996 57526
rect 215944 57462 215996 57468
rect 217968 57520 218020 57526
rect 217968 57462 218020 57468
rect 215024 56976 215076 56982
rect 215024 56918 215076 56924
rect 214564 21412 214616 21418
rect 214564 21354 214616 21360
rect 213932 16546 214512 16574
rect 213368 15428 213420 15434
rect 213368 15370 213420 15376
rect 209872 15360 209924 15366
rect 209872 15302 209924 15308
rect 209780 4072 209832 4078
rect 209780 4014 209832 4020
rect 209884 3482 209912 15302
rect 212172 9852 212224 9858
rect 212172 9794 212224 9800
rect 210976 4072 211028 4078
rect 210976 4014 211028 4020
rect 209792 3454 209912 3482
rect 209792 480 209820 3454
rect 210988 480 211016 4014
rect 212184 480 212212 9794
rect 213380 480 213408 15370
rect 214484 480 214512 16546
rect 215956 10130 215984 57462
rect 220084 57452 220136 57458
rect 220084 57394 220136 57400
rect 216036 57180 216088 57186
rect 216036 57122 216088 57128
rect 216048 24206 216076 57122
rect 217324 57112 217376 57118
rect 217324 57054 217376 57060
rect 216036 24200 216088 24206
rect 216036 24142 216088 24148
rect 217336 22778 217364 57054
rect 218060 55616 218112 55622
rect 218060 55558 218112 55564
rect 217324 22772 217376 22778
rect 217324 22714 217376 22720
rect 216864 15496 216916 15502
rect 216864 15438 216916 15444
rect 215668 10124 215720 10130
rect 215668 10066 215720 10072
rect 215944 10124 215996 10130
rect 215944 10066 215996 10072
rect 215680 480 215708 10066
rect 216876 480 216904 15438
rect 218072 480 218100 55558
rect 220096 20058 220124 57394
rect 223408 57186 223436 60044
rect 223684 59906 223712 60044
rect 223672 59900 223724 59906
rect 223672 59842 223724 59848
rect 223960 59430 223988 60044
rect 224236 59906 224264 60044
rect 224224 59900 224276 59906
rect 224224 59842 224276 59848
rect 223948 59424 224000 59430
rect 223948 59366 224000 59372
rect 224512 58070 224540 398754
rect 225420 397860 225472 397866
rect 225420 397802 225472 397808
rect 224960 397452 225012 397458
rect 224960 397394 225012 397400
rect 224776 396908 224828 396914
rect 224776 396850 224828 396856
rect 224590 232928 224646 232937
rect 224590 232863 224646 232872
rect 224604 60217 224632 232863
rect 224682 230072 224738 230081
rect 224682 230007 224738 230016
rect 224590 60208 224646 60217
rect 224590 60143 224646 60152
rect 224500 58064 224552 58070
rect 224500 58006 224552 58012
rect 224696 57934 224724 230007
rect 224788 225049 224816 396850
rect 224868 396364 224920 396370
rect 224868 396306 224920 396312
rect 224880 226681 224908 396306
rect 224866 226672 224922 226681
rect 224866 226607 224922 226616
rect 224774 225040 224830 225049
rect 224774 224975 224830 224984
rect 224972 59401 225000 397394
rect 225052 249280 225104 249286
rect 225052 249222 225104 249228
rect 224958 59392 225014 59401
rect 224958 59327 225014 59336
rect 224684 57928 224736 57934
rect 224684 57870 224736 57876
rect 223396 57180 223448 57186
rect 223396 57122 223448 57128
rect 220176 57044 220228 57050
rect 220176 56986 220228 56992
rect 220188 24138 220216 56986
rect 225064 56642 225092 249222
rect 225236 242140 225288 242146
rect 225236 242082 225288 242088
rect 225144 241936 225196 241942
rect 225144 241878 225196 241884
rect 225156 57866 225184 241878
rect 225144 57860 225196 57866
rect 225144 57802 225196 57808
rect 225248 57730 225276 242082
rect 225326 232792 225382 232801
rect 225326 232727 225382 232736
rect 225236 57724 225288 57730
rect 225236 57666 225288 57672
rect 225340 57089 225368 232727
rect 225432 222601 225460 397802
rect 226064 242888 226116 242894
rect 226064 242830 226116 242836
rect 225972 241256 226024 241262
rect 225972 241198 226024 241204
rect 225510 230480 225566 230489
rect 225510 230415 225566 230424
rect 225418 222592 225474 222601
rect 225418 222527 225474 222536
rect 225524 60081 225552 230415
rect 225602 229936 225658 229945
rect 225602 229871 225658 229880
rect 225510 60072 225566 60081
rect 225510 60007 225566 60016
rect 225616 57905 225644 229871
rect 225694 229800 225750 229809
rect 225694 229735 225750 229744
rect 225602 57896 225658 57905
rect 225602 57831 225658 57840
rect 225708 57798 225736 229735
rect 225878 227352 225934 227361
rect 225878 227287 225934 227296
rect 225786 226808 225842 226817
rect 225786 226743 225842 226752
rect 225800 59945 225828 226743
rect 225786 59936 225842 59945
rect 225786 59871 225842 59880
rect 225696 57792 225748 57798
rect 225892 57769 225920 227287
rect 225984 131209 226012 241198
rect 226076 141953 226104 242830
rect 226156 240712 226208 240718
rect 226156 240654 226208 240660
rect 226168 195673 226196 240654
rect 226246 230208 226302 230217
rect 226246 230143 226302 230152
rect 226154 195664 226210 195673
rect 226154 195599 226210 195608
rect 226062 141944 226118 141953
rect 226062 141879 226118 141888
rect 225970 131200 226026 131209
rect 225970 131135 226026 131144
rect 225696 57734 225748 57740
rect 225878 57760 225934 57769
rect 225878 57695 225934 57704
rect 226260 57633 226288 230143
rect 226352 109585 226380 399842
rect 230480 399832 230532 399838
rect 230480 399774 230532 399780
rect 227720 398744 227772 398750
rect 227720 398686 227772 398692
rect 226616 398608 226668 398614
rect 226616 398550 226668 398556
rect 226432 398064 226484 398070
rect 226432 398006 226484 398012
rect 226444 139233 226472 398006
rect 226524 397996 226576 398002
rect 226524 397938 226576 397944
rect 226536 149977 226564 397938
rect 226628 158001 226656 398550
rect 226708 398540 226760 398546
rect 226708 398482 226760 398488
rect 226720 182209 226748 398482
rect 226892 249620 226944 249626
rect 226892 249562 226944 249568
rect 226800 240168 226852 240174
rect 226800 240110 226852 240116
rect 226706 182200 226762 182209
rect 226706 182135 226762 182144
rect 226706 175264 226762 175273
rect 226706 175199 226762 175208
rect 226720 174185 226748 175199
rect 226706 174176 226762 174185
rect 226706 174111 226762 174120
rect 226706 169688 226762 169697
rect 226706 169623 226762 169632
rect 226720 168745 226748 169623
rect 226706 168736 226762 168745
rect 226706 168671 226762 168680
rect 226614 157992 226670 158001
rect 226614 157927 226670 157936
rect 226522 149968 226578 149977
rect 226522 149903 226578 149912
rect 226430 139224 226486 139233
rect 226430 139159 226486 139168
rect 226430 126984 226486 126993
rect 226430 126919 226486 126928
rect 226444 125769 226472 126919
rect 226430 125760 226486 125769
rect 226430 125695 226486 125704
rect 226338 109576 226394 109585
rect 226338 109511 226394 109520
rect 226430 73128 226486 73137
rect 226430 73063 226486 73072
rect 226444 72049 226472 73063
rect 226430 72040 226486 72049
rect 226430 71975 226486 71984
rect 226812 63889 226840 240110
rect 226904 88097 226932 249562
rect 226984 241052 227036 241058
rect 226984 240994 227036 241000
rect 226890 88088 226946 88097
rect 226890 88023 226946 88032
rect 226996 80073 227024 240994
rect 227074 235240 227130 235249
rect 227074 235175 227130 235184
rect 227088 128489 227116 235175
rect 227534 233200 227590 233209
rect 227534 233135 227590 233144
rect 227442 232656 227498 232665
rect 227442 232591 227498 232600
rect 227350 227216 227406 227225
rect 227350 227151 227406 227160
rect 227258 227080 227314 227089
rect 227258 227015 227314 227024
rect 227166 225040 227222 225049
rect 227166 224975 227222 224984
rect 227180 220969 227208 224975
rect 227166 220960 227222 220969
rect 227166 220895 227222 220904
rect 227166 220824 227222 220833
rect 227166 220759 227222 220768
rect 227180 219881 227208 220759
rect 227166 219872 227222 219881
rect 227166 219807 227222 219816
rect 227166 219736 227222 219745
rect 227166 219671 227222 219680
rect 227074 128480 227130 128489
rect 227074 128415 227130 128424
rect 227180 123049 227208 219671
rect 227272 144673 227300 227015
rect 227364 166161 227392 227151
rect 227456 198393 227484 232591
rect 227548 217161 227576 233135
rect 227626 228304 227682 228313
rect 227626 228239 227682 228248
rect 227640 219745 227668 228239
rect 227626 219736 227682 219745
rect 227626 219671 227682 219680
rect 227626 219600 227682 219609
rect 227626 219535 227682 219544
rect 227534 217152 227590 217161
rect 227534 217087 227590 217096
rect 227640 214577 227668 219535
rect 227626 214568 227682 214577
rect 227626 214503 227682 214512
rect 227534 212528 227590 212537
rect 227534 212463 227590 212472
rect 227548 211857 227576 212463
rect 227534 211848 227590 211857
rect 227534 211783 227590 211792
rect 227442 198384 227498 198393
rect 227442 198319 227498 198328
rect 227350 166152 227406 166161
rect 227350 166087 227406 166096
rect 227258 144664 227314 144673
rect 227258 144599 227314 144608
rect 227166 123040 227222 123049
rect 227166 122975 227222 122984
rect 226982 80064 227038 80073
rect 226982 79999 227038 80008
rect 226798 63880 226854 63889
rect 226798 63815 226854 63824
rect 227732 58138 227760 398686
rect 229284 398676 229336 398682
rect 229284 398618 229336 398624
rect 229192 398472 229244 398478
rect 229192 398414 229244 398420
rect 229100 398404 229152 398410
rect 229100 398346 229152 398352
rect 227812 398336 227864 398342
rect 227812 398278 227864 398284
rect 227824 59294 227852 398278
rect 228364 398268 228416 398274
rect 228364 398210 228416 398216
rect 228272 398200 228324 398206
rect 228272 398142 228324 398148
rect 228088 397928 228140 397934
rect 228088 397870 228140 397876
rect 227904 396568 227956 396574
rect 227904 396510 227956 396516
rect 227916 59362 227944 396510
rect 227996 395480 228048 395486
rect 227996 395422 228048 395428
rect 227904 59356 227956 59362
rect 227904 59298 227956 59304
rect 227812 59288 227864 59294
rect 227812 59230 227864 59236
rect 227720 58132 227772 58138
rect 227720 58074 227772 58080
rect 226246 57624 226302 57633
rect 228008 57594 228036 395422
rect 228100 163441 228128 397870
rect 228180 395412 228232 395418
rect 228180 395354 228232 395360
rect 228086 163432 228142 163441
rect 228086 163367 228142 163376
rect 228192 160721 228220 395354
rect 228284 171465 228312 398142
rect 228376 179625 228404 398210
rect 228640 398132 228692 398138
rect 228640 398074 228692 398080
rect 228456 397792 228508 397798
rect 228456 397734 228508 397740
rect 228468 184929 228496 397734
rect 228548 246288 228600 246294
rect 228548 246230 228600 246236
rect 228454 184920 228510 184929
rect 228454 184855 228510 184864
rect 228362 179616 228418 179625
rect 228362 179551 228418 179560
rect 228270 171456 228326 171465
rect 228270 171391 228326 171400
rect 228178 160712 228234 160721
rect 228178 160647 228234 160656
rect 228086 91760 228142 91769
rect 228086 91695 228142 91704
rect 228100 90817 228128 91695
rect 228086 90808 228142 90817
rect 228086 90743 228142 90752
rect 226246 57559 226302 57568
rect 227996 57588 228048 57594
rect 227996 57530 228048 57536
rect 228560 57526 228588 246230
rect 228652 209137 228680 398074
rect 228916 367804 228968 367810
rect 228916 367746 228968 367752
rect 228824 246900 228876 246906
rect 228824 246842 228876 246848
rect 228732 245472 228784 245478
rect 228732 245414 228784 245420
rect 228638 209128 228694 209137
rect 228638 209063 228694 209072
rect 228548 57520 228600 57526
rect 228548 57462 228600 57468
rect 225326 57080 225382 57089
rect 225326 57015 225382 57024
rect 228744 56982 228772 245414
rect 228836 74633 228864 246842
rect 228928 206417 228956 367746
rect 229008 241324 229060 241330
rect 229008 241266 229060 241272
rect 228914 206408 228970 206417
rect 228914 206343 228970 206352
rect 229020 176905 229048 241266
rect 229006 176896 229062 176905
rect 229006 176831 229062 176840
rect 228822 74624 228878 74633
rect 228822 74559 228878 74568
rect 229112 59022 229140 398346
rect 229100 59016 229152 59022
rect 229100 58958 229152 58964
rect 229204 58342 229232 398414
rect 229296 58546 229324 398618
rect 229376 397384 229428 397390
rect 229376 397326 229428 397332
rect 229284 58540 229336 58546
rect 229284 58482 229336 58488
rect 229388 58478 229416 397326
rect 229468 396636 229520 396642
rect 229468 396578 229520 396584
rect 229480 58750 229508 396578
rect 229652 261520 229704 261526
rect 229652 261462 229704 261468
rect 229558 226944 229614 226953
rect 229558 226879 229614 226888
rect 229468 58744 229520 58750
rect 229468 58686 229520 58692
rect 229376 58472 229428 58478
rect 229376 58414 229428 58420
rect 229192 58336 229244 58342
rect 229192 58278 229244 58284
rect 228732 56976 228784 56982
rect 228732 56918 228784 56924
rect 229572 56778 229600 226879
rect 229664 104281 229692 261462
rect 229744 248056 229796 248062
rect 229744 247998 229796 248004
rect 229650 104272 229706 104281
rect 229650 104207 229706 104216
rect 229756 98841 229784 247998
rect 229836 246968 229888 246974
rect 229836 246910 229888 246916
rect 229848 117745 229876 246910
rect 229926 233472 229982 233481
rect 229926 233407 229982 233416
rect 229940 151881 229968 233407
rect 229926 151872 229982 151881
rect 229926 151807 229982 151816
rect 229834 117736 229890 117745
rect 229834 117671 229890 117680
rect 229742 98832 229798 98841
rect 229742 98767 229798 98776
rect 230492 57118 230520 399774
rect 233240 399764 233292 399770
rect 233240 399706 233292 399712
rect 232044 399696 232096 399702
rect 232044 399638 232096 399644
rect 231952 399628 232004 399634
rect 231952 399570 232004 399576
rect 231860 396704 231912 396710
rect 231860 396646 231912 396652
rect 231124 395616 231176 395622
rect 231124 395558 231176 395564
rect 230664 249212 230716 249218
rect 230664 249154 230716 249160
rect 230572 242412 230624 242418
rect 230572 242354 230624 242360
rect 230480 57112 230532 57118
rect 230480 57054 230532 57060
rect 229560 56772 229612 56778
rect 229560 56714 229612 56720
rect 230584 56710 230612 242354
rect 230676 152697 230704 249154
rect 230756 241460 230808 241466
rect 230756 241402 230808 241408
rect 230768 190369 230796 241402
rect 230754 190360 230810 190369
rect 230754 190295 230810 190304
rect 230662 152688 230718 152697
rect 230662 152623 230718 152632
rect 231136 112305 231164 395558
rect 231214 234696 231270 234705
rect 231214 234631 231270 234640
rect 231228 178129 231256 234631
rect 231214 178120 231270 178129
rect 231214 178055 231270 178064
rect 231122 112296 231178 112305
rect 231122 112231 231178 112240
rect 231872 59158 231900 396646
rect 231964 61305 231992 399570
rect 232056 96257 232084 399638
rect 232504 395412 232556 395418
rect 232504 395354 232556 395360
rect 232320 245608 232372 245614
rect 232320 245550 232372 245556
rect 232228 244860 232280 244866
rect 232228 244802 232280 244808
rect 232136 241120 232188 241126
rect 232136 241062 232188 241068
rect 232042 96248 232098 96257
rect 232042 96183 232098 96192
rect 232148 93537 232176 241062
rect 232240 101561 232268 244802
rect 232332 120465 232360 245550
rect 232516 126993 232544 395354
rect 232688 250504 232740 250510
rect 232688 250446 232740 250452
rect 232594 232112 232650 232121
rect 232594 232047 232650 232056
rect 232502 126984 232558 126993
rect 232502 126919 232558 126928
rect 232318 120456 232374 120465
rect 232318 120391 232374 120400
rect 232226 101552 232282 101561
rect 232226 101487 232282 101496
rect 232134 93528 232190 93537
rect 232134 93463 232190 93472
rect 232608 71913 232636 232047
rect 232700 212537 232728 250446
rect 232686 212528 232742 212537
rect 232686 212463 232742 212472
rect 232594 71904 232650 71913
rect 232594 71839 232650 71848
rect 231950 61296 232006 61305
rect 231950 61231 232006 61240
rect 233252 60058 233280 399706
rect 235998 398168 236054 398177
rect 235998 398103 236054 398112
rect 265070 398168 265126 398177
rect 265070 398103 265126 398112
rect 300122 398168 300178 398177
rect 300122 398103 300178 398112
rect 315762 398168 315818 398177
rect 315762 398103 315818 398112
rect 325882 398168 325938 398177
rect 325882 398103 325938 398112
rect 233424 396840 233476 396846
rect 233424 396782 233476 396788
rect 233332 396772 233384 396778
rect 233332 396714 233384 396720
rect 233160 60030 233280 60058
rect 233160 59650 233188 60030
rect 233344 59906 233372 396714
rect 233240 59900 233292 59906
rect 233240 59842 233292 59848
rect 233332 59900 233384 59906
rect 233332 59842 233384 59848
rect 233252 59786 233280 59842
rect 233436 59786 233464 396782
rect 236012 396302 236040 398103
rect 237010 397352 237066 397361
rect 237010 397287 237066 397296
rect 238114 397352 238170 397361
rect 238114 397287 238170 397296
rect 239218 397352 239274 397361
rect 239218 397287 239274 397296
rect 240506 397352 240562 397361
rect 240506 397287 240562 397296
rect 241610 397352 241666 397361
rect 241610 397287 241666 397296
rect 247682 397352 247738 397361
rect 247682 397287 247738 397296
rect 249982 397352 250038 397361
rect 249982 397287 250038 397296
rect 251178 397352 251234 397361
rect 251178 397287 251234 397296
rect 252742 397352 252798 397361
rect 252742 397287 252798 397296
rect 259826 397352 259882 397361
rect 259826 397287 259882 397296
rect 262034 397352 262090 397361
rect 262034 397287 262090 397296
rect 237024 397186 237052 397287
rect 238024 397248 238076 397254
rect 238024 397190 238076 397196
rect 237012 397180 237064 397186
rect 237012 397122 237064 397128
rect 236000 396296 236052 396302
rect 236000 396238 236052 396244
rect 235264 395752 235316 395758
rect 235264 395694 235316 395700
rect 233516 395344 233568 395350
rect 233516 395286 233568 395292
rect 233528 77353 233556 395286
rect 233700 249144 233752 249150
rect 233700 249086 233752 249092
rect 233608 247036 233660 247042
rect 233608 246978 233660 246984
rect 233514 77344 233570 77353
rect 233514 77279 233570 77288
rect 233252 59758 233464 59786
rect 233160 59622 233280 59650
rect 231860 59152 231912 59158
rect 231860 59094 231912 59100
rect 233252 56846 233280 59622
rect 233620 57186 233648 246978
rect 233712 66609 233740 249086
rect 233882 193896 233938 193905
rect 233882 193831 233938 193840
rect 233896 192953 233924 193831
rect 233882 192944 233938 192953
rect 233882 192879 233938 192888
rect 235276 73137 235304 395694
rect 235356 240984 235408 240990
rect 235356 240926 235408 240932
rect 235368 203833 235396 240926
rect 235354 203824 235410 203833
rect 235354 203759 235410 203768
rect 235262 73128 235318 73137
rect 235262 73063 235318 73072
rect 233698 66600 233754 66609
rect 233698 66535 233754 66544
rect 238036 58614 238064 397190
rect 238128 397050 238156 397287
rect 239232 397254 239260 397287
rect 239220 397248 239272 397254
rect 239220 397190 239272 397196
rect 238116 397044 238168 397050
rect 238116 396986 238168 396992
rect 238208 396296 238260 396302
rect 238208 396238 238260 396244
rect 238116 395480 238168 395486
rect 238116 395422 238168 395428
rect 238128 133793 238156 395422
rect 238220 240650 238248 396238
rect 240520 396234 240548 397287
rect 240784 396772 240836 396778
rect 240784 396714 240836 396720
rect 240508 396228 240560 396234
rect 240508 396170 240560 396176
rect 238208 240644 238260 240650
rect 238208 240586 238260 240592
rect 238114 133784 238170 133793
rect 238114 133719 238170 133728
rect 240796 58818 240824 396714
rect 241624 395826 241652 397287
rect 247696 397118 247724 397287
rect 247684 397112 247736 397118
rect 247684 397054 247736 397060
rect 242898 396808 242954 396817
rect 242898 396743 242900 396752
rect 242952 396743 242954 396752
rect 244370 396808 244426 396817
rect 244370 396743 244426 396752
rect 245658 396808 245714 396817
rect 245658 396743 245714 396752
rect 247590 396808 247646 396817
rect 247590 396743 247646 396752
rect 248418 396808 248474 396817
rect 249798 396808 249854 396817
rect 248418 396743 248474 396752
rect 249064 396772 249116 396778
rect 242900 396714 242952 396720
rect 244278 396672 244334 396681
rect 244278 396607 244334 396616
rect 242256 396228 242308 396234
rect 242256 396170 242308 396176
rect 242164 396024 242216 396030
rect 242164 395966 242216 395972
rect 241612 395820 241664 395826
rect 241612 395762 241664 395768
rect 240876 395344 240928 395350
rect 240876 395286 240928 395292
rect 240888 155961 240916 395286
rect 240968 241528 241020 241534
rect 240968 241470 241020 241476
rect 240980 167006 241008 241470
rect 240968 167000 241020 167006
rect 240968 166942 241020 166948
rect 240874 155952 240930 155961
rect 240874 155887 240930 155896
rect 240784 58812 240836 58818
rect 240784 58754 240836 58760
rect 238024 58608 238076 58614
rect 238024 58550 238076 58556
rect 233608 57180 233660 57186
rect 233608 57122 233660 57128
rect 242176 56914 242204 395966
rect 242268 243506 242296 396170
rect 242256 243500 242308 243506
rect 242256 243442 242308 243448
rect 242256 241596 242308 241602
rect 242256 241538 242308 241544
rect 242268 206990 242296 241538
rect 242256 206984 242308 206990
rect 242256 206926 242308 206932
rect 244292 82793 244320 396607
rect 244384 240922 244412 396743
rect 244372 240916 244424 240922
rect 244372 240858 244424 240864
rect 244924 225616 244976 225622
rect 244924 225558 244976 225564
rect 244936 147665 244964 225558
rect 244922 147656 244978 147665
rect 244922 147591 244978 147600
rect 244278 82784 244334 82793
rect 244278 82719 244334 82728
rect 245672 58886 245700 396743
rect 246304 396568 246356 396574
rect 246304 396510 246356 396516
rect 246316 169697 246344 396510
rect 247604 396030 247632 396743
rect 247592 396024 247644 396030
rect 247592 395966 247644 395972
rect 246302 169688 246358 169697
rect 246302 169623 246358 169632
rect 248432 58954 248460 396743
rect 249798 396743 249854 396752
rect 249064 396714 249116 396720
rect 249076 241398 249104 396714
rect 249064 241392 249116 241398
rect 249064 241334 249116 241340
rect 249812 240854 249840 396743
rect 249996 395758 250024 397287
rect 249984 395752 250036 395758
rect 249984 395694 250036 395700
rect 249800 240848 249852 240854
rect 249800 240790 249852 240796
rect 248420 58948 248472 58954
rect 248420 58890 248472 58896
rect 245660 58880 245712 58886
rect 245660 58822 245712 58828
rect 251192 58206 251220 397287
rect 251270 397216 251326 397225
rect 251270 397151 251326 397160
rect 251284 396982 251312 397151
rect 251272 396976 251324 396982
rect 251272 396918 251324 396924
rect 252650 396808 252706 396817
rect 252650 396743 252706 396752
rect 252664 59838 252692 396743
rect 252756 396166 252784 397287
rect 258078 396944 258134 396953
rect 258078 396879 258134 396888
rect 254490 396808 254546 396817
rect 254490 396743 254546 396752
rect 255410 396808 255466 396817
rect 255410 396743 255466 396752
rect 256882 396808 256938 396817
rect 256882 396743 256884 396752
rect 254504 396710 254532 396743
rect 253204 396704 253256 396710
rect 253204 396646 253256 396652
rect 254492 396704 254544 396710
rect 254492 396646 254544 396652
rect 255318 396672 255374 396681
rect 252744 396160 252796 396166
rect 252744 396102 252796 396108
rect 253216 136649 253244 396646
rect 255318 396607 255374 396616
rect 253202 136640 253258 136649
rect 253202 136575 253258 136584
rect 255332 91769 255360 396607
rect 255424 225622 255452 396743
rect 256936 396743 256938 396752
rect 256884 396714 256936 396720
rect 255412 225616 255464 225622
rect 255412 225558 255464 225564
rect 255318 91760 255374 91769
rect 255318 91695 255374 91704
rect 252652 59832 252704 59838
rect 252652 59774 252704 59780
rect 258092 59770 258120 396879
rect 258170 396808 258226 396817
rect 258170 396743 258226 396752
rect 259550 396808 259606 396817
rect 259550 396743 259606 396752
rect 258184 241194 258212 396743
rect 259564 249082 259592 396743
rect 259840 396234 259868 397287
rect 260930 396808 260986 396817
rect 260930 396743 260986 396752
rect 260944 396710 260972 396743
rect 260104 396704 260156 396710
rect 260104 396646 260156 396652
rect 260932 396704 260984 396710
rect 260932 396646 260984 396652
rect 259828 396228 259880 396234
rect 259828 396170 259880 396176
rect 259552 249076 259604 249082
rect 259552 249018 259604 249024
rect 258172 241188 258224 241194
rect 258172 241130 258224 241136
rect 258080 59764 258132 59770
rect 258080 59706 258132 59712
rect 260116 58410 260144 396646
rect 262048 396574 262076 397287
rect 262218 396808 262274 396817
rect 262218 396743 262274 396752
rect 263598 396808 263654 396817
rect 263598 396743 263654 396752
rect 262036 396568 262088 396574
rect 262036 396510 262088 396516
rect 262232 175273 262260 396743
rect 262218 175264 262274 175273
rect 262218 175199 262274 175208
rect 260104 58404 260156 58410
rect 260104 58346 260156 58352
rect 263612 58274 263640 396743
rect 263690 396672 263746 396681
rect 263690 396607 263746 396616
rect 263704 242690 263732 396607
rect 265084 247926 265112 398103
rect 265898 397352 265954 397361
rect 265898 397287 265954 397296
rect 268290 397352 268346 397361
rect 268290 397287 268346 397296
rect 270866 397352 270922 397361
rect 270866 397287 270922 397296
rect 272246 397352 272302 397361
rect 272246 397287 272302 397296
rect 273442 397352 273498 397361
rect 273442 397287 273498 397296
rect 276202 397352 276258 397361
rect 276202 397287 276258 397296
rect 276386 397352 276442 397361
rect 276386 397287 276442 397296
rect 278042 397352 278098 397361
rect 278042 397287 278044 397296
rect 265912 395622 265940 397287
rect 266358 396808 266414 396817
rect 266358 396743 266414 396752
rect 267830 396808 267886 396817
rect 267830 396743 267886 396752
rect 265900 395616 265952 395622
rect 265900 395558 265952 395564
rect 265072 247920 265124 247926
rect 265072 247862 265124 247868
rect 263692 242684 263744 242690
rect 263692 242626 263744 242632
rect 266372 242350 266400 396743
rect 266450 396672 266506 396681
rect 266450 396607 266506 396616
rect 266464 245274 266492 396607
rect 266452 245268 266504 245274
rect 266452 245210 266504 245216
rect 266360 242344 266412 242350
rect 266360 242286 266412 242292
rect 267844 193905 267872 396743
rect 268304 395690 268332 397287
rect 269118 396808 269174 396817
rect 268384 396772 268436 396778
rect 269118 396743 269174 396752
rect 270590 396808 270646 396817
rect 270590 396743 270646 396752
rect 268384 396714 268436 396720
rect 268292 395684 268344 395690
rect 268292 395626 268344 395632
rect 267830 193896 267886 193905
rect 267830 193831 267886 193840
rect 268396 59090 268424 396714
rect 269132 59226 269160 396743
rect 270604 240990 270632 396743
rect 270880 395418 270908 397287
rect 272260 396302 272288 397287
rect 273350 397216 273406 397225
rect 273350 397151 273406 397160
rect 273258 396808 273314 396817
rect 273258 396743 273260 396752
rect 273312 396743 273314 396752
rect 273260 396714 273312 396720
rect 272248 396296 272300 396302
rect 272248 396238 272300 396244
rect 273364 395486 273392 397151
rect 273456 396438 273484 397287
rect 274638 396808 274694 396817
rect 274638 396743 274694 396752
rect 273444 396432 273496 396438
rect 273444 396374 273496 396380
rect 273352 395480 273404 395486
rect 273352 395422 273404 395428
rect 270868 395412 270920 395418
rect 270868 395354 270920 395360
rect 270592 240984 270644 240990
rect 270592 240926 270644 240932
rect 274652 240786 274680 396743
rect 276216 395554 276244 397287
rect 276400 396506 276428 397287
rect 278096 397287 278098 397296
rect 278962 397352 279018 397361
rect 278962 397287 279018 397296
rect 283194 397352 283250 397361
rect 283194 397287 283250 397296
rect 289818 397352 289874 397361
rect 289818 397287 289874 397296
rect 298466 397352 298522 397361
rect 298466 397287 298522 397296
rect 278044 397258 278096 397264
rect 277490 396808 277546 396817
rect 277490 396743 277546 396752
rect 276388 396500 276440 396506
rect 276388 396442 276440 396448
rect 276204 395548 276256 395554
rect 276204 395490 276256 395496
rect 277504 247858 277532 396743
rect 278976 396370 279004 397287
rect 280158 396808 280214 396817
rect 280158 396743 280214 396752
rect 278964 396364 279016 396370
rect 278964 396306 279016 396312
rect 277492 247852 277544 247858
rect 277492 247794 277544 247800
rect 280172 246838 280200 396743
rect 282184 396296 282236 396302
rect 282184 396238 282236 396244
rect 280160 246832 280212 246838
rect 280160 246774 280212 246780
rect 274640 240780 274692 240786
rect 274640 240722 274692 240728
rect 278042 230752 278098 230761
rect 278042 230687 278098 230696
rect 271142 229256 271198 229265
rect 271142 229191 271198 229200
rect 271156 126954 271184 229191
rect 278056 193186 278084 230687
rect 282196 220833 282224 396238
rect 283208 395350 283236 397287
rect 285678 396808 285734 396817
rect 285678 396743 285734 396752
rect 287058 396808 287114 396817
rect 287058 396743 287114 396752
rect 287704 396772 287756 396778
rect 284944 396228 284996 396234
rect 284944 396170 284996 396176
rect 283196 395344 283248 395350
rect 283196 395286 283248 395292
rect 284956 242554 284984 396170
rect 285692 244050 285720 396743
rect 287072 246770 287100 396743
rect 287704 396714 287756 396720
rect 287060 246764 287112 246770
rect 287060 246706 287112 246712
rect 287716 245410 287744 396714
rect 289832 396234 289860 397287
rect 298480 397254 298508 397287
rect 291844 397248 291896 397254
rect 291844 397190 291896 397196
rect 298468 397248 298520 397254
rect 298468 397190 298520 397196
rect 289820 396228 289872 396234
rect 289820 396170 289872 396176
rect 287704 245404 287756 245410
rect 287704 245346 287756 245352
rect 285680 244044 285732 244050
rect 285680 243986 285732 243992
rect 284944 242548 284996 242554
rect 284944 242490 284996 242496
rect 287702 230616 287758 230625
rect 287702 230551 287758 230560
rect 282182 220824 282238 220833
rect 282182 220759 282238 220768
rect 278044 193180 278096 193186
rect 278044 193122 278096 193128
rect 271144 126948 271196 126954
rect 271144 126890 271196 126896
rect 269120 59220 269172 59226
rect 269120 59162 269172 59168
rect 268384 59084 268436 59090
rect 268384 59026 268436 59032
rect 263600 58268 263652 58274
rect 263600 58210 263652 58216
rect 251180 58200 251232 58206
rect 251180 58142 251232 58148
rect 242164 56908 242216 56914
rect 242164 56850 242216 56856
rect 233240 56840 233292 56846
rect 233240 56782 233292 56788
rect 230572 56704 230624 56710
rect 230572 56646 230624 56652
rect 225052 56636 225104 56642
rect 225052 56578 225104 56584
rect 224960 55684 225012 55690
rect 224960 55626 225012 55632
rect 222844 54120 222896 54126
rect 222844 54062 222896 54068
rect 220176 24132 220228 24138
rect 220176 24074 220228 24080
rect 220084 20052 220136 20058
rect 220084 19994 220136 20000
rect 220820 18488 220872 18494
rect 220820 18430 220872 18436
rect 220832 16574 220860 18430
rect 220832 16546 221596 16574
rect 220452 15564 220504 15570
rect 220452 15506 220504 15512
rect 219256 9920 219308 9926
rect 219256 9862 219308 9868
rect 219268 480 219296 9862
rect 220464 480 220492 15506
rect 221568 480 221596 16546
rect 222752 9988 222804 9994
rect 222752 9930 222804 9936
rect 222764 480 222792 9930
rect 222856 4146 222884 54062
rect 224972 16574 225000 55626
rect 227720 55480 227772 55486
rect 227720 55422 227772 55428
rect 227732 16574 227760 55422
rect 231860 54188 231912 54194
rect 231860 54130 231912 54136
rect 229100 52760 229152 52766
rect 229100 52702 229152 52708
rect 229112 16574 229140 52702
rect 231872 16574 231900 54130
rect 258080 52964 258132 52970
rect 258080 52906 258132 52912
rect 251180 52896 251232 52902
rect 251180 52838 251232 52844
rect 233240 52828 233292 52834
rect 233240 52770 233292 52776
rect 233252 16574 233280 52770
rect 236000 51536 236052 51542
rect 236000 51478 236052 51484
rect 236012 16574 236040 51478
rect 240140 51468 240192 51474
rect 240140 51410 240192 51416
rect 238116 16584 238168 16590
rect 224972 16546 225184 16574
rect 227732 16546 228772 16574
rect 229112 16546 229876 16574
rect 231872 16546 232268 16574
rect 233252 16546 233464 16574
rect 236012 16546 237052 16574
rect 223948 15632 224000 15638
rect 223948 15574 224000 15580
rect 222844 4140 222896 4146
rect 222844 4082 222896 4088
rect 223960 480 223988 15574
rect 225156 480 225184 16546
rect 226340 15700 226392 15706
rect 226340 15642 226392 15648
rect 226352 4078 226380 15642
rect 226432 10056 226484 10062
rect 226432 9998 226484 10004
rect 226340 4072 226392 4078
rect 226340 4014 226392 4020
rect 226444 3482 226472 9998
rect 227536 4072 227588 4078
rect 227536 4014 227588 4020
rect 226352 3454 226472 3482
rect 226352 480 226380 3454
rect 227548 480 227576 4014
rect 228744 480 228772 16546
rect 229848 480 229876 16546
rect 231032 15768 231084 15774
rect 231032 15710 231084 15716
rect 231044 480 231072 15710
rect 232240 480 232268 16546
rect 233436 480 233464 16546
rect 234620 15836 234672 15842
rect 234620 15778 234672 15784
rect 234632 480 234660 15778
rect 235816 5636 235868 5642
rect 235816 5578 235868 5584
rect 235828 480 235856 5578
rect 237024 480 237052 16546
rect 240152 16574 240180 51410
rect 247040 18556 247092 18562
rect 247040 18498 247092 18504
rect 242900 17060 242952 17066
rect 242900 17002 242952 17008
rect 240152 16546 240548 16574
rect 238116 16526 238168 16532
rect 238128 480 238156 16526
rect 239312 5704 239364 5710
rect 239312 5646 239364 5652
rect 239324 480 239352 5646
rect 240520 480 240548 16546
rect 241704 16516 241756 16522
rect 241704 16458 241756 16464
rect 241716 480 241744 16458
rect 242912 3398 242940 17002
rect 247052 16574 247080 18498
rect 247052 16546 247632 16574
rect 245200 16448 245252 16454
rect 245200 16390 245252 16396
rect 242992 5772 243044 5778
rect 242992 5714 243044 5720
rect 242900 3392 242952 3398
rect 242900 3334 242952 3340
rect 243004 2938 243032 5714
rect 244096 3392 244148 3398
rect 244096 3334 244148 3340
rect 242912 2910 243032 2938
rect 242912 480 242940 2910
rect 244108 480 244136 3334
rect 245212 480 245240 16390
rect 246396 5840 246448 5846
rect 246396 5782 246448 5788
rect 246408 480 246436 5782
rect 247604 480 247632 16546
rect 248788 16380 248840 16386
rect 248788 16322 248840 16328
rect 248800 480 248828 16322
rect 249984 5908 250036 5914
rect 249984 5850 250036 5856
rect 249996 480 250024 5850
rect 251192 480 251220 52838
rect 253940 51604 253992 51610
rect 253940 51546 253992 51552
rect 253952 16574 253980 51546
rect 255320 17128 255372 17134
rect 255320 17070 255372 17076
rect 255332 16574 255360 17070
rect 258092 16574 258120 52906
rect 284300 50244 284352 50250
rect 284300 50186 284352 50192
rect 276020 48952 276072 48958
rect 276020 48894 276072 48900
rect 262220 17944 262272 17950
rect 262220 17886 262272 17892
rect 259460 17196 259512 17202
rect 259460 17138 259512 17144
rect 253952 16546 254716 16574
rect 255332 16546 255912 16574
rect 258092 16546 258304 16574
rect 252376 16312 252428 16318
rect 252376 16254 252428 16260
rect 252388 480 252416 16254
rect 253480 5976 253532 5982
rect 253480 5918 253532 5924
rect 253492 480 253520 5918
rect 254688 480 254716 16546
rect 255884 480 255912 16546
rect 257068 6044 257120 6050
rect 257068 5986 257120 5992
rect 257080 480 257108 5986
rect 258276 480 258304 16546
rect 259472 480 259500 17138
rect 262232 16574 262260 17886
rect 266360 17876 266412 17882
rect 266360 17818 266412 17824
rect 266372 16574 266400 17818
rect 269120 17808 269172 17814
rect 269120 17750 269172 17756
rect 269132 16574 269160 17750
rect 273260 17740 273312 17746
rect 273260 17682 273312 17688
rect 273272 16574 273300 17682
rect 262232 16546 262996 16574
rect 266372 16546 266584 16574
rect 269132 16546 270080 16574
rect 273272 16546 273668 16574
rect 261760 11212 261812 11218
rect 261760 11154 261812 11160
rect 260656 6112 260708 6118
rect 260656 6054 260708 6060
rect 260668 480 260696 6054
rect 261772 480 261800 11154
rect 262968 480 262996 16546
rect 265348 11280 265400 11286
rect 265348 11222 265400 11228
rect 264152 6860 264204 6866
rect 264152 6802 264204 6808
rect 264164 480 264192 6802
rect 265360 480 265388 11222
rect 266556 480 266584 16546
rect 268844 11348 268896 11354
rect 268844 11290 268896 11296
rect 267740 6792 267792 6798
rect 267740 6734 267792 6740
rect 267752 480 267780 6734
rect 268856 480 268884 11290
rect 270052 480 270080 16546
rect 272432 11416 272484 11422
rect 272432 11358 272484 11364
rect 271236 6724 271288 6730
rect 271236 6666 271288 6672
rect 271248 480 271276 6666
rect 272444 480 272472 11358
rect 273640 480 273668 16546
rect 274824 6656 274876 6662
rect 274824 6598 274876 6604
rect 274836 480 274864 6598
rect 276032 4146 276060 48894
rect 280160 17672 280212 17678
rect 280160 17614 280212 17620
rect 280172 16574 280200 17614
rect 280172 16546 280752 16574
rect 279516 11552 279568 11558
rect 279516 11494 279568 11500
rect 276112 11484 276164 11490
rect 276112 11426 276164 11432
rect 276020 4140 276072 4146
rect 276020 4082 276072 4088
rect 276124 3482 276152 11426
rect 278320 6588 278372 6594
rect 278320 6530 278372 6536
rect 277124 4140 277176 4146
rect 277124 4082 277176 4088
rect 276032 3454 276152 3482
rect 276032 480 276060 3454
rect 277136 480 277164 4082
rect 278332 480 278360 6530
rect 279528 480 279556 11494
rect 280724 480 280752 16546
rect 283104 11620 283156 11626
rect 283104 11562 283156 11568
rect 281908 6520 281960 6526
rect 281908 6462 281960 6468
rect 281920 480 281948 6462
rect 283116 480 283144 11562
rect 284312 480 284340 50186
rect 287716 46918 287744 230551
rect 291856 59702 291884 397190
rect 292946 396808 293002 396817
rect 292946 396743 293002 396752
rect 295890 396808 295946 396817
rect 295890 396743 295892 396752
rect 292960 396710 292988 396743
rect 295944 396743 295946 396752
rect 295892 396714 295944 396720
rect 291936 396704 291988 396710
rect 291936 396646 291988 396652
rect 292948 396704 293000 396710
rect 292948 396646 293000 396652
rect 291948 244186 291976 396646
rect 291936 244180 291988 244186
rect 291936 244122 291988 244128
rect 295982 226536 296038 226545
rect 295982 226471 296038 226480
rect 295996 60722 296024 226471
rect 300136 187649 300164 398103
rect 302238 396808 302294 396817
rect 302238 396743 302294 396752
rect 305274 396808 305330 396817
rect 307850 396808 307906 396817
rect 305274 396743 305330 396752
rect 307024 396772 307076 396778
rect 302252 244118 302280 396743
rect 305288 396710 305316 396743
rect 307850 396743 307852 396752
rect 307024 396714 307076 396720
rect 307904 396743 307906 396752
rect 310518 396808 310574 396817
rect 310518 396743 310574 396752
rect 313278 396808 313334 396817
rect 313278 396743 313334 396752
rect 307852 396714 307904 396720
rect 304264 396704 304316 396710
rect 304264 396646 304316 396652
rect 305276 396704 305328 396710
rect 305276 396646 305328 396652
rect 302240 244112 302292 244118
rect 302240 244054 302292 244060
rect 302882 227760 302938 227769
rect 302882 227695 302938 227704
rect 300122 187640 300178 187649
rect 300122 187575 300178 187584
rect 302896 100706 302924 227695
rect 302884 100700 302936 100706
rect 302884 100642 302936 100648
rect 295984 60716 296036 60722
rect 295984 60658 296036 60664
rect 291844 59696 291896 59702
rect 291844 59638 291896 59644
rect 304276 59634 304304 396646
rect 307036 201385 307064 396714
rect 309784 396704 309836 396710
rect 309784 396646 309836 396652
rect 307022 201376 307078 201385
rect 307022 201311 307078 201320
rect 304264 59628 304316 59634
rect 304264 59570 304316 59576
rect 309796 59566 309824 396646
rect 310532 247790 310560 396743
rect 310520 247784 310572 247790
rect 310520 247726 310572 247732
rect 309784 59560 309836 59566
rect 309784 59502 309836 59508
rect 313292 59498 313320 396743
rect 315776 396710 315804 398103
rect 317418 396808 317474 396817
rect 317418 396743 317474 396752
rect 320178 396808 320234 396817
rect 320178 396743 320234 396752
rect 323122 396808 323178 396817
rect 323122 396743 323178 396752
rect 315764 396704 315816 396710
rect 315764 396646 315816 396652
rect 316684 396160 316736 396166
rect 316684 396102 316736 396108
rect 316696 248130 316724 396102
rect 317432 250510 317460 396743
rect 317420 250504 317472 250510
rect 317420 250446 317472 250452
rect 316684 248124 316736 248130
rect 316684 248066 316736 248072
rect 320192 242486 320220 396743
rect 323136 396710 323164 396743
rect 322204 396704 322256 396710
rect 322204 396646 322256 396652
rect 323124 396704 323176 396710
rect 323124 396646 323176 396652
rect 320180 242480 320232 242486
rect 320180 242422 320232 242428
rect 313280 59492 313332 59498
rect 313280 59434 313332 59440
rect 322216 59430 322244 396646
rect 325896 396302 325924 398103
rect 343362 397352 343418 397361
rect 343362 397287 343418 397296
rect 342350 396808 342406 396817
rect 342350 396743 342406 396752
rect 325884 396296 325936 396302
rect 325884 396238 325936 396244
rect 342364 247994 342392 396743
rect 343376 396166 343404 397287
rect 343364 396160 343416 396166
rect 343364 396102 343416 396108
rect 342352 247988 342404 247994
rect 342352 247930 342404 247936
rect 322204 59424 322256 59430
rect 322204 59366 322256 59372
rect 356532 57225 356560 470566
rect 357452 60353 357480 479159
rect 358084 456816 358136 456822
rect 358084 456758 358136 456764
rect 357622 415848 357678 415857
rect 357622 415783 357678 415792
rect 357530 413128 357586 413137
rect 357530 413063 357586 413072
rect 357544 245342 357572 413063
rect 357636 399566 357664 415783
rect 357624 399560 357676 399566
rect 357624 399502 357676 399508
rect 357532 245336 357584 245342
rect 357532 245278 357584 245284
rect 358096 242282 358124 456758
rect 358818 418840 358874 418849
rect 358818 418775 358874 418784
rect 358084 242276 358136 242282
rect 358084 242218 358136 242224
rect 357438 60344 357494 60353
rect 357438 60279 357494 60288
rect 358832 59265 358860 418775
rect 358910 417208 358966 417217
rect 358910 417143 358966 417152
rect 358818 59256 358874 59265
rect 358818 59191 358874 59200
rect 358924 58682 358952 417143
rect 359002 414352 359058 414361
rect 359002 414287 359058 414296
rect 359016 399498 359044 414287
rect 359004 399492 359056 399498
rect 359004 399434 359056 399440
rect 360856 258806 360884 699654
rect 371884 696992 371936 696998
rect 371884 696934 371936 696940
rect 370504 643136 370556 643142
rect 370504 643078 370556 643084
rect 367744 590708 367796 590714
rect 367744 590650 367796 590656
rect 363604 484424 363656 484430
rect 363604 484366 363656 484372
rect 360844 258800 360896 258806
rect 360844 258742 360896 258748
rect 363616 243846 363644 484366
rect 367756 243914 367784 590650
rect 370516 245070 370544 643078
rect 370504 245064 370556 245070
rect 370504 245006 370556 245012
rect 371896 243982 371924 696934
rect 374656 245138 374684 700334
rect 376036 258738 376064 700470
rect 376024 258732 376076 258738
rect 376024 258674 376076 258680
rect 377416 245206 377444 700538
rect 388444 700460 388496 700466
rect 388444 700402 388496 700408
rect 385684 683188 385736 683194
rect 385684 683130 385736 683136
rect 382924 630692 382976 630698
rect 382924 630634 382976 630640
rect 381544 524476 381596 524482
rect 381544 524418 381596 524424
rect 378784 430636 378836 430642
rect 378784 430578 378836 430584
rect 378796 246498 378824 430578
rect 378784 246492 378836 246498
rect 378784 246434 378836 246440
rect 377404 245200 377456 245206
rect 377404 245142 377456 245148
rect 374644 245132 374696 245138
rect 374644 245074 374696 245080
rect 381556 245002 381584 524418
rect 382936 246634 382964 630634
rect 382924 246628 382976 246634
rect 382924 246570 382976 246576
rect 385696 246566 385724 683130
rect 388456 246702 388484 700402
rect 388444 246696 388496 246702
rect 388444 246638 388496 246644
rect 385684 246560 385736 246566
rect 385684 246502 385736 246508
rect 412652 246430 412680 703582
rect 413480 703474 413508 703582
rect 413622 703520 413734 704960
rect 429212 703582 429700 703610
rect 413664 703474 413692 703520
rect 413480 703446 413692 703474
rect 425704 404388 425756 404394
rect 425704 404330 425756 404336
rect 412640 246424 412692 246430
rect 412640 246366 412692 246372
rect 381544 244996 381596 245002
rect 381544 244938 381596 244944
rect 371884 243976 371936 243982
rect 371884 243918 371936 243924
rect 367744 243908 367796 243914
rect 367744 243850 367796 243856
rect 363604 243840 363656 243846
rect 363604 243782 363656 243788
rect 425716 243642 425744 404330
rect 429212 243778 429240 703582
rect 429672 703474 429700 703582
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 429856 703474 429884 703520
rect 429672 703446 429884 703474
rect 446404 700596 446456 700602
rect 446404 700538 446456 700544
rect 431224 536852 431276 536858
rect 431224 536794 431276 536800
rect 429200 243772 429252 243778
rect 429200 243714 429252 243720
rect 431236 243710 431264 536794
rect 443644 470620 443696 470626
rect 443644 470562 443696 470568
rect 443656 244934 443684 470562
rect 443644 244928 443696 244934
rect 443644 244870 443696 244876
rect 431224 243704 431276 243710
rect 431224 243646 431276 243652
rect 425704 243636 425756 243642
rect 425704 243578 425756 243584
rect 446416 242214 446444 700538
rect 462332 700534 462360 703520
rect 462320 700528 462372 700534
rect 462320 700470 462372 700476
rect 478524 700466 478552 703520
rect 494808 700602 494836 703520
rect 494796 700596 494848 700602
rect 494796 700538 494848 700544
rect 478512 700460 478564 700466
rect 478512 700402 478564 700408
rect 527192 700398 527220 703520
rect 543476 702434 543504 703520
rect 542372 702406 543504 702434
rect 527180 700392 527232 700398
rect 527180 700334 527232 700340
rect 449164 576904 449216 576910
rect 449164 576846 449216 576852
rect 449176 243574 449204 576846
rect 542372 246362 542400 702406
rect 559668 700330 559696 703520
rect 559656 700324 559708 700330
rect 559656 700266 559708 700272
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683194 580212 683839
rect 580172 683188 580224 683194
rect 580172 683130 580224 683136
rect 580172 670744 580224 670750
rect 580170 670712 580172 670721
rect 580224 670712 580226 670721
rect 580170 670647 580226 670656
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 580170 630864 580226 630873
rect 580170 630799 580226 630808
rect 580184 630698 580212 630799
rect 580172 630692 580224 630698
rect 580172 630634 580224 630640
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616894 580212 617471
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 579802 591016 579858 591025
rect 579802 590951 579858 590960
rect 579816 590714 579844 590951
rect 579804 590708 579856 590714
rect 579804 590650 579856 590656
rect 580170 577688 580226 577697
rect 580170 577623 580226 577632
rect 580184 576910 580212 577623
rect 580172 576904 580224 576910
rect 580172 576846 580224 576852
rect 579802 564360 579858 564369
rect 579802 564295 579858 564304
rect 579816 563106 579844 564295
rect 579804 563100 579856 563106
rect 579804 563042 579856 563048
rect 580170 537840 580226 537849
rect 580170 537775 580226 537784
rect 580184 536858 580212 537775
rect 580172 536852 580224 536858
rect 580172 536794 580224 536800
rect 580170 524512 580226 524521
rect 580170 524447 580172 524456
rect 580224 524447 580226 524456
rect 580172 524418 580224 524424
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 580184 510678 580212 511255
rect 580172 510672 580224 510678
rect 580172 510614 580224 510620
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 580184 484430 580212 484599
rect 580172 484424 580224 484430
rect 580172 484366 580224 484372
rect 579986 471472 580042 471481
rect 579986 471407 580042 471416
rect 580000 470626 580028 471407
rect 579988 470620 580040 470626
rect 579988 470562 580040 470568
rect 580170 458144 580226 458153
rect 580170 458079 580226 458088
rect 580184 456822 580212 458079
rect 580172 456816 580224 456822
rect 580172 456758 580224 456764
rect 580170 431624 580226 431633
rect 580170 431559 580226 431568
rect 580184 430642 580212 431559
rect 580172 430636 580224 430642
rect 580172 430578 580224 430584
rect 580262 418296 580318 418305
rect 580262 418231 580318 418240
rect 580170 404968 580226 404977
rect 580170 404903 580226 404912
rect 580184 404394 580212 404903
rect 580172 404388 580224 404394
rect 580172 404330 580224 404336
rect 580170 378448 580226 378457
rect 580170 378383 580226 378392
rect 580184 378214 580212 378383
rect 580172 378208 580224 378214
rect 580172 378150 580224 378156
rect 579618 365120 579674 365129
rect 579618 365055 579674 365064
rect 579632 364410 579660 365055
rect 579620 364404 579672 364410
rect 579620 364346 579672 364352
rect 580172 351960 580224 351966
rect 580170 351928 580172 351937
rect 580224 351928 580226 351937
rect 580170 351863 580226 351872
rect 580170 325272 580226 325281
rect 580170 325207 580226 325216
rect 580184 324358 580212 325207
rect 580172 324352 580224 324358
rect 580172 324294 580224 324300
rect 579986 312080 580042 312089
rect 579986 312015 580042 312024
rect 580000 311914 580028 312015
rect 579988 311908 580040 311914
rect 579988 311850 580040 311856
rect 580170 298752 580226 298761
rect 580170 298687 580226 298696
rect 580184 298178 580212 298687
rect 580172 298172 580224 298178
rect 580172 298114 580224 298120
rect 580170 272232 580226 272241
rect 580170 272167 580226 272176
rect 580184 271930 580212 272167
rect 580172 271924 580224 271930
rect 580172 271866 580224 271872
rect 580170 258904 580226 258913
rect 580170 258839 580226 258848
rect 580184 258126 580212 258839
rect 580172 258120 580224 258126
rect 580172 258062 580224 258068
rect 580276 247722 580304 418231
rect 580264 247716 580316 247722
rect 580264 247658 580316 247664
rect 542360 246356 542412 246362
rect 542360 246298 542412 246304
rect 579802 245576 579858 245585
rect 579802 245511 579858 245520
rect 579816 244322 579844 245511
rect 579804 244316 579856 244322
rect 579804 244258 579856 244264
rect 449164 243568 449216 243574
rect 449164 243510 449216 243516
rect 446404 242208 446456 242214
rect 446404 242150 446456 242156
rect 580262 229120 580318 229129
rect 580262 229055 580318 229064
rect 410522 226400 410578 226409
rect 410522 226335 410578 226344
rect 410536 139398 410564 226335
rect 580172 206984 580224 206990
rect 580172 206926 580224 206932
rect 580184 205737 580212 206926
rect 580170 205728 580226 205737
rect 580170 205663 580226 205672
rect 580172 193180 580224 193186
rect 580172 193122 580224 193128
rect 580184 192545 580212 193122
rect 580170 192536 580226 192545
rect 580170 192471 580226 192480
rect 580172 167000 580224 167006
rect 580172 166942 580224 166948
rect 580184 165889 580212 166942
rect 580170 165880 580226 165889
rect 580170 165815 580226 165824
rect 410524 139392 410576 139398
rect 580172 139392 580224 139398
rect 410524 139334 410576 139340
rect 580170 139360 580172 139369
rect 580224 139360 580226 139369
rect 580170 139295 580226 139304
rect 580172 126948 580224 126954
rect 580172 126890 580224 126896
rect 580184 126041 580212 126890
rect 580170 126032 580226 126041
rect 580170 125967 580226 125976
rect 580172 100700 580224 100706
rect 580172 100642 580224 100648
rect 580184 99521 580212 100642
rect 580170 99512 580226 99521
rect 580170 99447 580226 99456
rect 580276 86193 580304 229055
rect 580262 86184 580318 86193
rect 580262 86119 580318 86128
rect 580172 60716 580224 60722
rect 580172 60658 580224 60664
rect 580184 59673 580212 60658
rect 580170 59664 580226 59673
rect 580170 59599 580226 59608
rect 358912 58676 358964 58682
rect 358912 58618 358964 58624
rect 391204 57384 391256 57390
rect 391204 57326 391256 57332
rect 382924 57316 382976 57322
rect 382924 57258 382976 57264
rect 356518 57216 356574 57225
rect 356518 57151 356574 57160
rect 316040 55208 316092 55214
rect 316040 55150 316092 55156
rect 313280 54460 313332 54466
rect 313280 54402 313332 54408
rect 309140 54392 309192 54398
rect 309140 54334 309192 54340
rect 306380 54324 306432 54330
rect 306380 54266 306432 54272
rect 302240 54256 302292 54262
rect 302240 54198 302292 54204
rect 291200 49700 291252 49706
rect 291200 49642 291252 49648
rect 287704 46912 287756 46918
rect 287704 46854 287756 46860
rect 287060 19304 287112 19310
rect 287060 19246 287112 19252
rect 287072 16574 287100 19246
rect 291212 16574 291240 49642
rect 298100 49632 298152 49638
rect 298100 49574 298152 49580
rect 293960 49564 294012 49570
rect 293960 49506 294012 49512
rect 293972 16574 294000 49506
rect 298112 16574 298140 49574
rect 300860 17468 300912 17474
rect 300860 17410 300912 17416
rect 300872 16574 300900 17410
rect 302252 16574 302280 54198
rect 305000 49428 305052 49434
rect 305000 49370 305052 49376
rect 305012 16574 305040 49370
rect 306392 16574 306420 54266
rect 307760 17400 307812 17406
rect 307760 17342 307812 17348
rect 287072 16546 287836 16574
rect 291212 16546 291424 16574
rect 293972 16546 294920 16574
rect 298112 16546 298508 16574
rect 300872 16546 302004 16574
rect 302252 16546 303200 16574
rect 305012 16546 305592 16574
rect 306392 16546 306788 16574
rect 286600 11688 286652 11694
rect 286600 11630 286652 11636
rect 285404 6452 285456 6458
rect 285404 6394 285456 6400
rect 285416 480 285444 6394
rect 286612 480 286640 11630
rect 287808 480 287836 16546
rect 290188 12436 290240 12442
rect 290188 12378 290240 12384
rect 288992 6384 289044 6390
rect 288992 6326 289044 6332
rect 289004 480 289032 6326
rect 290200 480 290228 12378
rect 291396 480 291424 16546
rect 293684 12368 293736 12374
rect 293684 12310 293736 12316
rect 292580 6316 292632 6322
rect 292580 6258 292632 6264
rect 292592 480 292620 6258
rect 293696 480 293724 12310
rect 294892 480 294920 16546
rect 297272 12300 297324 12306
rect 297272 12242 297324 12248
rect 296076 6248 296128 6254
rect 296076 6190 296128 6196
rect 296088 480 296116 6190
rect 297284 480 297312 12242
rect 298480 480 298508 16546
rect 299480 12232 299532 12238
rect 299480 12174 299532 12180
rect 299492 1698 299520 12174
rect 299664 6180 299716 6186
rect 299664 6122 299716 6128
rect 299480 1692 299532 1698
rect 299480 1634 299532 1640
rect 299676 480 299704 6122
rect 300768 1692 300820 1698
rect 300768 1634 300820 1640
rect 300780 480 300808 1634
rect 301976 480 302004 16546
rect 303172 480 303200 16546
rect 304356 12164 304408 12170
rect 304356 12106 304408 12112
rect 304368 480 304396 12106
rect 305564 480 305592 16546
rect 306760 480 306788 16546
rect 307772 3398 307800 17342
rect 309152 16574 309180 54334
rect 311900 49496 311952 49502
rect 311900 49438 311952 49444
rect 311912 16574 311940 49438
rect 313292 16574 313320 54402
rect 309152 16546 310284 16574
rect 311912 16546 312676 16574
rect 313292 16546 313872 16574
rect 307944 12096 307996 12102
rect 307944 12038 307996 12044
rect 307760 3392 307812 3398
rect 307760 3334 307812 3340
rect 307956 480 307984 12038
rect 309048 3392 309100 3398
rect 309048 3334 309100 3340
rect 309060 480 309088 3334
rect 310256 480 310284 16546
rect 311440 12028 311492 12034
rect 311440 11970 311492 11976
rect 311452 480 311480 11970
rect 312648 480 312676 16546
rect 313844 480 313872 16546
rect 315028 11960 315080 11966
rect 315028 11902 315080 11908
rect 315040 480 315068 11902
rect 316052 3398 316080 55150
rect 320180 55140 320232 55146
rect 320180 55082 320232 55088
rect 316132 49224 316184 49230
rect 316132 49166 316184 49172
rect 316144 16574 316172 49166
rect 318800 17604 318852 17610
rect 318800 17546 318852 17552
rect 318812 16574 318840 17546
rect 320192 16574 320220 55082
rect 324320 55072 324372 55078
rect 324320 55014 324372 55020
rect 322940 50312 322992 50318
rect 322940 50254 322992 50260
rect 322952 16574 322980 50254
rect 324332 16574 324360 55014
rect 327080 55004 327132 55010
rect 327080 54946 327132 54952
rect 325700 17536 325752 17542
rect 325700 17478 325752 17484
rect 325712 16574 325740 17478
rect 327092 16574 327120 54946
rect 353300 53780 353352 53786
rect 353300 53722 353352 53728
rect 331220 53032 331272 53038
rect 331220 52974 331272 52980
rect 328460 51672 328512 51678
rect 328460 51614 328512 51620
rect 328472 16574 328500 51614
rect 329840 49292 329892 49298
rect 329840 49234 329892 49240
rect 329852 16574 329880 49234
rect 331232 16574 331260 52974
rect 335360 52420 335412 52426
rect 335360 52362 335412 52368
rect 332600 19100 332652 19106
rect 332600 19042 332652 19048
rect 316144 16546 316264 16574
rect 318812 16546 319760 16574
rect 320192 16546 320956 16574
rect 322952 16546 323348 16574
rect 324332 16546 324452 16574
rect 325712 16546 326844 16574
rect 327092 16546 328040 16574
rect 328472 16546 329236 16574
rect 329852 16546 330432 16574
rect 331232 16546 331628 16574
rect 316040 3392 316092 3398
rect 316040 3334 316092 3340
rect 316236 480 316264 16546
rect 318524 11892 318576 11898
rect 318524 11834 318576 11840
rect 317328 3392 317380 3398
rect 317328 3334 317380 3340
rect 317340 480 317368 3334
rect 318536 480 318564 11834
rect 319732 480 319760 16546
rect 320928 480 320956 16546
rect 322112 11824 322164 11830
rect 322112 11766 322164 11772
rect 322124 480 322152 11766
rect 323320 480 323348 16546
rect 324424 480 324452 16546
rect 325608 11756 325660 11762
rect 325608 11698 325660 11704
rect 325620 480 325648 11698
rect 326816 480 326844 16546
rect 328012 480 328040 16546
rect 329208 480 329236 16546
rect 330404 480 330432 16546
rect 331600 480 331628 16546
rect 332612 3398 332640 19042
rect 332692 17332 332744 17338
rect 332692 17274 332744 17280
rect 332600 3392 332652 3398
rect 332600 3334 332652 3340
rect 332704 480 332732 17274
rect 335372 16574 335400 52362
rect 339500 52352 339552 52358
rect 339500 52294 339552 52300
rect 336740 19168 336792 19174
rect 336740 19110 336792 19116
rect 336752 16574 336780 19110
rect 339512 16574 339540 52294
rect 342260 52284 342312 52290
rect 342260 52226 342312 52232
rect 340880 49360 340932 49366
rect 340880 49302 340932 49308
rect 340892 16574 340920 49302
rect 342272 16574 342300 52226
rect 346400 52216 346452 52222
rect 346400 52158 346452 52164
rect 343640 19032 343692 19038
rect 343640 18974 343692 18980
rect 343652 16574 343680 18974
rect 346412 16574 346440 52158
rect 349160 52148 349212 52154
rect 349160 52090 349212 52096
rect 347780 18964 347832 18970
rect 347780 18906 347832 18912
rect 347792 16574 347820 18906
rect 335372 16546 336320 16574
rect 336752 16546 337516 16574
rect 339512 16546 339908 16574
rect 340892 16546 341012 16574
rect 342272 16546 343404 16574
rect 343652 16546 344600 16574
rect 346412 16546 346992 16574
rect 347792 16546 348096 16574
rect 335084 7064 335136 7070
rect 335084 7006 335136 7012
rect 333888 3392 333940 3398
rect 333888 3334 333940 3340
rect 333900 480 333928 3334
rect 335096 480 335124 7006
rect 336292 480 336320 16546
rect 337488 480 337516 16546
rect 338672 7132 338724 7138
rect 338672 7074 338724 7080
rect 338684 480 338712 7074
rect 339880 480 339908 16546
rect 340984 480 341012 16546
rect 342168 7200 342220 7206
rect 342168 7142 342220 7148
rect 342180 480 342208 7142
rect 343376 480 343404 16546
rect 344572 480 344600 16546
rect 345756 7268 345808 7274
rect 345756 7210 345808 7216
rect 345768 480 345796 7210
rect 346964 480 346992 16546
rect 348068 480 348096 16546
rect 349172 3398 349200 52090
rect 350540 18896 350592 18902
rect 350540 18838 350592 18844
rect 350552 16574 350580 18838
rect 353312 16574 353340 53722
rect 357440 52080 357492 52086
rect 357440 52022 357492 52028
rect 354680 18828 354732 18834
rect 354680 18770 354732 18776
rect 354692 16574 354720 18770
rect 350552 16546 351684 16574
rect 353312 16546 354076 16574
rect 354692 16546 355272 16574
rect 349252 7336 349304 7342
rect 349252 7278 349304 7284
rect 349160 3392 349212 3398
rect 349160 3334 349212 3340
rect 349264 480 349292 7278
rect 350448 3392 350500 3398
rect 350448 3334 350500 3340
rect 350460 480 350488 3334
rect 351656 480 351684 16546
rect 352840 7404 352892 7410
rect 352840 7346 352892 7352
rect 352852 480 352880 7346
rect 354048 480 354076 16546
rect 355244 480 355272 16546
rect 356336 7472 356388 7478
rect 356336 7414 356388 7420
rect 356348 480 356376 7414
rect 357452 6914 357480 52022
rect 375380 49156 375432 49162
rect 375380 49098 375432 49104
rect 357532 20256 357584 20262
rect 357532 20198 357584 20204
rect 357544 11762 357572 20198
rect 365720 19236 365772 19242
rect 365720 19178 365772 19184
rect 361580 18760 361632 18766
rect 361580 18702 361632 18708
rect 361592 16574 361620 18702
rect 365732 16574 365760 19178
rect 368480 18692 368532 18698
rect 368480 18634 368532 18640
rect 368492 16574 368520 18634
rect 375392 16574 375420 49098
rect 382280 49088 382332 49094
rect 382280 49030 382332 49036
rect 361592 16546 362356 16574
rect 365732 16546 365852 16574
rect 368492 16546 369440 16574
rect 375392 16546 376524 16574
rect 361120 12572 361172 12578
rect 361120 12514 361172 12520
rect 357532 11756 357584 11762
rect 357532 11698 357584 11704
rect 358728 11756 358780 11762
rect 358728 11698 358780 11704
rect 357452 6886 357572 6914
rect 357544 480 357572 6886
rect 358740 480 358768 11698
rect 359924 7540 359976 7546
rect 359924 7482 359976 7488
rect 359936 480 359964 7482
rect 361132 480 361160 12514
rect 362328 480 362356 16546
rect 364616 12640 364668 12646
rect 364616 12582 364668 12588
rect 363512 8288 363564 8294
rect 363512 8230 363564 8236
rect 363524 480 363552 8230
rect 364628 480 364656 12582
rect 365824 480 365852 16546
rect 368204 12708 368256 12714
rect 368204 12650 368256 12656
rect 367008 8220 367060 8226
rect 367008 8162 367060 8168
rect 367020 480 367048 8162
rect 368216 480 368244 12650
rect 369412 480 369440 16546
rect 374000 12844 374052 12850
rect 374000 12786 374052 12792
rect 371700 12776 371752 12782
rect 371700 12718 371752 12724
rect 370596 8152 370648 8158
rect 370596 8094 370648 8100
rect 370608 480 370636 8094
rect 371712 480 371740 12718
rect 372896 10124 372948 10130
rect 372896 10066 372948 10072
rect 372908 480 372936 10066
rect 374012 3398 374040 12786
rect 374092 8084 374144 8090
rect 374092 8026 374144 8032
rect 374000 3392 374052 3398
rect 374000 3334 374052 3340
rect 374104 480 374132 8026
rect 375288 3392 375340 3398
rect 375288 3334 375340 3340
rect 375300 480 375328 3334
rect 376496 480 376524 16546
rect 378876 12912 378928 12918
rect 378876 12854 378928 12860
rect 377680 8016 377732 8022
rect 377680 7958 377732 7964
rect 377692 480 377720 7958
rect 378888 480 378916 12854
rect 381176 7948 381228 7954
rect 381176 7890 381228 7896
rect 379980 4072 380032 4078
rect 379980 4014 380032 4020
rect 379992 480 380020 4014
rect 381188 480 381216 7890
rect 382292 3330 382320 49030
rect 382372 12980 382424 12986
rect 382372 12922 382424 12928
rect 382280 3324 382332 3330
rect 382280 3266 382332 3272
rect 382384 480 382412 12922
rect 382936 3398 382964 57258
rect 387064 57248 387116 57254
rect 387064 57190 387116 57196
rect 386420 20120 386472 20126
rect 386420 20062 386472 20068
rect 386432 16574 386460 20062
rect 386432 16546 387012 16574
rect 385960 13048 386012 13054
rect 385960 12990 386012 12996
rect 384764 7880 384816 7886
rect 384764 7822 384816 7828
rect 382924 3392 382976 3398
rect 382924 3334 382976 3340
rect 383568 3324 383620 3330
rect 383568 3266 383620 3272
rect 383580 480 383608 3266
rect 384776 480 384804 7822
rect 385972 480 386000 12990
rect 386984 3482 387012 16546
rect 387076 4146 387104 57190
rect 388444 48000 388496 48006
rect 388444 47942 388496 47948
rect 388260 7812 388312 7818
rect 388260 7754 388312 7760
rect 387064 4140 387116 4146
rect 387064 4082 387116 4088
rect 386984 3454 387196 3482
rect 387168 480 387196 3454
rect 388272 480 388300 7754
rect 388456 3262 388484 47942
rect 389456 13796 389508 13802
rect 389456 13738 389508 13744
rect 388444 3256 388496 3262
rect 388444 3198 388496 3204
rect 389468 480 389496 13738
rect 391216 4078 391244 57326
rect 436744 56568 436796 56574
rect 436744 56510 436796 56516
rect 425704 55820 425756 55826
rect 425704 55762 425756 55768
rect 407764 55752 407816 55758
rect 407764 55694 407816 55700
rect 405740 54936 405792 54942
rect 405740 54878 405792 54884
rect 393320 51060 393372 51066
rect 393320 51002 393372 51008
rect 393332 16574 393360 51002
rect 396724 49020 396776 49026
rect 396724 48962 396776 48968
rect 393332 16546 394280 16574
rect 393044 13728 393096 13734
rect 393044 13670 393096 13676
rect 391848 7744 391900 7750
rect 391848 7686 391900 7692
rect 391204 4072 391256 4078
rect 391204 4014 391256 4020
rect 390652 3256 390704 3262
rect 390652 3198 390704 3204
rect 390664 480 390692 3198
rect 391860 480 391888 7686
rect 393056 480 393084 13670
rect 394252 480 394280 16546
rect 396540 13660 396592 13666
rect 396540 13602 396592 13608
rect 395344 7676 395396 7682
rect 395344 7618 395396 7624
rect 395356 480 395384 7618
rect 396552 480 396580 13602
rect 396736 3194 396764 48962
rect 400220 47864 400272 47870
rect 400220 47806 400272 47812
rect 400232 16574 400260 47806
rect 404360 20188 404412 20194
rect 404360 20130 404412 20136
rect 401600 18624 401652 18630
rect 401600 18566 401652 18572
rect 401612 16574 401640 18566
rect 404372 16574 404400 20130
rect 405752 16574 405780 54878
rect 407120 47796 407172 47802
rect 407120 47738 407172 47744
rect 400232 16546 401364 16574
rect 401612 16546 402560 16574
rect 404372 16546 404860 16574
rect 405752 16546 406056 16574
rect 398840 13592 398892 13598
rect 398840 13534 398892 13540
rect 398852 3330 398880 13534
rect 398932 7608 398984 7614
rect 398932 7550 398984 7556
rect 398840 3324 398892 3330
rect 398840 3266 398892 3272
rect 396724 3188 396776 3194
rect 396724 3130 396776 3136
rect 397736 3188 397788 3194
rect 397736 3130 397788 3136
rect 397748 480 397776 3130
rect 398944 480 398972 7550
rect 400128 3324 400180 3330
rect 400128 3266 400180 3272
rect 400140 480 400168 3266
rect 401336 480 401364 16546
rect 402532 480 402560 16546
rect 403624 13524 403676 13530
rect 403624 13466 403676 13472
rect 403636 480 403664 13466
rect 404832 480 404860 16546
rect 406028 480 406056 16546
rect 407132 3262 407160 47738
rect 407212 13456 407264 13462
rect 407212 13398 407264 13404
rect 407120 3256 407172 3262
rect 407120 3198 407172 3204
rect 407224 480 407252 13398
rect 407776 3330 407804 55694
rect 412640 54868 412692 54874
rect 412640 54810 412692 54816
rect 411260 47932 411312 47938
rect 411260 47874 411312 47880
rect 411272 16574 411300 47874
rect 412652 16574 412680 54810
rect 414664 54800 414716 54806
rect 414664 54742 414716 54748
rect 411272 16546 411944 16574
rect 412652 16546 413140 16574
rect 410800 13388 410852 13394
rect 410800 13330 410852 13336
rect 407764 3324 407816 3330
rect 407764 3266 407816 3272
rect 409604 3324 409656 3330
rect 409604 3266 409656 3272
rect 408408 3256 408460 3262
rect 408408 3198 408460 3204
rect 408420 480 408448 3198
rect 409616 480 409644 3266
rect 410812 480 410840 13330
rect 411916 480 411944 16546
rect 413112 480 413140 16546
rect 414296 13320 414348 13326
rect 414296 13262 414348 13268
rect 414308 480 414336 13262
rect 414676 3330 414704 54742
rect 418804 53712 418856 53718
rect 418804 53654 418856 53660
rect 418160 47592 418212 47598
rect 418160 47534 418212 47540
rect 415492 17264 415544 17270
rect 415492 17206 415544 17212
rect 414664 3324 414716 3330
rect 414664 3266 414716 3272
rect 415504 480 415532 17206
rect 418172 16574 418200 47534
rect 418172 16546 418752 16574
rect 417884 13252 417936 13258
rect 417884 13194 417936 13200
rect 416688 3324 416740 3330
rect 416688 3266 416740 3272
rect 416700 480 416728 3266
rect 417896 480 417924 13194
rect 418724 3074 418752 16546
rect 418816 3262 418844 53654
rect 421564 53644 421616 53650
rect 421564 53586 421616 53592
rect 421380 13184 421432 13190
rect 421380 13126 421432 13132
rect 418804 3256 418856 3262
rect 418804 3198 418856 3204
rect 420184 3256 420236 3262
rect 420184 3198 420236 3204
rect 418724 3046 419028 3074
rect 419000 480 419028 3046
rect 420196 480 420224 3198
rect 421392 480 421420 13126
rect 421576 2922 421604 53586
rect 425060 20052 425112 20058
rect 425060 19994 425112 20000
rect 422300 19984 422352 19990
rect 422300 19926 422352 19932
rect 422312 16574 422340 19926
rect 422312 16546 422616 16574
rect 421564 2916 421616 2922
rect 421564 2858 421616 2864
rect 422588 480 422616 16546
rect 423772 13116 423824 13122
rect 423772 13058 423824 13064
rect 423784 3330 423812 13058
rect 425072 6914 425100 19994
rect 425716 16574 425744 55762
rect 427820 54732 427872 54738
rect 427820 54674 427872 54680
rect 427832 16574 427860 54674
rect 430580 53508 430632 53514
rect 430580 53450 430632 53456
rect 430592 16574 430620 53450
rect 431960 52012 432012 52018
rect 431960 51954 432012 51960
rect 425716 16546 425836 16574
rect 427832 16546 428504 16574
rect 430592 16546 430896 16574
rect 425072 6886 425744 6914
rect 423772 3324 423824 3330
rect 423772 3266 423824 3272
rect 424968 3324 425020 3330
rect 424968 3266 425020 3272
rect 423772 2916 423824 2922
rect 423772 2858 423824 2864
rect 423784 480 423812 2858
rect 424980 480 425008 3266
rect 425716 2938 425744 6886
rect 425808 3058 425836 16546
rect 425796 3052 425848 3058
rect 425796 2994 425848 3000
rect 427268 3052 427320 3058
rect 427268 2994 427320 3000
rect 425716 2910 426204 2938
rect 426176 480 426204 2910
rect 427280 480 427308 2994
rect 428476 480 428504 16546
rect 429660 4004 429712 4010
rect 429660 3946 429712 3952
rect 429672 480 429700 3946
rect 430868 480 430896 16546
rect 431972 6914 432000 51954
rect 434720 51944 434772 51950
rect 434720 51886 434772 51892
rect 432052 47728 432104 47734
rect 432052 47670 432104 47676
rect 432064 11762 432092 47670
rect 434732 16574 434760 51886
rect 436756 16574 436784 56510
rect 454684 56500 454736 56506
rect 454684 56442 454736 56448
rect 447784 53576 447836 53582
rect 447784 53518 447836 53524
rect 445760 53372 445812 53378
rect 445760 53314 445812 53320
rect 438860 50992 438912 50998
rect 438860 50934 438912 50940
rect 438872 16574 438900 50934
rect 443644 50924 443696 50930
rect 443644 50866 443696 50872
rect 440240 21412 440292 21418
rect 440240 21354 440292 21360
rect 440252 16574 440280 21354
rect 434732 16546 435588 16574
rect 436756 16546 436876 16574
rect 438872 16546 439176 16574
rect 440252 16546 440372 16574
rect 432052 11756 432104 11762
rect 432052 11698 432104 11704
rect 433248 11756 433300 11762
rect 433248 11698 433300 11704
rect 431972 6886 432092 6914
rect 432064 480 432092 6886
rect 433260 480 433288 11698
rect 434444 8424 434496 8430
rect 434444 8366 434496 8372
rect 434456 480 434484 8366
rect 435560 480 435588 16546
rect 436848 4010 436876 16546
rect 437940 8492 437992 8498
rect 437940 8434 437992 8440
rect 436836 4004 436888 4010
rect 436836 3946 436888 3952
rect 436744 3936 436796 3942
rect 436744 3878 436796 3884
rect 436756 480 436784 3878
rect 437952 480 437980 8434
rect 439148 480 439176 16546
rect 440344 480 440372 16546
rect 441528 8560 441580 8566
rect 441528 8502 441580 8508
rect 441540 480 441568 8502
rect 442632 4004 442684 4010
rect 442632 3946 442684 3952
rect 442644 480 442672 3946
rect 443656 3194 443684 50866
rect 445772 16574 445800 53314
rect 447140 24200 447192 24206
rect 447140 24142 447192 24148
rect 447152 16574 447180 24142
rect 445772 16546 446260 16574
rect 447152 16546 447456 16574
rect 445024 8628 445076 8634
rect 445024 8570 445076 8576
rect 443828 3868 443880 3874
rect 443828 3810 443880 3816
rect 443644 3188 443696 3194
rect 443644 3130 443696 3136
rect 443840 480 443868 3810
rect 445036 480 445064 8570
rect 446232 480 446260 16546
rect 447428 480 447456 16546
rect 447796 4010 447824 53518
rect 450544 53440 450596 53446
rect 450544 53382 450596 53388
rect 448612 8696 448664 8702
rect 448612 8638 448664 8644
rect 447784 4004 447836 4010
rect 447784 3946 447836 3952
rect 448624 480 448652 8638
rect 450556 3874 450584 53382
rect 452660 51876 452712 51882
rect 452660 51818 452712 51824
rect 452672 16574 452700 51818
rect 454040 22772 454092 22778
rect 454040 22714 454092 22720
rect 454052 16574 454080 22714
rect 452672 16546 453344 16574
rect 454052 16546 454540 16574
rect 452108 8764 452160 8770
rect 452108 8706 452160 8712
rect 450544 3868 450596 3874
rect 450544 3810 450596 3816
rect 450912 3800 450964 3806
rect 450912 3742 450964 3748
rect 449808 3188 449860 3194
rect 449808 3130 449860 3136
rect 449820 480 449848 3130
rect 450924 480 450952 3742
rect 452120 480 452148 8706
rect 453316 480 453344 16546
rect 454512 480 454540 16546
rect 454696 3942 454724 56442
rect 468484 56432 468536 56438
rect 468484 56374 468536 56380
rect 461584 56364 461636 56370
rect 461584 56306 461636 56312
rect 456892 50856 456944 50862
rect 456892 50798 456944 50804
rect 455696 8832 455748 8838
rect 455696 8774 455748 8780
rect 454684 3936 454736 3942
rect 454684 3878 454736 3884
rect 455708 480 455736 8774
rect 456904 480 456932 50798
rect 460940 47660 460992 47666
rect 460940 47602 460992 47608
rect 460388 13932 460440 13938
rect 460388 13874 460440 13880
rect 459192 8900 459244 8906
rect 459192 8842 459244 8848
rect 458088 3732 458140 3738
rect 458088 3674 458140 3680
rect 458100 480 458128 3674
rect 459204 480 459232 8842
rect 460400 480 460428 13874
rect 460952 6914 460980 47602
rect 461596 16574 461624 56306
rect 467840 24132 467892 24138
rect 467840 24074 467892 24080
rect 467852 16574 467880 24074
rect 461596 16546 461716 16574
rect 467852 16546 468432 16574
rect 460952 6886 461624 6914
rect 461596 480 461624 6886
rect 461688 3738 461716 16546
rect 467472 14068 467524 14074
rect 467472 14010 467524 14016
rect 463976 14000 464028 14006
rect 463976 13942 464028 13948
rect 462780 9648 462832 9654
rect 462780 9590 462832 9596
rect 461676 3732 461728 3738
rect 461676 3674 461728 3680
rect 462792 480 462820 9590
rect 463988 480 464016 13942
rect 466276 9580 466328 9586
rect 466276 9522 466328 9528
rect 465172 3664 465224 3670
rect 465172 3606 465224 3612
rect 465184 480 465212 3606
rect 466288 480 466316 9522
rect 467484 480 467512 14010
rect 468404 3074 468432 16546
rect 468496 3262 468524 56374
rect 472624 56296 472676 56302
rect 472624 56238 472676 56244
rect 471060 14136 471112 14142
rect 471060 14078 471112 14084
rect 469864 9512 469916 9518
rect 469864 9454 469916 9460
rect 468484 3256 468536 3262
rect 468484 3198 468536 3204
rect 468404 3046 468708 3074
rect 468680 480 468708 3046
rect 469876 480 469904 9454
rect 471072 480 471100 14078
rect 472636 3670 472664 56238
rect 475384 56228 475436 56234
rect 475384 56170 475436 56176
rect 473360 14204 473412 14210
rect 473360 14146 473412 14152
rect 472624 3664 472676 3670
rect 472624 3606 472676 3612
rect 473372 3602 473400 14146
rect 473452 9444 473504 9450
rect 473452 9386 473504 9392
rect 472256 3596 472308 3602
rect 472256 3538 472308 3544
rect 473360 3596 473412 3602
rect 473360 3538 473412 3544
rect 472268 480 472296 3538
rect 473464 480 473492 9386
rect 474556 3596 474608 3602
rect 474556 3538 474608 3544
rect 474568 480 474596 3538
rect 475396 3330 475424 56170
rect 479524 56160 479576 56166
rect 479524 56102 479576 56108
rect 478144 14272 478196 14278
rect 478144 14214 478196 14220
rect 476948 9376 477000 9382
rect 476948 9318 477000 9324
rect 475752 3392 475804 3398
rect 475752 3334 475804 3340
rect 475384 3324 475436 3330
rect 475384 3266 475436 3272
rect 475764 480 475792 3334
rect 476960 480 476988 9318
rect 478156 480 478184 14214
rect 479340 4140 479392 4146
rect 479340 4082 479392 4088
rect 479352 480 479380 4082
rect 479536 4010 479564 56102
rect 483020 56092 483072 56098
rect 483020 56034 483072 56040
rect 483032 16574 483060 56034
rect 500960 56024 501012 56030
rect 500960 55966 501012 55972
rect 485044 54664 485096 54670
rect 485044 54606 485096 54612
rect 483032 16546 484072 16574
rect 481640 14340 481692 14346
rect 481640 14282 481692 14288
rect 479524 4004 479576 4010
rect 479524 3946 479576 3952
rect 480536 3936 480588 3942
rect 480536 3878 480588 3884
rect 480548 480 480576 3878
rect 481652 3602 481680 14282
rect 481732 9308 481784 9314
rect 481732 9250 481784 9256
rect 481640 3596 481692 3602
rect 481640 3538 481692 3544
rect 481744 480 481772 9250
rect 482836 3596 482888 3602
rect 482836 3538 482888 3544
rect 482848 480 482876 3538
rect 484044 480 484072 16546
rect 485056 3670 485084 54606
rect 489184 50788 489236 50794
rect 489184 50730 489236 50736
rect 486424 14408 486476 14414
rect 486424 14350 486476 14356
rect 485228 9240 485280 9246
rect 485228 9182 485280 9188
rect 485044 3664 485096 3670
rect 485044 3606 485096 3612
rect 485240 480 485268 9182
rect 486436 480 486464 14350
rect 488816 9172 488868 9178
rect 488816 9114 488868 9120
rect 487620 3732 487672 3738
rect 487620 3674 487672 3680
rect 487632 480 487660 3674
rect 488828 480 488856 9114
rect 489196 3602 489224 50730
rect 500972 16574 501000 55966
rect 580264 55956 580316 55962
rect 580264 55898 580316 55904
rect 512644 55888 512696 55894
rect 512644 55830 512696 55836
rect 507860 54596 507912 54602
rect 507860 54538 507912 54544
rect 502340 53304 502392 53310
rect 502340 53246 502392 53252
rect 502352 16574 502380 53246
rect 507872 16574 507900 54538
rect 500972 16546 501828 16574
rect 502352 16546 503024 16574
rect 507872 16546 508912 16574
rect 489920 15156 489972 15162
rect 489920 15098 489972 15104
rect 489184 3596 489236 3602
rect 489184 3538 489236 3544
rect 489932 480 489960 15098
rect 493508 15088 493560 15094
rect 493508 15030 493560 15036
rect 492312 9104 492364 9110
rect 492312 9046 492364 9052
rect 491116 3256 491168 3262
rect 491116 3198 491168 3204
rect 491128 480 491156 3198
rect 492324 480 492352 9046
rect 493520 480 493548 15030
rect 497096 15020 497148 15026
rect 497096 14962 497148 14968
rect 495900 9036 495952 9042
rect 495900 8978 495952 8984
rect 494704 3324 494756 3330
rect 494704 3266 494756 3272
rect 494716 480 494744 3266
rect 495912 480 495940 8978
rect 497108 480 497136 14962
rect 500592 14952 500644 14958
rect 500592 14894 500644 14900
rect 499396 8968 499448 8974
rect 499396 8910 499448 8916
rect 498200 3392 498252 3398
rect 498200 3334 498252 3340
rect 498212 480 498240 3334
rect 499408 480 499436 8910
rect 500604 480 500632 14894
rect 501800 480 501828 16546
rect 502996 480 503024 16546
rect 504180 14884 504232 14890
rect 504180 14826 504232 14832
rect 504192 480 504220 14826
rect 507676 14816 507728 14822
rect 507676 14758 507728 14764
rect 505376 4004 505428 4010
rect 505376 3946 505428 3952
rect 505388 480 505416 3946
rect 506480 3800 506532 3806
rect 506480 3742 506532 3748
rect 506492 480 506520 3742
rect 507688 480 507716 14758
rect 508884 480 508912 16546
rect 511264 14748 511316 14754
rect 511264 14690 511316 14696
rect 510068 3868 510120 3874
rect 510068 3810 510120 3816
rect 510080 480 510108 3810
rect 511276 480 511304 14690
rect 512460 4276 512512 4282
rect 512460 4218 512512 4224
rect 512472 480 512500 4218
rect 512656 3398 512684 55830
rect 530584 54528 530636 54534
rect 530584 54470 530636 54476
rect 519544 53236 519596 53242
rect 519544 53178 519596 53184
rect 519556 16574 519584 53178
rect 520280 53168 520332 53174
rect 520280 53110 520332 53116
rect 520292 16574 520320 53110
rect 526444 53100 526496 53106
rect 526444 53042 526496 53048
rect 519556 16546 519676 16574
rect 520292 16546 520780 16574
rect 514760 14680 514812 14686
rect 514760 14622 514812 14628
rect 512644 3392 512696 3398
rect 512644 3334 512696 3340
rect 513564 3392 513616 3398
rect 513564 3334 513616 3340
rect 513576 480 513604 3334
rect 514772 480 514800 14622
rect 518348 14612 518400 14618
rect 518348 14554 518400 14560
rect 515956 4344 516008 4350
rect 515956 4286 516008 4292
rect 515968 480 515996 4286
rect 517152 3664 517204 3670
rect 517152 3606 517204 3612
rect 517164 480 517192 3606
rect 518360 480 518388 14554
rect 519544 4412 519596 4418
rect 519544 4354 519596 4360
rect 519556 480 519584 4354
rect 519648 3262 519676 16546
rect 519636 3256 519688 3262
rect 519636 3198 519688 3204
rect 520752 480 520780 16546
rect 521844 14544 521896 14550
rect 521844 14486 521896 14492
rect 521856 480 521884 14486
rect 525432 14476 525484 14482
rect 525432 14418 525484 14424
rect 523040 4480 523092 4486
rect 523040 4422 523092 4428
rect 523052 480 523080 4422
rect 524236 3256 524288 3262
rect 524236 3198 524288 3204
rect 524248 480 524276 3198
rect 525444 480 525472 14418
rect 526456 3398 526484 53042
rect 528560 51808 528612 51814
rect 528560 51750 528612 51756
rect 528572 16574 528600 51750
rect 528572 16546 529060 16574
rect 526628 4548 526680 4554
rect 526628 4490 526680 4496
rect 526444 3392 526496 3398
rect 526444 3334 526496 3340
rect 526640 480 526668 4490
rect 527824 3392 527876 3398
rect 527824 3334 527876 3340
rect 527836 480 527864 3334
rect 529032 480 529060 16546
rect 530124 4616 530176 4622
rect 530124 4558 530176 4564
rect 530136 480 530164 4558
rect 530596 3602 530624 54470
rect 544384 51740 544436 51746
rect 544384 51682 544436 51688
rect 533344 50720 533396 50726
rect 533344 50662 533396 50668
rect 532516 3664 532568 3670
rect 532516 3606 532568 3612
rect 530584 3596 530636 3602
rect 530584 3538 530636 3544
rect 531320 3596 531372 3602
rect 531320 3538 531372 3544
rect 531332 480 531360 3538
rect 532528 480 532556 3606
rect 533356 3602 533384 50662
rect 537484 50652 537536 50658
rect 537484 50594 537536 50600
rect 535460 50584 535512 50590
rect 535460 50526 535512 50532
rect 535472 16574 535500 50526
rect 535472 16546 536144 16574
rect 534908 10192 534960 10198
rect 534908 10134 534960 10140
rect 533712 4684 533764 4690
rect 533712 4626 533764 4632
rect 533344 3596 533396 3602
rect 533344 3538 533396 3544
rect 533724 480 533752 4626
rect 534920 480 534948 10134
rect 536116 480 536144 16546
rect 537208 4752 537260 4758
rect 537208 4694 537260 4700
rect 537220 480 537248 4694
rect 537496 3670 537524 50594
rect 539600 50516 539652 50522
rect 539600 50458 539652 50464
rect 538404 10260 538456 10266
rect 538404 10202 538456 10208
rect 537484 3664 537536 3670
rect 537484 3606 537536 3612
rect 538416 480 538444 10202
rect 539612 480 539640 50458
rect 542360 50448 542412 50454
rect 542360 50390 542412 50396
rect 542372 16574 542400 50390
rect 542372 16546 543228 16574
rect 541992 11008 542044 11014
rect 541992 10950 542044 10956
rect 540796 5500 540848 5506
rect 540796 5442 540848 5448
rect 540808 480 540836 5442
rect 542004 480 542032 10950
rect 543200 480 543228 16546
rect 544292 5432 544344 5438
rect 544292 5374 544344 5380
rect 544304 1034 544332 5374
rect 544396 3738 544424 51682
rect 546500 50380 546552 50386
rect 546500 50322 546552 50328
rect 546512 16574 546540 50322
rect 580172 46912 580224 46918
rect 580172 46854 580224 46860
rect 580184 46345 580212 46854
rect 580170 46336 580226 46345
rect 580170 46271 580226 46280
rect 580170 33144 580226 33153
rect 580170 33079 580172 33088
rect 580224 33079 580226 33088
rect 580172 33050 580224 33056
rect 580172 20664 580224 20670
rect 580172 20606 580224 20612
rect 580184 19825 580212 20606
rect 580170 19816 580226 19825
rect 580170 19751 580226 19760
rect 546512 16546 546724 16574
rect 545488 10940 545540 10946
rect 545488 10882 545540 10888
rect 544384 3732 544436 3738
rect 544384 3674 544436 3680
rect 544304 1006 544424 1034
rect 544396 480 544424 1006
rect 545500 480 545528 10882
rect 546696 480 546724 16546
rect 560852 16244 560904 16250
rect 560852 16186 560904 16192
rect 547880 10872 547932 10878
rect 547880 10814 547932 10820
rect 547892 3398 547920 10814
rect 552664 10804 552716 10810
rect 552664 10746 552716 10752
rect 547972 5364 548024 5370
rect 547972 5306 548024 5312
rect 547880 3392 547932 3398
rect 547880 3334 547932 3340
rect 547984 2666 548012 5306
rect 551468 5296 551520 5302
rect 551468 5238 551520 5244
rect 550272 3596 550324 3602
rect 550272 3538 550324 3544
rect 549076 3392 549128 3398
rect 549076 3334 549128 3340
rect 547892 2638 548012 2666
rect 547892 480 547920 2638
rect 549088 480 549116 3334
rect 550284 480 550312 3538
rect 551480 480 551508 5238
rect 552676 480 552704 10746
rect 556160 10736 556212 10742
rect 556160 10678 556212 10684
rect 554964 5228 555016 5234
rect 554964 5170 555016 5176
rect 553768 3664 553820 3670
rect 553768 3606 553820 3612
rect 553780 480 553808 3606
rect 554976 480 555004 5170
rect 556172 480 556200 10678
rect 559748 10668 559800 10674
rect 559748 10610 559800 10616
rect 558552 5160 558604 5166
rect 558552 5102 558604 5108
rect 557356 3732 557408 3738
rect 557356 3674 557408 3680
rect 557368 480 557396 3674
rect 558564 480 558592 5102
rect 559760 480 559788 10610
rect 560864 480 560892 16186
rect 564440 16176 564492 16182
rect 564440 16118 564492 16124
rect 563244 10600 563296 10606
rect 563244 10542 563296 10548
rect 562048 5092 562100 5098
rect 562048 5034 562100 5040
rect 562060 480 562088 5034
rect 563256 480 563284 10542
rect 564452 480 564480 16118
rect 568028 16108 568080 16114
rect 568028 16050 568080 16056
rect 566832 10532 566884 10538
rect 566832 10474 566884 10480
rect 565636 5024 565688 5030
rect 565636 4966 565688 4972
rect 565648 480 565676 4966
rect 566844 480 566872 10474
rect 568040 480 568068 16050
rect 571524 16040 571576 16046
rect 571524 15982 571576 15988
rect 570328 10464 570380 10470
rect 570328 10406 570380 10412
rect 569132 4956 569184 4962
rect 569132 4898 569184 4904
rect 569144 480 569172 4898
rect 570340 480 570368 10406
rect 571536 480 571564 15982
rect 575112 15972 575164 15978
rect 575112 15914 575164 15920
rect 572720 10396 572772 10402
rect 572720 10338 572772 10344
rect 572732 3602 572760 10338
rect 572812 4888 572864 4894
rect 572812 4830 572864 4836
rect 572720 3596 572772 3602
rect 572720 3538 572772 3544
rect 572824 2530 572852 4830
rect 573916 3596 573968 3602
rect 573916 3538 573968 3544
rect 572732 2502 572852 2530
rect 572732 480 572760 2502
rect 573928 480 573956 3538
rect 575124 480 575152 15914
rect 578608 15904 578660 15910
rect 578608 15846 578660 15852
rect 577412 10328 577464 10334
rect 577412 10270 577464 10276
rect 576308 4820 576360 4826
rect 576308 4762 576360 4768
rect 576320 480 576348 4762
rect 577424 480 577452 10270
rect 578620 480 578648 15846
rect 580276 6633 580304 55898
rect 580262 6624 580318 6633
rect 580262 6559 580318 6568
rect 582196 4072 582248 4078
rect 582196 4014 582248 4020
rect 581000 3528 581052 3534
rect 581000 3470 581052 3476
rect 581012 480 581040 3470
rect 582208 480 582236 4014
rect 583392 3460 583444 3466
rect 583392 3402 583444 3408
rect 583404 480 583432 3402
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3514 671200 3570 671256
rect 3422 658144 3478 658200
rect 3422 632068 3424 632088
rect 3424 632068 3476 632088
rect 3476 632068 3478 632088
rect 3422 632032 3478 632068
rect 3146 619112 3202 619168
rect 3238 606056 3294 606112
rect 3330 579944 3386 580000
rect 3422 566888 3478 566944
rect 3422 553832 3478 553888
rect 3422 527856 3478 527912
rect 3422 514820 3478 514856
rect 3422 514800 3424 514820
rect 3424 514800 3476 514820
rect 3476 514800 3478 514820
rect 2778 501744 2834 501800
rect 3422 475632 3478 475688
rect 3238 462576 3294 462632
rect 3146 449520 3202 449576
rect 3422 423544 3478 423600
rect 3146 410488 3202 410544
rect 3422 397468 3424 397488
rect 3424 397468 3476 397488
rect 3476 397468 3478 397488
rect 3422 397432 3478 397468
rect 3422 371320 3478 371376
rect 3146 358400 3202 358456
rect 3330 345344 3386 345400
rect 3422 319232 3478 319288
rect 3238 306176 3294 306232
rect 3422 293120 3478 293176
rect 3054 267144 3110 267200
rect 3422 254088 3478 254144
rect 52366 504192 52422 504248
rect 50986 504056 51042 504112
rect 3422 241032 3478 241088
rect 33782 234776 33838 234832
rect 15842 232328 15898 232384
rect 14462 230832 14518 230888
rect 11702 229472 11758 229528
rect 7562 229336 7618 229392
rect 3422 226888 3478 226944
rect 3054 201864 3110 201920
rect 2778 188844 2780 188864
rect 2780 188844 2832 188864
rect 2832 188844 2834 188864
rect 2778 188808 2834 188844
rect 3238 162832 3294 162888
rect 3146 110608 3202 110664
rect 3054 58520 3110 58576
rect 4802 226616 4858 226672
rect 3514 214920 3570 214976
rect 3514 149776 3570 149832
rect 3514 136720 3570 136776
rect 17222 232192 17278 232248
rect 3514 97552 3570 97608
rect 22742 230968 22798 231024
rect 21362 229608 21418 229664
rect 18602 228520 18658 228576
rect 3514 84632 3570 84688
rect 3514 71576 3570 71632
rect 3514 45500 3516 45520
rect 3516 45500 3568 45520
rect 3568 45500 3570 45520
rect 3514 45464 3570 45500
rect 3514 32408 3570 32464
rect 3514 19352 3570 19408
rect 3422 6432 3478 6488
rect 25502 227976 25558 228032
rect 29642 226752 29698 226808
rect 40682 228248 40738 228304
rect 36542 228112 36598 228168
rect 50894 503784 50950 503840
rect 53746 503920 53802 503976
rect 55678 226344 55734 226400
rect 55770 226072 55826 226128
rect 55862 192888 55918 192944
rect 55954 176840 56010 176896
rect 56046 139168 56102 139224
rect 56414 225256 56470 225312
rect 56322 222536 56378 222592
rect 57242 435920 57298 435976
rect 57150 432792 57206 432848
rect 57058 409944 57114 410000
rect 56966 407496 57022 407552
rect 57426 433744 57482 433800
rect 57334 429936 57390 429992
rect 57242 242120 57298 242176
rect 56506 203768 56562 203824
rect 56874 179560 56930 179616
rect 57242 160656 57298 160712
rect 57518 217096 57574 217152
rect 57702 436872 57758 436928
rect 57610 211792 57666 211848
rect 57610 198328 57666 198384
rect 57610 195608 57666 195664
rect 57610 190304 57666 190360
rect 57610 184884 57666 184920
rect 57610 184864 57612 184884
rect 57612 184864 57664 184884
rect 57664 184864 57666 184884
rect 57610 182144 57666 182200
rect 57610 171400 57666 171456
rect 57610 168680 57666 168736
rect 57610 166096 57666 166152
rect 57610 163376 57666 163432
rect 57610 157936 57666 157992
rect 57610 152632 57666 152688
rect 57610 149912 57666 149968
rect 57610 144608 57666 144664
rect 57610 141888 57666 141944
rect 57610 136448 57666 136504
rect 57610 133728 57666 133784
rect 57610 131144 57666 131200
rect 57886 431024 57942 431080
rect 57886 408176 57942 408232
rect 57886 225936 57942 225992
rect 57886 219816 57942 219872
rect 58162 174120 58218 174176
rect 57794 122984 57850 123040
rect 57702 120400 57758 120456
rect 57610 117680 57666 117736
rect 57610 114960 57666 115016
rect 59082 428168 59138 428224
rect 59082 397976 59138 398032
rect 58346 228384 58402 228440
rect 58346 225528 58402 225584
rect 58254 112240 58310 112296
rect 57610 109520 57666 109576
rect 57610 106936 57666 106992
rect 57610 104216 57666 104272
rect 57610 101496 57666 101552
rect 57150 96192 57206 96248
rect 57610 90752 57666 90808
rect 57610 88032 57666 88088
rect 57610 85312 57666 85368
rect 57610 80028 57666 80064
rect 57610 80008 57612 80028
rect 57612 80008 57664 80028
rect 57664 80008 57666 80028
rect 57610 77288 57666 77344
rect 57610 74568 57666 74624
rect 57610 69264 57666 69320
rect 56230 66544 56286 66600
rect 58438 209072 58494 209128
rect 58530 206352 58586 206408
rect 58530 98776 58586 98832
rect 58714 201048 58770 201104
rect 58806 187584 58862 187640
rect 58898 155352 58954 155408
rect 58990 147192 59046 147248
rect 59082 128424 59138 128480
rect 59266 93472 59322 93528
rect 59634 214512 59690 214568
rect 59542 125704 59598 125760
rect 59450 82728 59506 82784
rect 91006 505144 91062 505200
rect 89626 503512 89682 503568
rect 96526 503512 96582 503568
rect 98550 503512 98606 503568
rect 101310 503512 101366 503568
rect 103886 503512 103942 503568
rect 104070 503548 104072 503568
rect 104072 503548 104124 503568
rect 104124 503548 104126 503568
rect 104070 503512 104126 503548
rect 113546 503512 113602 503568
rect 129646 504328 129702 504384
rect 117226 503648 117282 503704
rect 128634 503648 128690 503704
rect 123574 503532 123630 503568
rect 123574 503512 123576 503532
rect 123576 503512 123628 503532
rect 123628 503512 123630 503532
rect 123758 503512 123814 503568
rect 129738 503512 129794 503568
rect 108302 491000 108358 491056
rect 89534 490320 89590 490376
rect 91558 490320 91614 490376
rect 143354 503512 143410 503568
rect 144458 503512 144514 503568
rect 148506 503648 148562 503704
rect 146574 503512 146630 503568
rect 149518 503512 149574 503568
rect 111982 488280 112038 488336
rect 176842 503648 176898 503704
rect 156050 503512 156106 503568
rect 158626 503512 158682 503568
rect 160098 503512 160154 503568
rect 164054 503512 164110 503568
rect 165618 503512 165674 503568
rect 133602 491816 133658 491872
rect 153014 491680 153070 491736
rect 196714 486240 196770 486296
rect 118514 485152 118570 485208
rect 143078 484064 143134 484120
rect 180246 484064 180302 484120
rect 111430 483656 111486 483712
rect 85486 398112 85542 398168
rect 92386 398112 92442 398168
rect 95974 398112 96030 398168
rect 99378 398112 99434 398168
rect 78310 397296 78366 397352
rect 80978 397296 81034 397352
rect 81990 397296 82046 397352
rect 83370 397296 83426 397352
rect 85026 397296 85082 397352
rect 87602 397296 87658 397352
rect 88798 397296 88854 397352
rect 90730 397296 90786 397352
rect 91282 397296 91338 397352
rect 77206 396752 77262 396808
rect 77114 396616 77170 396672
rect 60002 232464 60058 232520
rect 61106 226072 61162 226128
rect 70306 233416 70362 233472
rect 67546 233280 67602 233336
rect 64602 232056 64658 232112
rect 63314 230560 63370 230616
rect 66166 229064 66222 229120
rect 69018 229200 69074 229256
rect 68006 227704 68062 227760
rect 74170 234640 74226 234696
rect 72790 230696 72846 230752
rect 75734 231920 75790 231976
rect 74998 227432 75054 227488
rect 78770 396752 78826 396808
rect 76930 236000 76986 236056
rect 75826 227432 75882 227488
rect 86866 396752 86922 396808
rect 65430 226480 65486 226536
rect 62118 226344 62174 226400
rect 71134 226344 71190 226400
rect 84566 227432 84622 227488
rect 88338 396752 88394 396808
rect 91006 396752 91062 396808
rect 85486 227432 85542 227488
rect 94226 397296 94282 397352
rect 93674 396752 93730 396808
rect 93766 396616 93822 396672
rect 97630 397296 97686 397352
rect 96342 396752 96398 396808
rect 100758 397296 100814 397352
rect 102046 397296 102102 397352
rect 104070 397296 104126 397352
rect 106462 397296 106518 397352
rect 109498 397296 109554 397352
rect 111246 397296 111302 397352
rect 112074 397296 112130 397352
rect 99194 396752 99250 396808
rect 99286 396616 99342 396672
rect 101954 396752 102010 396808
rect 103426 396752 103482 396808
rect 104714 396752 104770 396808
rect 105726 396752 105782 396808
rect 106094 396752 106150 396808
rect 107566 396752 107622 396808
rect 108946 396752 109002 396808
rect 111706 396752 111762 396808
rect 95974 230288 96030 230344
rect 96526 230288 96582 230344
rect 99654 230288 99710 230344
rect 100666 230288 100722 230344
rect 102230 228928 102286 228984
rect 103334 228928 103390 228984
rect 105358 230288 105414 230344
rect 106922 233824 106978 233880
rect 106186 230288 106242 230344
rect 108854 396616 108910 396672
rect 108762 231104 108818 231160
rect 108946 231104 109002 231160
rect 107934 228928 107990 228984
rect 108854 228928 108910 228984
rect 113638 398112 113694 398168
rect 113178 397296 113234 397352
rect 113730 397296 113786 397352
rect 115846 397296 115902 397352
rect 117134 397296 117190 397352
rect 118330 397296 118386 397352
rect 118606 397296 118662 397352
rect 117042 396752 117098 396808
rect 119894 396752 119950 396808
rect 120078 396752 120134 396808
rect 121274 237904 121330 237960
rect 146022 398112 146078 398168
rect 123482 397296 123538 397352
rect 125966 397296 126022 397352
rect 136270 397296 136326 397352
rect 138386 397296 138442 397352
rect 129738 396752 129794 396808
rect 133786 396752 133842 396808
rect 129646 396072 129702 396128
rect 123206 228384 123262 228440
rect 125046 232464 125102 232520
rect 126978 230288 127034 230344
rect 127530 230288 127586 230344
rect 129738 233960 129794 234016
rect 130382 233960 130438 234016
rect 140778 396752 140834 396808
rect 132498 233960 132554 234016
rect 133142 233960 133198 234016
rect 135902 237904 135958 237960
rect 138018 227432 138074 227488
rect 138938 227432 138994 227488
rect 144826 396752 144882 396808
rect 156418 397296 156474 397352
rect 163870 397296 163926 397352
rect 147678 396752 147734 396808
rect 151726 396752 151782 396808
rect 154486 396752 154542 396808
rect 144918 227432 144974 227488
rect 145746 227432 145802 227488
rect 158626 396752 158682 396808
rect 161386 396752 161442 396808
rect 152278 233824 152334 233880
rect 165618 396752 165674 396808
rect 167366 234776 167422 234832
rect 157982 232328 158038 232384
rect 157430 229472 157486 229528
rect 154578 229336 154634 229392
rect 156602 227840 156658 227896
rect 156602 226888 156658 226944
rect 156418 226752 156474 226808
rect 155130 226616 155186 226672
rect 160742 232192 160798 232248
rect 160282 230832 160338 230888
rect 159270 228520 159326 228576
rect 165986 230968 166042 231024
rect 163134 229608 163190 229664
rect 162122 227976 162178 228032
rect 164054 228248 164110 228304
rect 164974 228112 165030 228168
rect 166906 227840 166962 227896
rect 170678 228248 170734 228304
rect 172886 226616 172942 226672
rect 174542 228384 174598 228440
rect 173806 226616 173862 226672
rect 175830 227432 175886 227488
rect 176566 227432 176622 227488
rect 179234 228520 179290 228576
rect 182178 396752 182234 396808
rect 183466 396752 183522 396808
rect 180890 226616 180946 226672
rect 183098 227840 183154 227896
rect 181810 226616 181866 226672
rect 184938 228656 184994 228712
rect 184202 227840 184258 227896
rect 191654 227840 191710 227896
rect 197358 228520 197414 228576
rect 196714 228384 196770 228440
rect 197542 413616 197598 413672
rect 197450 227840 197506 227896
rect 198738 479168 198794 479224
rect 198830 419328 198886 419384
rect 198922 417696 198978 417752
rect 199474 416336 199530 416392
rect 199382 414840 199438 414896
rect 200762 228656 200818 228712
rect 203430 230288 203486 230344
rect 204166 230288 204222 230344
rect 206466 228248 206522 228304
rect 212538 230288 212594 230344
rect 213090 230288 213146 230344
rect 215298 232872 215354 232928
rect 215574 235184 215630 235240
rect 215666 233008 215722 233064
rect 215850 232736 215906 232792
rect 215758 232600 215814 232656
rect 215482 232464 215538 232520
rect 215758 227432 215814 227488
rect 216126 230016 216182 230072
rect 216310 229744 216366 229800
rect 216494 229880 216550 229936
rect 216402 228792 216458 228848
rect 216218 228656 216274 228712
rect 217690 435920 217746 435976
rect 217598 433744 217654 433800
rect 217414 432792 217470 432848
rect 216678 431024 216734 431080
rect 216678 429936 216734 429992
rect 217230 409944 217286 410000
rect 216678 408176 216734 408232
rect 216770 408040 216826 408096
rect 217966 436872 218022 436928
rect 217874 428168 217930 428224
rect 217322 230832 217378 230888
rect 216586 227432 216642 227488
rect 216034 226888 216090 226944
rect 217966 228248 218022 228304
rect 218794 230152 218850 230208
rect 218978 233144 219034 233200
rect 218886 227432 218942 227488
rect 218702 227296 218758 227352
rect 252558 504056 252614 504112
rect 245842 503512 245898 503568
rect 260838 503512 260894 503568
rect 277398 503648 277454 503704
rect 265714 503512 265770 503568
rect 267738 503512 267794 503568
rect 270498 503512 270554 503568
rect 273258 503512 273314 503568
rect 277306 503512 277362 503568
rect 280158 503512 280214 503568
rect 288438 503648 288494 503704
rect 285678 503532 285734 503568
rect 285678 503512 285680 503532
rect 285680 503512 285732 503532
rect 285732 503512 285734 503532
rect 286874 503512 286930 503568
rect 292578 503512 292634 503568
rect 295338 503512 295394 503568
rect 219806 485968 219862 486024
rect 322938 503512 322994 503568
rect 298098 492632 298154 492688
rect 300858 492632 300914 492688
rect 302238 492632 302294 492688
rect 304998 492632 305054 492688
rect 307758 492632 307814 492688
rect 310518 492632 310574 492688
rect 313278 492632 313334 492688
rect 316038 492632 316094 492688
rect 317418 492632 317474 492688
rect 320178 492632 320234 492688
rect 339406 492632 339462 492688
rect 339498 492632 339554 492688
rect 326618 488280 326674 488336
rect 253294 487600 253350 487656
rect 263690 487600 263746 487656
rect 284390 487600 284446 487656
rect 356794 485424 356850 485480
rect 219806 480936 219862 480992
rect 219254 227160 219310 227216
rect 219070 227024 219126 227080
rect 219898 230424 219954 230480
rect 357438 479168 357494 479224
rect 220082 230832 220138 230888
rect 220174 228792 220230 228848
rect 219990 226752 220046 226808
rect 222014 228656 222070 228712
rect 222842 227840 222898 227896
rect 224222 226616 224278 226672
rect 61750 225936 61806 225992
rect 78862 225936 78918 225992
rect 223670 225936 223726 225992
rect 59726 71984 59782 72040
rect 59174 61240 59230 61296
rect 221738 60152 221794 60208
rect 58714 57840 58770 57896
rect 207294 57296 207350 57352
rect 208766 57160 208822 57216
rect 208490 56888 208546 56944
rect 210238 59200 210294 59256
rect 212354 59336 212410 59392
rect 211158 57432 211214 57488
rect 214746 57840 214802 57896
rect 213826 57024 213882 57080
rect 216494 57704 216550 57760
rect 218242 57840 218298 57896
rect 219530 57840 219586 57896
rect 219714 57840 219770 57896
rect 222934 60016 222990 60072
rect 223302 59880 223358 59936
rect 219530 57568 219586 57624
rect 224590 232872 224646 232928
rect 224682 230016 224738 230072
rect 224590 60152 224646 60208
rect 224866 226616 224922 226672
rect 224774 224984 224830 225040
rect 224958 59336 225014 59392
rect 225326 232736 225382 232792
rect 225510 230424 225566 230480
rect 225418 222536 225474 222592
rect 225602 229880 225658 229936
rect 225510 60016 225566 60072
rect 225694 229744 225750 229800
rect 225602 57840 225658 57896
rect 225878 227296 225934 227352
rect 225786 226752 225842 226808
rect 225786 59880 225842 59936
rect 226246 230152 226302 230208
rect 226154 195608 226210 195664
rect 226062 141888 226118 141944
rect 225970 131144 226026 131200
rect 225878 57704 225934 57760
rect 226706 182144 226762 182200
rect 226706 175208 226762 175264
rect 226706 174120 226762 174176
rect 226706 169632 226762 169688
rect 226706 168680 226762 168736
rect 226614 157936 226670 157992
rect 226522 149912 226578 149968
rect 226430 139168 226486 139224
rect 226430 126928 226486 126984
rect 226430 125704 226486 125760
rect 226338 109520 226394 109576
rect 226430 73072 226486 73128
rect 226430 71984 226486 72040
rect 226890 88032 226946 88088
rect 227074 235184 227130 235240
rect 227534 233144 227590 233200
rect 227442 232600 227498 232656
rect 227350 227160 227406 227216
rect 227258 227024 227314 227080
rect 227166 224984 227222 225040
rect 227166 220904 227222 220960
rect 227166 220768 227222 220824
rect 227166 219816 227222 219872
rect 227166 219680 227222 219736
rect 227074 128424 227130 128480
rect 227626 228248 227682 228304
rect 227626 219680 227682 219736
rect 227626 219544 227682 219600
rect 227534 217096 227590 217152
rect 227626 214512 227682 214568
rect 227534 212472 227590 212528
rect 227534 211792 227590 211848
rect 227442 198328 227498 198384
rect 227350 166096 227406 166152
rect 227258 144608 227314 144664
rect 227166 122984 227222 123040
rect 226982 80008 227038 80064
rect 226798 63824 226854 63880
rect 226246 57568 226302 57624
rect 228086 163376 228142 163432
rect 228454 184864 228510 184920
rect 228362 179560 228418 179616
rect 228270 171400 228326 171456
rect 228178 160656 228234 160712
rect 228086 91704 228142 91760
rect 228086 90752 228142 90808
rect 228638 209072 228694 209128
rect 225326 57024 225382 57080
rect 228914 206352 228970 206408
rect 229006 176840 229062 176896
rect 228822 74568 228878 74624
rect 229558 226888 229614 226944
rect 229650 104216 229706 104272
rect 229926 233416 229982 233472
rect 229926 151816 229982 151872
rect 229834 117680 229890 117736
rect 229742 98776 229798 98832
rect 230754 190304 230810 190360
rect 230662 152632 230718 152688
rect 231214 234640 231270 234696
rect 231214 178064 231270 178120
rect 231122 112240 231178 112296
rect 232042 96192 232098 96248
rect 232594 232056 232650 232112
rect 232502 126928 232558 126984
rect 232318 120400 232374 120456
rect 232226 101496 232282 101552
rect 232134 93472 232190 93528
rect 232686 212472 232742 212528
rect 232594 71848 232650 71904
rect 231950 61240 232006 61296
rect 235998 398112 236054 398168
rect 265070 398112 265126 398168
rect 300122 398112 300178 398168
rect 315762 398112 315818 398168
rect 325882 398112 325938 398168
rect 237010 397296 237066 397352
rect 238114 397296 238170 397352
rect 239218 397296 239274 397352
rect 240506 397296 240562 397352
rect 241610 397296 241666 397352
rect 247682 397296 247738 397352
rect 249982 397296 250038 397352
rect 251178 397296 251234 397352
rect 252742 397296 252798 397352
rect 259826 397296 259882 397352
rect 262034 397296 262090 397352
rect 233514 77288 233570 77344
rect 233882 193840 233938 193896
rect 233882 192888 233938 192944
rect 235354 203768 235410 203824
rect 235262 73072 235318 73128
rect 233698 66544 233754 66600
rect 238114 133728 238170 133784
rect 242898 396772 242954 396808
rect 242898 396752 242900 396772
rect 242900 396752 242952 396772
rect 242952 396752 242954 396772
rect 244370 396752 244426 396808
rect 245658 396752 245714 396808
rect 247590 396752 247646 396808
rect 248418 396752 248474 396808
rect 244278 396616 244334 396672
rect 240874 155896 240930 155952
rect 244922 147600 244978 147656
rect 244278 82728 244334 82784
rect 246302 169632 246358 169688
rect 249798 396752 249854 396808
rect 251270 397160 251326 397216
rect 252650 396752 252706 396808
rect 258078 396888 258134 396944
rect 254490 396752 254546 396808
rect 255410 396752 255466 396808
rect 256882 396772 256938 396808
rect 256882 396752 256884 396772
rect 256884 396752 256936 396772
rect 256936 396752 256938 396772
rect 255318 396616 255374 396672
rect 253202 136584 253258 136640
rect 255318 91704 255374 91760
rect 258170 396752 258226 396808
rect 259550 396752 259606 396808
rect 260930 396752 260986 396808
rect 262218 396752 262274 396808
rect 263598 396752 263654 396808
rect 262218 175208 262274 175264
rect 263690 396616 263746 396672
rect 265898 397296 265954 397352
rect 268290 397296 268346 397352
rect 270866 397296 270922 397352
rect 272246 397296 272302 397352
rect 273442 397296 273498 397352
rect 276202 397296 276258 397352
rect 276386 397296 276442 397352
rect 278042 397316 278098 397352
rect 278042 397296 278044 397316
rect 278044 397296 278096 397316
rect 278096 397296 278098 397316
rect 266358 396752 266414 396808
rect 267830 396752 267886 396808
rect 266450 396616 266506 396672
rect 269118 396752 269174 396808
rect 270590 396752 270646 396808
rect 267830 193840 267886 193896
rect 273350 397160 273406 397216
rect 273258 396772 273314 396808
rect 273258 396752 273260 396772
rect 273260 396752 273312 396772
rect 273312 396752 273314 396772
rect 274638 396752 274694 396808
rect 278962 397296 279018 397352
rect 283194 397296 283250 397352
rect 289818 397296 289874 397352
rect 298466 397296 298522 397352
rect 277490 396752 277546 396808
rect 280158 396752 280214 396808
rect 278042 230696 278098 230752
rect 271142 229200 271198 229256
rect 285678 396752 285734 396808
rect 287058 396752 287114 396808
rect 287702 230560 287758 230616
rect 282182 220768 282238 220824
rect 292946 396752 293002 396808
rect 295890 396772 295946 396808
rect 295890 396752 295892 396772
rect 295892 396752 295944 396772
rect 295944 396752 295946 396772
rect 295982 226480 296038 226536
rect 302238 396752 302294 396808
rect 305274 396752 305330 396808
rect 307850 396772 307906 396808
rect 307850 396752 307852 396772
rect 307852 396752 307904 396772
rect 307904 396752 307906 396772
rect 310518 396752 310574 396808
rect 313278 396752 313334 396808
rect 302882 227704 302938 227760
rect 300122 187584 300178 187640
rect 307022 201320 307078 201376
rect 317418 396752 317474 396808
rect 320178 396752 320234 396808
rect 323122 396752 323178 396808
rect 343362 397296 343418 397352
rect 342350 396752 342406 396808
rect 357622 415792 357678 415848
rect 357530 413072 357586 413128
rect 358818 418784 358874 418840
rect 357438 60288 357494 60344
rect 358910 417152 358966 417208
rect 358818 59200 358874 59256
rect 359002 414296 359058 414352
rect 580170 697176 580226 697232
rect 580170 683848 580226 683904
rect 580170 670692 580172 670712
rect 580172 670692 580224 670712
rect 580224 670692 580226 670712
rect 580170 670656 580226 670692
rect 580170 644000 580226 644056
rect 580170 630808 580226 630864
rect 580170 617480 580226 617536
rect 579802 590960 579858 591016
rect 580170 577632 580226 577688
rect 579802 564304 579858 564360
rect 580170 537784 580226 537840
rect 580170 524476 580226 524512
rect 580170 524456 580172 524476
rect 580172 524456 580224 524476
rect 580224 524456 580226 524476
rect 580170 511264 580226 511320
rect 580170 484608 580226 484664
rect 579986 471416 580042 471472
rect 580170 458088 580226 458144
rect 580170 431568 580226 431624
rect 580262 418240 580318 418296
rect 580170 404912 580226 404968
rect 580170 378392 580226 378448
rect 579618 365064 579674 365120
rect 580170 351908 580172 351928
rect 580172 351908 580224 351928
rect 580224 351908 580226 351928
rect 580170 351872 580226 351908
rect 580170 325216 580226 325272
rect 579986 312024 580042 312080
rect 580170 298696 580226 298752
rect 580170 272176 580226 272232
rect 580170 258848 580226 258904
rect 579802 245520 579858 245576
rect 580262 229064 580318 229120
rect 410522 226344 410578 226400
rect 580170 205672 580226 205728
rect 580170 192480 580226 192536
rect 580170 165824 580226 165880
rect 580170 139340 580172 139360
rect 580172 139340 580224 139360
rect 580224 139340 580226 139360
rect 580170 139304 580226 139340
rect 580170 125976 580226 126032
rect 580170 99456 580226 99512
rect 580262 86128 580318 86184
rect 580170 59608 580226 59664
rect 356518 57160 356574 57216
rect 580170 46280 580226 46336
rect 580170 33108 580226 33144
rect 580170 33088 580172 33108
rect 580172 33088 580224 33108
rect 580224 33088 580226 33108
rect 580170 19760 580226 19816
rect 580262 6568 580318 6624
<< metal3 >>
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3417 658202 3483 658205
rect -960 658200 3483 658202
rect -960 658144 3422 658200
rect 3478 658144 3483 658200
rect -960 658142 3483 658144
rect -960 658052 480 658142
rect 3417 658139 3483 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3417 632090 3483 632093
rect -960 632088 3483 632090
rect -960 632032 3422 632088
rect 3478 632032 3483 632088
rect -960 632030 3483 632032
rect -960 631940 480 632030
rect 3417 632027 3483 632030
rect 580165 630866 580231 630869
rect 583520 630866 584960 630956
rect 580165 630864 584960 630866
rect 580165 630808 580170 630864
rect 580226 630808 584960 630864
rect 580165 630806 584960 630808
rect 580165 630803 580231 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3141 619170 3207 619173
rect -960 619168 3207 619170
rect -960 619112 3146 619168
rect 3202 619112 3207 619168
rect -960 619110 3207 619112
rect -960 619020 480 619110
rect 3141 619107 3207 619110
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3233 606114 3299 606117
rect -960 606112 3299 606114
rect -960 606056 3238 606112
rect 3294 606056 3299 606112
rect -960 606054 3299 606056
rect -960 605964 480 606054
rect 3233 606051 3299 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 579797 591018 579863 591021
rect 583520 591018 584960 591108
rect 579797 591016 584960 591018
rect 579797 590960 579802 591016
rect 579858 590960 584960 591016
rect 579797 590958 584960 590960
rect 579797 590955 579863 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 3325 580002 3391 580005
rect -960 580000 3391 580002
rect -960 579944 3330 580000
rect 3386 579944 3391 580000
rect -960 579942 3391 579944
rect -960 579852 480 579942
rect 3325 579939 3391 579942
rect 580165 577690 580231 577693
rect 583520 577690 584960 577780
rect 580165 577688 584960 577690
rect 580165 577632 580170 577688
rect 580226 577632 584960 577688
rect 580165 577630 584960 577632
rect 580165 577627 580231 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3417 566946 3483 566949
rect -960 566944 3483 566946
rect -960 566888 3422 566944
rect 3478 566888 3483 566944
rect -960 566886 3483 566888
rect -960 566796 480 566886
rect 3417 566883 3483 566886
rect 579797 564362 579863 564365
rect 583520 564362 584960 564452
rect 579797 564360 584960 564362
rect 579797 564304 579802 564360
rect 579858 564304 584960 564360
rect 579797 564302 584960 564304
rect 579797 564299 579863 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 3417 553890 3483 553893
rect -960 553888 3483 553890
rect -960 553832 3422 553888
rect 3478 553832 3483 553888
rect -960 553830 3483 553832
rect -960 553740 480 553830
rect 3417 553827 3483 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 580165 537842 580231 537845
rect 583520 537842 584960 537932
rect 580165 537840 584960 537842
rect 580165 537784 580170 537840
rect 580226 537784 584960 537840
rect 580165 537782 584960 537784
rect 580165 537779 580231 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 3417 527914 3483 527917
rect -960 527912 3483 527914
rect -960 527856 3422 527912
rect 3478 527856 3483 527912
rect -960 527854 3483 527856
rect -960 527764 480 527854
rect 3417 527851 3483 527854
rect 580165 524514 580231 524517
rect 583520 524514 584960 524604
rect 580165 524512 584960 524514
rect 580165 524456 580170 524512
rect 580226 524456 584960 524512
rect 580165 524454 584960 524456
rect 580165 524451 580231 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 3417 514858 3483 514861
rect -960 514856 3483 514858
rect -960 514800 3422 514856
rect 3478 514800 3483 514856
rect -960 514798 3483 514800
rect -960 514708 480 514798
rect 3417 514795 3483 514798
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect 91001 505202 91067 505205
rect 218646 505202 218652 505204
rect 91001 505200 218652 505202
rect 91001 505144 91006 505200
rect 91062 505144 218652 505200
rect 91001 505142 218652 505144
rect 91001 505139 91067 505142
rect 218646 505140 218652 505142
rect 218716 505140 218722 505204
rect 128670 504324 128676 504388
rect 128740 504386 128746 504388
rect 129641 504386 129707 504389
rect 128740 504384 129707 504386
rect 128740 504328 129646 504384
rect 129702 504328 129707 504384
rect 128740 504326 129707 504328
rect 128740 504324 128746 504326
rect 129641 504323 129707 504326
rect 52361 504250 52427 504253
rect 248454 504250 248460 504252
rect 52361 504248 248460 504250
rect 52361 504192 52366 504248
rect 52422 504192 248460 504248
rect 52361 504190 248460 504192
rect 52361 504187 52427 504190
rect 248454 504188 248460 504190
rect 248524 504188 248530 504252
rect 50981 504114 51047 504117
rect 252553 504114 252619 504117
rect 50981 504112 252619 504114
rect 50981 504056 50986 504112
rect 51042 504056 252558 504112
rect 252614 504056 252619 504112
rect 50981 504054 252619 504056
rect 50981 504051 51047 504054
rect 252553 504051 252619 504054
rect 53741 503978 53807 503981
rect 258390 503978 258396 503980
rect 53741 503976 258396 503978
rect 53741 503920 53746 503976
rect 53802 503920 258396 503976
rect 53741 503918 258396 503920
rect 53741 503915 53807 503918
rect 258390 503916 258396 503918
rect 258460 503916 258466 503980
rect 50889 503842 50955 503845
rect 256182 503842 256188 503844
rect 50889 503840 256188 503842
rect 50889 503784 50894 503840
rect 50950 503784 256188 503840
rect 50889 503782 256188 503784
rect 50889 503779 50955 503782
rect 256182 503780 256188 503782
rect 256252 503780 256258 503844
rect 116158 503644 116164 503708
rect 116228 503706 116234 503708
rect 117221 503706 117287 503709
rect 116228 503704 117287 503706
rect 116228 503648 117226 503704
rect 117282 503648 117287 503704
rect 116228 503646 117287 503648
rect 116228 503644 116234 503646
rect 117221 503643 117287 503646
rect 128629 503706 128695 503709
rect 134926 503706 134932 503708
rect 128629 503704 134932 503706
rect 128629 503648 128634 503704
rect 128690 503648 134932 503704
rect 128629 503646 134932 503648
rect 128629 503643 128695 503646
rect 134926 503644 134932 503646
rect 134996 503644 135002 503708
rect 148501 503706 148567 503709
rect 151118 503706 151124 503708
rect 148501 503704 151124 503706
rect 148501 503648 148506 503704
rect 148562 503648 151124 503704
rect 148501 503646 151124 503648
rect 148501 503643 148567 503646
rect 151118 503644 151124 503646
rect 151188 503644 151194 503708
rect 176837 503706 176903 503709
rect 178534 503706 178540 503708
rect 176837 503704 178540 503706
rect 176837 503648 176842 503704
rect 176898 503648 178540 503704
rect 176837 503646 178540 503648
rect 176837 503643 176903 503646
rect 178534 503644 178540 503646
rect 178604 503644 178610 503708
rect 277393 503706 277459 503709
rect 278446 503706 278452 503708
rect 277393 503704 278452 503706
rect 277393 503648 277398 503704
rect 277454 503648 278452 503704
rect 277393 503646 278452 503648
rect 277393 503643 277459 503646
rect 278446 503644 278452 503646
rect 278516 503644 278522 503708
rect 288433 503706 288499 503709
rect 288566 503706 288572 503708
rect 288433 503704 288572 503706
rect 288433 503648 288438 503704
rect 288494 503648 288572 503704
rect 288433 503646 288572 503648
rect 288433 503643 288499 503646
rect 288566 503644 288572 503646
rect 288636 503644 288642 503708
rect 88742 503508 88748 503572
rect 88812 503570 88818 503572
rect 89621 503570 89687 503573
rect 96521 503572 96587 503573
rect 98545 503572 98611 503573
rect 101305 503572 101371 503573
rect 103881 503572 103947 503573
rect 96470 503570 96476 503572
rect 88812 503568 89687 503570
rect 88812 503512 89626 503568
rect 89682 503512 89687 503568
rect 88812 503510 89687 503512
rect 96430 503510 96476 503570
rect 96540 503568 96587 503572
rect 98494 503570 98500 503572
rect 96582 503512 96587 503568
rect 88812 503508 88818 503510
rect 89621 503507 89687 503510
rect 96470 503508 96476 503510
rect 96540 503508 96587 503512
rect 98454 503510 98500 503570
rect 98564 503568 98611 503572
rect 101254 503570 101260 503572
rect 98606 503512 98611 503568
rect 98494 503508 98500 503510
rect 98564 503508 98611 503512
rect 101214 503510 101260 503570
rect 101324 503568 101371 503572
rect 103830 503570 103836 503572
rect 101366 503512 101371 503568
rect 101254 503508 101260 503510
rect 101324 503508 101371 503512
rect 103790 503510 103836 503570
rect 103900 503568 103947 503572
rect 103942 503512 103947 503568
rect 103830 503508 103836 503510
rect 103900 503508 103947 503512
rect 96521 503507 96587 503508
rect 98545 503507 98611 503508
rect 101305 503507 101371 503508
rect 103881 503507 103947 503508
rect 104065 503570 104131 503573
rect 106038 503570 106044 503572
rect 104065 503568 106044 503570
rect 104065 503512 104070 503568
rect 104126 503512 106044 503568
rect 104065 503510 106044 503512
rect 104065 503507 104131 503510
rect 106038 503508 106044 503510
rect 106108 503508 106114 503572
rect 113541 503570 113607 503573
rect 123569 503572 123635 503573
rect 118182 503570 118188 503572
rect 113541 503568 118188 503570
rect 113541 503512 113546 503568
rect 113602 503512 118188 503568
rect 113541 503510 118188 503512
rect 113541 503507 113607 503510
rect 118182 503508 118188 503510
rect 118252 503508 118258 503572
rect 123518 503570 123524 503572
rect 123478 503510 123524 503570
rect 123588 503568 123635 503572
rect 123630 503512 123635 503568
rect 123518 503508 123524 503510
rect 123588 503508 123635 503512
rect 123569 503507 123635 503508
rect 123753 503570 123819 503573
rect 129733 503572 129799 503573
rect 123886 503570 123892 503572
rect 123753 503568 123892 503570
rect 123753 503512 123758 503568
rect 123814 503512 123892 503568
rect 123753 503510 123892 503512
rect 123753 503507 123819 503510
rect 123886 503508 123892 503510
rect 123956 503508 123962 503572
rect 129733 503570 129780 503572
rect 129688 503568 129780 503570
rect 129688 503512 129738 503568
rect 129688 503510 129780 503512
rect 129733 503508 129780 503510
rect 129844 503508 129850 503572
rect 143206 503508 143212 503572
rect 143276 503570 143282 503572
rect 143349 503570 143415 503573
rect 143276 503568 143415 503570
rect 143276 503512 143354 503568
rect 143410 503512 143415 503568
rect 143276 503510 143415 503512
rect 143276 503508 143282 503510
rect 129733 503507 129799 503508
rect 143349 503507 143415 503510
rect 144453 503570 144519 503573
rect 146569 503572 146635 503573
rect 144862 503570 144868 503572
rect 144453 503568 144868 503570
rect 144453 503512 144458 503568
rect 144514 503512 144868 503568
rect 144453 503510 144868 503512
rect 144453 503507 144519 503510
rect 144862 503508 144868 503510
rect 144932 503508 144938 503572
rect 146518 503570 146524 503572
rect 146478 503510 146524 503570
rect 146588 503568 146635 503572
rect 146630 503512 146635 503568
rect 146518 503508 146524 503510
rect 146588 503508 146635 503512
rect 148358 503508 148364 503572
rect 148428 503570 148434 503572
rect 149513 503570 149579 503573
rect 148428 503568 149579 503570
rect 148428 503512 149518 503568
rect 149574 503512 149579 503568
rect 148428 503510 149579 503512
rect 148428 503508 148434 503510
rect 146569 503507 146635 503508
rect 149513 503507 149579 503510
rect 155902 503508 155908 503572
rect 155972 503570 155978 503572
rect 156045 503570 156111 503573
rect 155972 503568 156111 503570
rect 155972 503512 156050 503568
rect 156106 503512 156111 503568
rect 155972 503510 156111 503512
rect 155972 503508 155978 503510
rect 156045 503507 156111 503510
rect 158621 503572 158687 503573
rect 160093 503572 160159 503573
rect 158621 503568 158668 503572
rect 158732 503570 158738 503572
rect 160093 503570 160140 503572
rect 158621 503512 158626 503568
rect 158621 503508 158668 503512
rect 158732 503510 158778 503570
rect 160048 503568 160140 503570
rect 160048 503512 160098 503568
rect 160048 503510 160140 503512
rect 158732 503508 158738 503510
rect 160093 503508 160140 503510
rect 160204 503508 160210 503572
rect 163446 503508 163452 503572
rect 163516 503570 163522 503572
rect 164049 503570 164115 503573
rect 165613 503572 165679 503573
rect 165613 503570 165660 503572
rect 163516 503568 164115 503570
rect 163516 503512 164054 503568
rect 164110 503512 164115 503568
rect 163516 503510 164115 503512
rect 165568 503568 165660 503570
rect 165568 503512 165618 503568
rect 165568 503510 165660 503512
rect 163516 503508 163522 503510
rect 158621 503507 158687 503508
rect 160093 503507 160159 503508
rect 164049 503507 164115 503510
rect 165613 503508 165660 503510
rect 165724 503508 165730 503572
rect 245837 503570 245903 503573
rect 251030 503570 251036 503572
rect 245837 503568 251036 503570
rect 245837 503512 245842 503568
rect 245898 503512 251036 503568
rect 245837 503510 251036 503512
rect 165613 503507 165679 503508
rect 245837 503507 245903 503510
rect 251030 503508 251036 503510
rect 251100 503508 251106 503572
rect 260833 503570 260899 503573
rect 260966 503570 260972 503572
rect 260833 503568 260972 503570
rect 260833 503512 260838 503568
rect 260894 503512 260972 503568
rect 260833 503510 260972 503512
rect 260833 503507 260899 503510
rect 260966 503508 260972 503510
rect 261036 503508 261042 503572
rect 265709 503570 265775 503573
rect 267733 503572 267799 503573
rect 270493 503572 270559 503573
rect 273253 503572 273319 503573
rect 266118 503570 266124 503572
rect 265709 503568 266124 503570
rect 265709 503512 265714 503568
rect 265770 503512 266124 503568
rect 265709 503510 266124 503512
rect 265709 503507 265775 503510
rect 266118 503508 266124 503510
rect 266188 503508 266194 503572
rect 267733 503570 267780 503572
rect 267688 503568 267780 503570
rect 267688 503512 267738 503568
rect 267688 503510 267780 503512
rect 267733 503508 267780 503510
rect 267844 503508 267850 503572
rect 270493 503570 270540 503572
rect 270448 503568 270540 503570
rect 270448 503512 270498 503568
rect 270448 503510 270540 503512
rect 270493 503508 270540 503510
rect 270604 503508 270610 503572
rect 273253 503568 273300 503572
rect 273364 503570 273370 503572
rect 273253 503512 273258 503568
rect 273253 503508 273300 503512
rect 273364 503510 273410 503570
rect 273364 503508 273370 503510
rect 276238 503508 276244 503572
rect 276308 503570 276314 503572
rect 277301 503570 277367 503573
rect 280153 503572 280219 503573
rect 285673 503572 285739 503573
rect 276308 503568 277367 503570
rect 276308 503512 277306 503568
rect 277362 503512 277367 503568
rect 276308 503510 277367 503512
rect 276308 503508 276314 503510
rect 267733 503507 267799 503508
rect 270493 503507 270559 503508
rect 273253 503507 273319 503508
rect 277301 503507 277367 503510
rect 280102 503508 280108 503572
rect 280172 503570 280219 503572
rect 280172 503568 280264 503570
rect 280214 503512 280264 503568
rect 280172 503510 280264 503512
rect 280172 503508 280219 503510
rect 285622 503508 285628 503572
rect 285692 503570 285739 503572
rect 286869 503570 286935 503573
rect 292573 503572 292639 503573
rect 295333 503572 295399 503573
rect 290958 503570 290964 503572
rect 285692 503568 285784 503570
rect 285734 503512 285784 503568
rect 285692 503510 285784 503512
rect 286869 503568 290964 503570
rect 286869 503512 286874 503568
rect 286930 503512 290964 503568
rect 286869 503510 290964 503512
rect 285692 503508 285739 503510
rect 280153 503507 280219 503508
rect 285673 503507 285739 503508
rect 286869 503507 286935 503510
rect 290958 503508 290964 503510
rect 291028 503508 291034 503572
rect 292573 503568 292620 503572
rect 292684 503570 292690 503572
rect 295333 503570 295380 503572
rect 292573 503512 292578 503568
rect 292573 503508 292620 503512
rect 292684 503510 292730 503570
rect 295288 503568 295380 503570
rect 295288 503512 295338 503568
rect 295288 503510 295380 503512
rect 292684 503508 292690 503510
rect 295333 503508 295380 503510
rect 295444 503508 295450 503572
rect 322933 503570 322999 503573
rect 323342 503570 323348 503572
rect 322933 503568 323348 503570
rect 322933 503512 322938 503568
rect 322994 503512 323348 503568
rect 322933 503510 323348 503512
rect 292573 503507 292639 503508
rect 295333 503507 295399 503508
rect 322933 503507 322999 503510
rect 323342 503508 323348 503510
rect 323412 503508 323418 503572
rect -960 501802 480 501892
rect 2773 501802 2839 501805
rect -960 501800 2839 501802
rect -960 501744 2778 501800
rect 2834 501744 2839 501800
rect -960 501742 2839 501744
rect -960 501652 480 501742
rect 2773 501739 2839 501742
rect 583520 497844 584960 498084
rect 298093 492692 298159 492693
rect 300853 492692 300919 492693
rect 302233 492692 302299 492693
rect 304993 492692 305059 492693
rect 307753 492692 307819 492693
rect 310513 492692 310579 492693
rect 313273 492692 313339 492693
rect 316033 492692 316099 492693
rect 298093 492688 298140 492692
rect 298204 492690 298210 492692
rect 298093 492632 298098 492688
rect 298093 492628 298140 492632
rect 298204 492630 298250 492690
rect 300853 492688 300900 492692
rect 300964 492690 300970 492692
rect 300853 492632 300858 492688
rect 298204 492628 298210 492630
rect 300853 492628 300900 492632
rect 300964 492630 301010 492690
rect 300964 492628 300970 492630
rect 302182 492628 302188 492692
rect 302252 492690 302299 492692
rect 302252 492688 302344 492690
rect 302294 492632 302344 492688
rect 302252 492630 302344 492632
rect 302252 492628 302299 492630
rect 304942 492628 304948 492692
rect 305012 492690 305059 492692
rect 305012 492688 305104 492690
rect 305054 492632 305104 492688
rect 305012 492630 305104 492632
rect 305012 492628 305059 492630
rect 307702 492628 307708 492692
rect 307772 492690 307819 492692
rect 307772 492688 307864 492690
rect 307814 492632 307864 492688
rect 307772 492630 307864 492632
rect 307772 492628 307819 492630
rect 310462 492628 310468 492692
rect 310532 492690 310579 492692
rect 310532 492688 310624 492690
rect 310574 492632 310624 492688
rect 310532 492630 310624 492632
rect 310532 492628 310579 492630
rect 313222 492628 313228 492692
rect 313292 492690 313339 492692
rect 313292 492688 313384 492690
rect 313334 492632 313384 492688
rect 313292 492630 313384 492632
rect 313292 492628 313339 492630
rect 316016 492628 316022 492692
rect 316086 492690 316099 492692
rect 317413 492692 317479 492693
rect 320173 492692 320239 492693
rect 339401 492692 339467 492693
rect 316086 492688 316178 492690
rect 316094 492632 316178 492688
rect 316086 492630 316178 492632
rect 317413 492688 317460 492692
rect 317524 492690 317530 492692
rect 317413 492632 317418 492688
rect 316086 492628 316099 492630
rect 298093 492627 298159 492628
rect 300853 492627 300919 492628
rect 302233 492627 302299 492628
rect 304993 492627 305059 492628
rect 307753 492627 307819 492628
rect 310513 492627 310579 492628
rect 313273 492627 313339 492628
rect 316033 492627 316099 492628
rect 317413 492628 317460 492632
rect 317524 492630 317570 492690
rect 320173 492688 320220 492692
rect 320284 492690 320290 492692
rect 320173 492632 320178 492688
rect 317524 492628 317530 492630
rect 320173 492628 320220 492632
rect 320284 492630 320330 492690
rect 320284 492628 320290 492630
rect 339350 492628 339356 492692
rect 339420 492690 339467 492692
rect 339493 492692 339559 492693
rect 339493 492690 339540 492692
rect 339420 492688 339540 492690
rect 339604 492690 339610 492692
rect 339462 492632 339498 492688
rect 339420 492630 339540 492632
rect 339420 492628 339467 492630
rect 317413 492627 317479 492628
rect 320173 492627 320239 492628
rect 339401 492627 339467 492628
rect 339493 492628 339540 492630
rect 339604 492630 339650 492690
rect 339604 492628 339610 492630
rect 339493 492627 339559 492628
rect 133597 491876 133663 491877
rect 133592 491874 133598 491876
rect 133506 491814 133598 491874
rect 133592 491812 133598 491814
rect 133662 491812 133668 491876
rect 133597 491811 133663 491812
rect 153009 491740 153075 491741
rect 153004 491676 153010 491740
rect 153074 491738 153080 491740
rect 153074 491678 153166 491738
rect 153074 491676 153080 491678
rect 153009 491675 153075 491676
rect 108297 491060 108363 491061
rect 108292 490996 108298 491060
rect 108362 491058 108368 491060
rect 108362 490998 108454 491058
rect 108362 490996 108368 490998
rect 108297 490995 108363 490996
rect 89529 490380 89595 490381
rect 91553 490380 91619 490381
rect 89524 490316 89530 490380
rect 89594 490378 89600 490380
rect 89594 490318 89686 490378
rect 89594 490316 89600 490318
rect 91548 490316 91554 490380
rect 91618 490378 91624 490380
rect 91618 490318 91710 490378
rect 91618 490316 91624 490318
rect 89529 490315 89595 490316
rect 91553 490315 91619 490316
rect -960 488596 480 488836
rect 111977 488340 112043 488341
rect 326613 488340 326679 488341
rect 111972 488276 111978 488340
rect 112042 488338 112048 488340
rect 326608 488338 326614 488340
rect 112042 488278 112134 488338
rect 326522 488278 326614 488338
rect 112042 488276 112048 488278
rect 326608 488276 326614 488278
rect 326678 488276 326684 488340
rect 111977 488275 112043 488276
rect 326613 488275 326679 488276
rect 253289 487660 253355 487661
rect 263685 487660 263751 487661
rect 284385 487660 284451 487661
rect 253284 487596 253290 487660
rect 253354 487658 253360 487660
rect 263680 487658 263686 487660
rect 253354 487598 253446 487658
rect 263594 487598 263686 487658
rect 253354 487596 253360 487598
rect 263680 487596 263686 487598
rect 263750 487596 263756 487660
rect 284380 487596 284386 487660
rect 284450 487658 284456 487660
rect 284450 487598 284542 487658
rect 284450 487596 284456 487598
rect 253289 487595 253355 487596
rect 263685 487595 263751 487596
rect 284385 487595 284451 487596
rect 196709 486300 196775 486301
rect 196709 486296 196756 486300
rect 196820 486298 196826 486300
rect 196709 486240 196714 486296
rect 196709 486236 196756 486240
rect 196820 486238 196866 486298
rect 196820 486236 196826 486238
rect 196709 486235 196775 486236
rect 219801 486028 219867 486029
rect 219750 486026 219756 486028
rect 219710 485966 219756 486026
rect 219820 486024 219867 486028
rect 219862 485968 219867 486024
rect 219750 485964 219756 485966
rect 219820 485964 219867 485968
rect 219801 485963 219867 485964
rect 356789 485484 356855 485485
rect 356789 485480 356836 485484
rect 356900 485482 356906 485484
rect 356789 485424 356794 485480
rect 356789 485420 356836 485424
rect 356900 485422 356946 485482
rect 356900 485420 356906 485422
rect 356789 485419 356855 485420
rect 118509 485212 118575 485213
rect 118504 485210 118510 485212
rect 118418 485150 118510 485210
rect 118504 485148 118510 485150
rect 118574 485148 118580 485212
rect 118509 485147 118575 485148
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 583520 484516 584960 484606
rect 143073 484124 143139 484125
rect 180241 484124 180307 484125
rect 143022 484060 143028 484124
rect 143092 484122 143139 484124
rect 143092 484120 143184 484122
rect 143134 484064 143184 484120
rect 143092 484062 143184 484064
rect 143092 484060 143139 484062
rect 180190 484060 180196 484124
rect 180260 484122 180307 484124
rect 180260 484120 180352 484122
rect 180302 484064 180352 484120
rect 180260 484062 180352 484064
rect 180260 484060 180307 484062
rect 143073 484059 143139 484060
rect 180241 484059 180307 484060
rect 111425 483716 111491 483717
rect 111374 483652 111380 483716
rect 111444 483714 111491 483716
rect 111444 483712 111536 483714
rect 111486 483656 111536 483712
rect 111444 483654 111536 483656
rect 111444 483652 111491 483654
rect 111425 483651 111491 483652
rect 219801 480996 219867 480997
rect 219750 480994 219756 480996
rect 219710 480934 219756 480994
rect 219820 480992 219867 480996
rect 219862 480936 219867 480992
rect 219750 480932 219756 480934
rect 219820 480932 219867 480936
rect 219801 480931 219867 480932
rect 198733 479226 198799 479229
rect 357433 479226 357499 479229
rect 197126 479224 198799 479226
rect 197126 479220 198738 479224
rect 196604 479168 198738 479220
rect 198794 479168 198799 479224
rect 357206 479224 357499 479226
rect 357206 479220 357438 479224
rect 196604 479166 198799 479168
rect 196604 479160 197186 479166
rect 198733 479163 198799 479166
rect 356592 479168 357438 479220
rect 357494 479168 357499 479224
rect 356592 479166 357499 479168
rect 356592 479160 357266 479166
rect 357433 479163 357499 479166
rect -960 475690 480 475780
rect 3417 475690 3483 475693
rect -960 475688 3483 475690
rect -960 475632 3422 475688
rect 3478 475632 3483 475688
rect -960 475630 3483 475632
rect -960 475540 480 475630
rect 3417 475627 3483 475630
rect 579981 471474 580047 471477
rect 583520 471474 584960 471564
rect 579981 471472 584960 471474
rect 579981 471416 579986 471472
rect 580042 471416 584960 471472
rect 579981 471414 584960 471416
rect 579981 471411 580047 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 3233 462634 3299 462637
rect -960 462632 3299 462634
rect -960 462576 3238 462632
rect 3294 462576 3299 462632
rect -960 462574 3299 462576
rect -960 462484 480 462574
rect 3233 462571 3299 462574
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 580165 458083 580231 458086
rect 583520 457996 584960 458086
rect -960 449578 480 449668
rect 3141 449578 3207 449581
rect -960 449576 3207 449578
rect -960 449520 3146 449576
rect 3202 449520 3207 449576
rect -960 449518 3207 449520
rect -960 449428 480 449518
rect 3141 449515 3207 449518
rect 583520 444668 584960 444908
rect 57697 436930 57763 436933
rect 217961 436930 218027 436933
rect 57697 436928 59554 436930
rect 57697 436872 57702 436928
rect 57758 436924 59554 436928
rect 217961 436928 219450 436930
rect 57758 436872 60032 436924
rect 57697 436870 60032 436872
rect 57697 436867 57763 436870
rect 59494 436864 60032 436870
rect 217961 436872 217966 436928
rect 218022 436924 219450 436928
rect 218022 436872 220064 436924
rect 217961 436870 220064 436872
rect 217961 436867 218027 436870
rect 219390 436864 220064 436870
rect -960 436508 480 436748
rect 57237 435978 57303 435981
rect 217685 435978 217751 435981
rect 57237 435976 59554 435978
rect 57237 435920 57242 435976
rect 57298 435972 59554 435976
rect 217685 435976 219450 435978
rect 57298 435920 60032 435972
rect 57237 435918 60032 435920
rect 57237 435915 57303 435918
rect 59494 435912 60032 435918
rect 217685 435920 217690 435976
rect 217746 435972 219450 435976
rect 217746 435920 220064 435972
rect 217685 435918 220064 435920
rect 217685 435915 217751 435918
rect 219390 435912 220064 435918
rect 57421 433802 57487 433805
rect 217593 433802 217659 433805
rect 57421 433800 59554 433802
rect 57421 433744 57426 433800
rect 57482 433796 59554 433800
rect 217593 433800 219450 433802
rect 57482 433744 60032 433796
rect 57421 433742 60032 433744
rect 57421 433739 57487 433742
rect 59494 433736 60032 433742
rect 217593 433744 217598 433800
rect 217654 433796 219450 433800
rect 217654 433744 220064 433796
rect 217593 433742 220064 433744
rect 217593 433739 217659 433742
rect 219390 433736 220064 433742
rect 57145 432850 57211 432853
rect 217409 432850 217475 432853
rect 57145 432848 59554 432850
rect 57145 432792 57150 432848
rect 57206 432844 59554 432848
rect 217409 432848 219450 432850
rect 57206 432792 60032 432844
rect 57145 432790 60032 432792
rect 57145 432787 57211 432790
rect 59494 432784 60032 432790
rect 217409 432792 217414 432848
rect 217470 432844 219450 432848
rect 217470 432792 220064 432844
rect 217409 432790 220064 432792
rect 217409 432787 217475 432790
rect 219390 432784 220064 432790
rect 580165 431626 580231 431629
rect 583520 431626 584960 431716
rect 580165 431624 584960 431626
rect 580165 431568 580170 431624
rect 580226 431568 584960 431624
rect 580165 431566 584960 431568
rect 580165 431563 580231 431566
rect 583520 431476 584960 431566
rect 57881 431082 57947 431085
rect 216673 431082 216739 431085
rect 57881 431080 59554 431082
rect 57881 431024 57886 431080
rect 57942 431076 59554 431080
rect 216673 431080 219450 431082
rect 57942 431024 60032 431076
rect 57881 431022 60032 431024
rect 57881 431019 57947 431022
rect 59494 431016 60032 431022
rect 216673 431024 216678 431080
rect 216734 431076 219450 431080
rect 216734 431024 220064 431076
rect 216673 431022 220064 431024
rect 216673 431019 216739 431022
rect 219390 431016 220064 431022
rect 57329 429994 57395 429997
rect 216673 429994 216739 429997
rect 57329 429992 59554 429994
rect 57329 429936 57334 429992
rect 57390 429988 59554 429992
rect 216673 429992 219450 429994
rect 57390 429936 60032 429988
rect 57329 429934 60032 429936
rect 57329 429931 57395 429934
rect 59494 429928 60032 429934
rect 216673 429936 216678 429992
rect 216734 429988 219450 429992
rect 216734 429936 220064 429988
rect 216673 429934 220064 429936
rect 216673 429931 216739 429934
rect 219390 429928 220064 429934
rect 59077 428226 59143 428229
rect 217869 428226 217935 428229
rect 59077 428224 59554 428226
rect 59077 428168 59082 428224
rect 59138 428220 59554 428224
rect 217869 428224 219450 428226
rect 59138 428168 60032 428220
rect 59077 428166 60032 428168
rect 59077 428163 59143 428166
rect 59494 428160 60032 428166
rect 217869 428168 217874 428224
rect 217930 428220 219450 428224
rect 217930 428168 220064 428220
rect 217869 428166 220064 428168
rect 217869 428163 217935 428166
rect 219390 428160 220064 428166
rect -960 423602 480 423692
rect 3417 423602 3483 423605
rect -960 423600 3483 423602
rect -960 423544 3422 423600
rect 3478 423544 3483 423600
rect -960 423542 3483 423544
rect -960 423452 480 423542
rect 3417 423539 3483 423542
rect 198825 419386 198891 419389
rect 197126 419384 198891 419386
rect 197126 419380 198830 419384
rect 196604 419328 198830 419380
rect 198886 419328 198891 419384
rect 196604 419326 198891 419328
rect 196604 419320 197186 419326
rect 198825 419323 198891 419326
rect 356562 418842 356622 419350
rect 358813 418842 358879 418845
rect 356562 418840 358879 418842
rect 356562 418784 358818 418840
rect 358874 418784 358879 418840
rect 356562 418782 358879 418784
rect 358813 418779 358879 418782
rect 580257 418298 580323 418301
rect 583520 418298 584960 418388
rect 580257 418296 584960 418298
rect 580257 418240 580262 418296
rect 580318 418240 584960 418296
rect 580257 418238 584960 418240
rect 580257 418235 580323 418238
rect 583520 418148 584960 418238
rect 198917 417754 198983 417757
rect 197126 417752 198983 417754
rect 197126 417748 198922 417752
rect 196604 417696 198922 417748
rect 198978 417696 198983 417752
rect 196604 417694 198983 417696
rect 196604 417688 197186 417694
rect 198917 417691 198983 417694
rect 356562 417210 356622 417718
rect 358905 417210 358971 417213
rect 356562 417208 358971 417210
rect 356562 417152 358910 417208
rect 358966 417152 358971 417208
rect 356562 417150 358971 417152
rect 358905 417147 358971 417150
rect 199469 416394 199535 416397
rect 197126 416392 199535 416394
rect 197126 416388 199474 416392
rect 196604 416336 199474 416388
rect 199530 416336 199535 416392
rect 196604 416334 199535 416336
rect 196604 416328 197186 416334
rect 199469 416331 199535 416334
rect 356562 415850 356622 416358
rect 357617 415850 357683 415853
rect 356562 415848 357683 415850
rect 356562 415792 357622 415848
rect 357678 415792 357683 415848
rect 356562 415790 357683 415792
rect 357617 415787 357683 415790
rect 199377 414898 199443 414901
rect 197126 414896 199443 414898
rect 197126 414892 199382 414896
rect 196604 414840 199382 414892
rect 199438 414840 199443 414896
rect 196604 414838 199443 414840
rect 196604 414832 197186 414838
rect 199377 414835 199443 414838
rect 356562 414354 356622 414862
rect 358997 414354 359063 414357
rect 356562 414352 359063 414354
rect 356562 414296 359002 414352
rect 359058 414296 359063 414352
rect 356562 414294 359063 414296
rect 358997 414291 359063 414294
rect 197537 413674 197603 413677
rect 196942 413672 197603 413674
rect 196942 413668 197542 413672
rect 196604 413616 197542 413668
rect 197598 413616 197603 413672
rect 196604 413614 197603 413616
rect 196604 413608 197002 413614
rect 197537 413611 197603 413614
rect 356562 413130 356622 413638
rect 357525 413130 357591 413133
rect 356562 413128 357591 413130
rect 356562 413072 357530 413128
rect 357586 413072 357591 413128
rect 356562 413070 357591 413072
rect 357525 413067 357591 413070
rect -960 410546 480 410636
rect 3141 410546 3207 410549
rect -960 410544 3207 410546
rect -960 410488 3146 410544
rect 3202 410488 3207 410544
rect -960 410486 3207 410488
rect -960 410396 480 410486
rect 3141 410483 3207 410486
rect 57053 410002 57119 410005
rect 217225 410002 217291 410005
rect 57053 410000 60062 410002
rect 57053 409944 57058 410000
rect 57114 409944 60062 410000
rect 57053 409942 60062 409944
rect 217225 410000 219450 410002
rect 217225 409944 217230 410000
rect 217286 409996 219450 410000
rect 217286 409944 220064 409996
rect 217225 409942 220064 409944
rect 57053 409939 57119 409942
rect 217225 409939 217291 409942
rect 219390 409936 220064 409942
rect 57881 408234 57947 408237
rect 60002 408234 60062 408334
rect 57881 408232 60062 408234
rect 57881 408176 57886 408232
rect 57942 408176 60062 408232
rect 57881 408174 60062 408176
rect 216673 408234 216739 408237
rect 220034 408234 220094 408334
rect 216673 408232 220094 408234
rect 216673 408176 216678 408232
rect 216734 408176 220094 408232
rect 216673 408174 220094 408176
rect 57881 408171 57947 408174
rect 216673 408171 216739 408174
rect 216765 408098 216831 408101
rect 216765 408096 220094 408098
rect 56961 407554 57027 407557
rect 60002 407554 60062 408062
rect 216765 408040 216770 408096
rect 216826 408040 220094 408096
rect 216765 408038 220094 408040
rect 216765 408035 216831 408038
rect 56961 407552 60062 407554
rect 56961 407496 56966 407552
rect 57022 407496 60062 407552
rect 56961 407494 60062 407496
rect 56961 407491 57027 407494
rect 580165 404970 580231 404973
rect 583520 404970 584960 405060
rect 580165 404968 584960 404970
rect 580165 404912 580170 404968
rect 580226 404912 584960 404968
rect 580165 404910 584960 404912
rect 580165 404907 580231 404910
rect 583520 404820 584960 404910
rect 85481 398172 85547 398173
rect 85430 398170 85436 398172
rect 85390 398110 85436 398170
rect 85500 398168 85547 398172
rect 85542 398112 85547 398168
rect 85430 398108 85436 398110
rect 85500 398108 85547 398112
rect 85481 398107 85547 398108
rect 92381 398172 92447 398173
rect 95969 398172 96035 398173
rect 92381 398168 92428 398172
rect 92492 398170 92498 398172
rect 95918 398170 95924 398172
rect 92381 398112 92386 398168
rect 92381 398108 92428 398112
rect 92492 398110 92538 398170
rect 95878 398110 95924 398170
rect 95988 398168 96035 398172
rect 96030 398112 96035 398168
rect 92492 398108 92498 398110
rect 95918 398108 95924 398110
rect 95988 398108 96035 398112
rect 92381 398107 92447 398108
rect 95969 398107 96035 398108
rect 99373 398172 99439 398173
rect 113633 398172 113699 398173
rect 146017 398172 146083 398173
rect 235993 398172 236059 398173
rect 99373 398168 99420 398172
rect 99484 398170 99490 398172
rect 113582 398170 113588 398172
rect 99373 398112 99378 398168
rect 99373 398108 99420 398112
rect 99484 398110 99530 398170
rect 113542 398110 113588 398170
rect 113652 398168 113699 398172
rect 145966 398170 145972 398172
rect 113694 398112 113699 398168
rect 99484 398108 99490 398110
rect 113582 398108 113588 398110
rect 113652 398108 113699 398112
rect 145926 398110 145972 398170
rect 146036 398168 146083 398172
rect 235942 398170 235948 398172
rect 146078 398112 146083 398168
rect 145966 398108 145972 398110
rect 146036 398108 146083 398112
rect 235902 398110 235948 398170
rect 236012 398168 236059 398172
rect 236054 398112 236059 398168
rect 235942 398108 235948 398110
rect 236012 398108 236059 398112
rect 99373 398107 99439 398108
rect 113633 398107 113699 398108
rect 146017 398107 146083 398108
rect 235993 398107 236059 398108
rect 265065 398170 265131 398173
rect 265198 398170 265204 398172
rect 265065 398168 265204 398170
rect 265065 398112 265070 398168
rect 265126 398112 265204 398168
rect 265065 398110 265204 398112
rect 265065 398107 265131 398110
rect 265198 398108 265204 398110
rect 265268 398108 265274 398172
rect 300117 398170 300183 398173
rect 315757 398172 315823 398173
rect 325877 398172 325943 398173
rect 300894 398170 300900 398172
rect 300117 398168 300900 398170
rect 300117 398112 300122 398168
rect 300178 398112 300900 398168
rect 300117 398110 300900 398112
rect 300117 398107 300183 398110
rect 300894 398108 300900 398110
rect 300964 398108 300970 398172
rect 315757 398168 315804 398172
rect 315868 398170 315874 398172
rect 315757 398112 315762 398168
rect 315757 398108 315804 398112
rect 315868 398110 315914 398170
rect 325877 398168 325924 398172
rect 325988 398170 325994 398172
rect 325877 398112 325882 398168
rect 315868 398108 315874 398110
rect 325877 398108 325924 398112
rect 325988 398110 326034 398170
rect 325988 398108 325994 398110
rect 315757 398107 315823 398108
rect 325877 398107 325943 398108
rect 59077 398034 59143 398037
rect 226374 398034 226380 398036
rect 59077 398032 226380 398034
rect 59077 397976 59082 398032
rect 59138 397976 226380 398032
rect 59077 397974 226380 397976
rect 59077 397971 59143 397974
rect 226374 397972 226380 397974
rect 226444 397972 226450 398036
rect -960 397490 480 397580
rect 3417 397490 3483 397493
rect -960 397488 3483 397490
rect -960 397432 3422 397488
rect 3478 397432 3483 397488
rect -960 397430 3483 397432
rect -960 397340 480 397430
rect 3417 397427 3483 397430
rect 78305 397356 78371 397357
rect 78254 397354 78260 397356
rect 78214 397294 78260 397354
rect 78324 397352 78371 397356
rect 78366 397296 78371 397352
rect 78254 397292 78260 397294
rect 78324 397292 78371 397296
rect 80646 397292 80652 397356
rect 80716 397354 80722 397356
rect 80973 397354 81039 397357
rect 81985 397356 82051 397357
rect 81934 397354 81940 397356
rect 80716 397352 81039 397354
rect 80716 397296 80978 397352
rect 81034 397296 81039 397352
rect 80716 397294 81039 397296
rect 81894 397294 81940 397354
rect 82004 397352 82051 397356
rect 82046 397296 82051 397352
rect 80716 397292 80722 397294
rect 78305 397291 78371 397292
rect 80973 397291 81039 397294
rect 81934 397292 81940 397294
rect 82004 397292 82051 397296
rect 83222 397292 83228 397356
rect 83292 397354 83298 397356
rect 83365 397354 83431 397357
rect 83292 397352 83431 397354
rect 83292 397296 83370 397352
rect 83426 397296 83431 397352
rect 83292 397294 83431 397296
rect 83292 397292 83298 397294
rect 81985 397291 82051 397292
rect 83365 397291 83431 397294
rect 84326 397292 84332 397356
rect 84396 397354 84402 397356
rect 85021 397354 85087 397357
rect 84396 397352 85087 397354
rect 84396 397296 85026 397352
rect 85082 397296 85087 397352
rect 84396 397294 85087 397296
rect 84396 397292 84402 397294
rect 85021 397291 85087 397294
rect 87597 397356 87663 397357
rect 88793 397356 88859 397357
rect 87597 397352 87644 397356
rect 87708 397354 87714 397356
rect 88742 397354 88748 397356
rect 87597 397296 87602 397352
rect 87597 397292 87644 397296
rect 87708 397294 87754 397354
rect 88702 397294 88748 397354
rect 88812 397352 88859 397356
rect 88854 397296 88859 397352
rect 87708 397292 87714 397294
rect 88742 397292 88748 397294
rect 88812 397292 88859 397296
rect 90030 397292 90036 397356
rect 90100 397354 90106 397356
rect 90725 397354 90791 397357
rect 90100 397352 90791 397354
rect 90100 397296 90730 397352
rect 90786 397296 90791 397352
rect 90100 397294 90791 397296
rect 90100 397292 90106 397294
rect 87597 397291 87663 397292
rect 88793 397291 88859 397292
rect 90725 397291 90791 397294
rect 91277 397356 91343 397357
rect 91277 397352 91324 397356
rect 91388 397354 91394 397356
rect 94221 397354 94287 397357
rect 94446 397354 94452 397356
rect 91277 397296 91282 397352
rect 91277 397292 91324 397296
rect 91388 397294 91434 397354
rect 94221 397352 94452 397354
rect 94221 397296 94226 397352
rect 94282 397296 94452 397352
rect 94221 397294 94452 397296
rect 91388 397292 91394 397294
rect 91277 397291 91343 397292
rect 94221 397291 94287 397294
rect 94446 397292 94452 397294
rect 94516 397292 94522 397356
rect 97022 397292 97028 397356
rect 97092 397354 97098 397356
rect 97625 397354 97691 397357
rect 100753 397356 100819 397357
rect 100702 397354 100708 397356
rect 97092 397352 97691 397354
rect 97092 397296 97630 397352
rect 97686 397296 97691 397352
rect 97092 397294 97691 397296
rect 100662 397294 100708 397354
rect 100772 397352 100819 397356
rect 100814 397296 100819 397352
rect 97092 397292 97098 397294
rect 97625 397291 97691 397294
rect 100702 397292 100708 397294
rect 100772 397292 100819 397296
rect 101806 397292 101812 397356
rect 101876 397354 101882 397356
rect 102041 397354 102107 397357
rect 104065 397356 104131 397357
rect 106457 397356 106523 397357
rect 104014 397354 104020 397356
rect 101876 397352 102107 397354
rect 101876 397296 102046 397352
rect 102102 397296 102107 397352
rect 101876 397294 102107 397296
rect 103974 397294 104020 397354
rect 104084 397352 104131 397356
rect 106406 397354 106412 397356
rect 104126 397296 104131 397352
rect 101876 397292 101882 397294
rect 100753 397291 100819 397292
rect 102041 397291 102107 397294
rect 104014 397292 104020 397294
rect 104084 397292 104131 397296
rect 106366 397294 106412 397354
rect 106476 397352 106523 397356
rect 106518 397296 106523 397352
rect 106406 397292 106412 397294
rect 106476 397292 106523 397296
rect 104065 397291 104131 397292
rect 106457 397291 106523 397292
rect 109493 397356 109559 397357
rect 111241 397356 111307 397357
rect 109493 397352 109540 397356
rect 109604 397354 109610 397356
rect 111190 397354 111196 397356
rect 109493 397296 109498 397352
rect 109493 397292 109540 397296
rect 109604 397294 109650 397354
rect 111150 397294 111196 397354
rect 111260 397352 111307 397356
rect 111302 397296 111307 397352
rect 109604 397292 109610 397294
rect 111190 397292 111196 397294
rect 111260 397292 111307 397296
rect 109493 397291 109559 397292
rect 111241 397291 111307 397292
rect 112069 397356 112135 397357
rect 113173 397356 113239 397357
rect 112069 397352 112116 397356
rect 112180 397354 112186 397356
rect 112069 397296 112074 397352
rect 112069 397292 112116 397296
rect 112180 397294 112226 397354
rect 113173 397352 113220 397356
rect 113284 397354 113290 397356
rect 113725 397354 113791 397357
rect 115841 397356 115907 397357
rect 117129 397356 117195 397357
rect 114318 397354 114324 397356
rect 113173 397296 113178 397352
rect 112180 397292 112186 397294
rect 113173 397292 113220 397296
rect 113284 397294 113330 397354
rect 113725 397352 114324 397354
rect 113725 397296 113730 397352
rect 113786 397296 114324 397352
rect 113725 397294 114324 397296
rect 113284 397292 113290 397294
rect 112069 397291 112135 397292
rect 113173 397291 113239 397292
rect 113725 397291 113791 397294
rect 114318 397292 114324 397294
rect 114388 397292 114394 397356
rect 115790 397354 115796 397356
rect 115750 397294 115796 397354
rect 115860 397352 115907 397356
rect 117078 397354 117084 397356
rect 115902 397296 115907 397352
rect 115790 397292 115796 397294
rect 115860 397292 115907 397296
rect 117038 397294 117084 397354
rect 117148 397352 117195 397356
rect 117190 397296 117195 397352
rect 117078 397292 117084 397294
rect 117148 397292 117195 397296
rect 118182 397292 118188 397356
rect 118252 397354 118258 397356
rect 118325 397354 118391 397357
rect 118601 397356 118667 397357
rect 118252 397352 118391 397354
rect 118252 397296 118330 397352
rect 118386 397296 118391 397352
rect 118252 397294 118391 397296
rect 118252 397292 118258 397294
rect 115841 397291 115907 397292
rect 117129 397291 117195 397292
rect 118325 397291 118391 397294
rect 118550 397292 118556 397356
rect 118620 397354 118667 397356
rect 123477 397356 123543 397357
rect 125961 397356 126027 397357
rect 118620 397352 118712 397354
rect 118662 397296 118712 397352
rect 118620 397294 118712 397296
rect 123477 397352 123524 397356
rect 123588 397354 123594 397356
rect 125910 397354 125916 397356
rect 123477 397296 123482 397352
rect 118620 397292 118667 397294
rect 118601 397291 118667 397292
rect 123477 397292 123524 397296
rect 123588 397294 123634 397354
rect 125870 397294 125916 397354
rect 125980 397352 126027 397356
rect 126022 397296 126027 397352
rect 123588 397292 123594 397294
rect 125910 397292 125916 397294
rect 125980 397292 126027 397296
rect 136030 397292 136036 397356
rect 136100 397354 136106 397356
rect 136265 397354 136331 397357
rect 136100 397352 136331 397354
rect 136100 397296 136270 397352
rect 136326 397296 136331 397352
rect 136100 397294 136331 397296
rect 136100 397292 136106 397294
rect 123477 397291 123543 397292
rect 125961 397291 126027 397292
rect 136265 397291 136331 397294
rect 138381 397356 138447 397357
rect 138381 397352 138428 397356
rect 138492 397354 138498 397356
rect 138381 397296 138386 397352
rect 138381 397292 138428 397296
rect 138492 397294 138538 397354
rect 138492 397292 138498 397294
rect 155902 397292 155908 397356
rect 155972 397354 155978 397356
rect 156413 397354 156479 397357
rect 155972 397352 156479 397354
rect 155972 397296 156418 397352
rect 156474 397296 156479 397352
rect 155972 397294 156479 397296
rect 155972 397292 155978 397294
rect 138381 397291 138447 397292
rect 156413 397291 156479 397294
rect 163446 397292 163452 397356
rect 163516 397354 163522 397356
rect 163865 397354 163931 397357
rect 163516 397352 163931 397354
rect 163516 397296 163870 397352
rect 163926 397296 163931 397352
rect 163516 397294 163931 397296
rect 163516 397292 163522 397294
rect 163865 397291 163931 397294
rect 237005 397356 237071 397357
rect 238109 397356 238175 397357
rect 239213 397356 239279 397357
rect 240501 397356 240567 397357
rect 241605 397356 241671 397357
rect 247677 397356 247743 397357
rect 237005 397352 237052 397356
rect 237116 397354 237122 397356
rect 237005 397296 237010 397352
rect 237005 397292 237052 397296
rect 237116 397294 237162 397354
rect 238109 397352 238156 397356
rect 238220 397354 238226 397356
rect 238109 397296 238114 397352
rect 237116 397292 237122 397294
rect 238109 397292 238156 397296
rect 238220 397294 238266 397354
rect 239213 397352 239260 397356
rect 239324 397354 239330 397356
rect 239213 397296 239218 397352
rect 238220 397292 238226 397294
rect 239213 397292 239260 397296
rect 239324 397294 239370 397354
rect 240501 397352 240548 397356
rect 240612 397354 240618 397356
rect 240501 397296 240506 397352
rect 239324 397292 239330 397294
rect 240501 397292 240548 397296
rect 240612 397294 240658 397354
rect 241605 397352 241652 397356
rect 241716 397354 241722 397356
rect 241605 397296 241610 397352
rect 240612 397292 240618 397294
rect 241605 397292 241652 397296
rect 241716 397294 241762 397354
rect 247677 397352 247724 397356
rect 247788 397354 247794 397356
rect 249977 397354 250043 397357
rect 250662 397354 250668 397356
rect 247677 397296 247682 397352
rect 241716 397292 241722 397294
rect 247677 397292 247724 397296
rect 247788 397294 247834 397354
rect 249977 397352 250668 397354
rect 249977 397296 249982 397352
rect 250038 397296 250668 397352
rect 249977 397294 250668 397296
rect 247788 397292 247794 397294
rect 237005 397291 237071 397292
rect 238109 397291 238175 397292
rect 239213 397291 239279 397292
rect 240501 397291 240567 397292
rect 241605 397291 241671 397292
rect 247677 397291 247743 397292
rect 249977 397291 250043 397294
rect 250662 397292 250668 397294
rect 250732 397292 250738 397356
rect 251173 397354 251239 397357
rect 252318 397354 252324 397356
rect 251173 397352 252324 397354
rect 251173 397296 251178 397352
rect 251234 397296 252324 397352
rect 251173 397294 252324 397296
rect 251173 397291 251239 397294
rect 252318 397292 252324 397294
rect 252388 397292 252394 397356
rect 252737 397354 252803 397357
rect 253422 397354 253428 397356
rect 252737 397352 253428 397354
rect 252737 397296 252742 397352
rect 252798 397296 253428 397352
rect 252737 397294 253428 397296
rect 252737 397291 252803 397294
rect 253422 397292 253428 397294
rect 253492 397292 253498 397356
rect 259821 397354 259887 397357
rect 262029 397356 262095 397357
rect 265893 397356 265959 397357
rect 268285 397356 268351 397357
rect 270861 397356 270927 397357
rect 260598 397354 260604 397356
rect 259821 397352 260604 397354
rect 259821 397296 259826 397352
rect 259882 397296 260604 397352
rect 259821 397294 260604 397296
rect 259821 397291 259887 397294
rect 260598 397292 260604 397294
rect 260668 397292 260674 397356
rect 262029 397352 262076 397356
rect 262140 397354 262146 397356
rect 262029 397296 262034 397352
rect 262029 397292 262076 397296
rect 262140 397294 262186 397354
rect 265893 397352 265940 397356
rect 266004 397354 266010 397356
rect 265893 397296 265898 397352
rect 262140 397292 262146 397294
rect 265893 397292 265940 397296
rect 266004 397294 266050 397354
rect 268285 397352 268332 397356
rect 268396 397354 268402 397356
rect 268285 397296 268290 397352
rect 266004 397292 266010 397294
rect 268285 397292 268332 397296
rect 268396 397294 268442 397354
rect 270861 397352 270908 397356
rect 270972 397354 270978 397356
rect 272241 397354 272307 397357
rect 272558 397354 272564 397356
rect 270861 397296 270866 397352
rect 268396 397292 268402 397294
rect 270861 397292 270908 397296
rect 270972 397294 271018 397354
rect 272241 397352 272564 397354
rect 272241 397296 272246 397352
rect 272302 397296 272564 397352
rect 272241 397294 272564 397296
rect 270972 397292 270978 397294
rect 262029 397291 262095 397292
rect 265893 397291 265959 397292
rect 268285 397291 268351 397292
rect 270861 397291 270927 397292
rect 272241 397291 272307 397294
rect 272558 397292 272564 397294
rect 272628 397292 272634 397356
rect 273437 397354 273503 397357
rect 276197 397356 276263 397357
rect 274398 397354 274404 397356
rect 273437 397352 274404 397354
rect 273437 397296 273442 397352
rect 273498 397296 274404 397352
rect 273437 397294 274404 397296
rect 273437 397291 273503 397294
rect 274398 397292 274404 397294
rect 274468 397292 274474 397356
rect 276197 397354 276244 397356
rect 276152 397352 276244 397354
rect 276152 397296 276202 397352
rect 276152 397294 276244 397296
rect 276197 397292 276244 397294
rect 276308 397292 276314 397356
rect 276381 397354 276447 397357
rect 278037 397356 278103 397357
rect 278957 397356 279023 397357
rect 276974 397354 276980 397356
rect 276381 397352 276980 397354
rect 276381 397296 276386 397352
rect 276442 397296 276980 397352
rect 276381 397294 276980 397296
rect 276197 397291 276263 397292
rect 276381 397291 276447 397294
rect 276974 397292 276980 397294
rect 277044 397292 277050 397356
rect 278037 397352 278084 397356
rect 278148 397354 278154 397356
rect 278037 397296 278042 397352
rect 278037 397292 278084 397296
rect 278148 397294 278194 397354
rect 278957 397352 279004 397356
rect 279068 397354 279074 397356
rect 283189 397354 283255 397357
rect 283782 397354 283788 397356
rect 278957 397296 278962 397352
rect 278148 397292 278154 397294
rect 278957 397292 279004 397296
rect 279068 397294 279114 397354
rect 283189 397352 283788 397354
rect 283189 397296 283194 397352
rect 283250 397296 283788 397352
rect 283189 397294 283788 397296
rect 279068 397292 279074 397294
rect 278037 397291 278103 397292
rect 278957 397291 279023 397292
rect 283189 397291 283255 397294
rect 283782 397292 283788 397294
rect 283852 397292 283858 397356
rect 289813 397354 289879 397357
rect 298461 397356 298527 397357
rect 343357 397356 343423 397357
rect 290958 397354 290964 397356
rect 289813 397352 290964 397354
rect 289813 397296 289818 397352
rect 289874 397296 290964 397352
rect 289813 397294 290964 397296
rect 289813 397291 289879 397294
rect 290958 397292 290964 397294
rect 291028 397292 291034 397356
rect 298461 397352 298508 397356
rect 298572 397354 298578 397356
rect 298461 397296 298466 397352
rect 298461 397292 298508 397296
rect 298572 397294 298618 397354
rect 343357 397352 343404 397356
rect 343468 397354 343474 397356
rect 343357 397296 343362 397352
rect 298572 397292 298578 397294
rect 343357 397292 343404 397296
rect 343468 397294 343514 397354
rect 343468 397292 343474 397294
rect 298461 397291 298527 397292
rect 343357 397291 343423 397292
rect 251265 397220 251331 397221
rect 251214 397218 251220 397220
rect 251174 397158 251220 397218
rect 251284 397216 251331 397220
rect 251326 397160 251331 397216
rect 251214 397156 251220 397158
rect 251284 397156 251331 397160
rect 251265 397155 251331 397156
rect 273345 397218 273411 397221
rect 273478 397218 273484 397220
rect 273345 397216 273484 397218
rect 273345 397160 273350 397216
rect 273406 397160 273484 397216
rect 273345 397158 273484 397160
rect 273345 397155 273411 397158
rect 273478 397156 273484 397158
rect 273548 397156 273554 397220
rect 258073 396946 258139 396949
rect 258390 396946 258396 396948
rect 258073 396944 258396 396946
rect 258073 396888 258078 396944
rect 258134 396888 258396 396944
rect 258073 396886 258396 396888
rect 258073 396883 258139 396886
rect 258390 396884 258396 396886
rect 258460 396884 258466 396948
rect 77201 396812 77267 396813
rect 77150 396810 77156 396812
rect 77110 396750 77156 396810
rect 77220 396808 77267 396812
rect 77262 396752 77267 396808
rect 77150 396748 77156 396750
rect 77220 396748 77267 396752
rect 77201 396747 77267 396748
rect 78765 396810 78831 396813
rect 79542 396810 79548 396812
rect 78765 396808 79548 396810
rect 78765 396752 78770 396808
rect 78826 396752 79548 396808
rect 78765 396750 79548 396752
rect 78765 396747 78831 396750
rect 79542 396748 79548 396750
rect 79612 396748 79618 396812
rect 86534 396748 86540 396812
rect 86604 396810 86610 396812
rect 86861 396810 86927 396813
rect 86604 396808 86927 396810
rect 86604 396752 86866 396808
rect 86922 396752 86927 396808
rect 86604 396750 86927 396752
rect 86604 396748 86610 396750
rect 86861 396747 86927 396750
rect 88333 396812 88399 396813
rect 88333 396808 88380 396812
rect 88444 396810 88450 396812
rect 88333 396752 88338 396808
rect 88333 396748 88380 396752
rect 88444 396750 88490 396810
rect 88444 396748 88450 396750
rect 90766 396748 90772 396812
rect 90836 396810 90842 396812
rect 91001 396810 91067 396813
rect 90836 396808 91067 396810
rect 90836 396752 91006 396808
rect 91062 396752 91067 396808
rect 90836 396750 91067 396752
rect 90836 396748 90842 396750
rect 88333 396747 88399 396748
rect 91001 396747 91067 396750
rect 93669 396812 93735 396813
rect 96337 396812 96403 396813
rect 93669 396808 93716 396812
rect 93780 396810 93786 396812
rect 96286 396810 96292 396812
rect 93669 396752 93674 396808
rect 93669 396748 93716 396752
rect 93780 396750 93826 396810
rect 96246 396750 96292 396810
rect 96356 396808 96403 396812
rect 96398 396752 96403 396808
rect 93780 396748 93786 396750
rect 96286 396748 96292 396750
rect 96356 396748 96403 396752
rect 98494 396748 98500 396812
rect 98564 396810 98570 396812
rect 99189 396810 99255 396813
rect 98564 396808 99255 396810
rect 98564 396752 99194 396808
rect 99250 396752 99255 396808
rect 98564 396750 99255 396752
rect 98564 396748 98570 396750
rect 93669 396747 93735 396748
rect 96337 396747 96403 396748
rect 99189 396747 99255 396750
rect 101070 396748 101076 396812
rect 101140 396810 101146 396812
rect 101949 396810 102015 396813
rect 101140 396808 102015 396810
rect 101140 396752 101954 396808
rect 102010 396752 102015 396808
rect 101140 396750 102015 396752
rect 101140 396748 101146 396750
rect 101949 396747 102015 396750
rect 102726 396748 102732 396812
rect 102796 396810 102802 396812
rect 103421 396810 103487 396813
rect 102796 396808 103487 396810
rect 102796 396752 103426 396808
rect 103482 396752 103487 396808
rect 102796 396750 103487 396752
rect 102796 396748 102802 396750
rect 103421 396747 103487 396750
rect 103830 396748 103836 396812
rect 103900 396810 103906 396812
rect 104709 396810 104775 396813
rect 103900 396808 104775 396810
rect 103900 396752 104714 396808
rect 104770 396752 104775 396808
rect 103900 396750 104775 396752
rect 103900 396748 103906 396750
rect 104709 396747 104775 396750
rect 105302 396748 105308 396812
rect 105372 396810 105378 396812
rect 105721 396810 105787 396813
rect 106089 396812 106155 396813
rect 107561 396812 107627 396813
rect 106038 396810 106044 396812
rect 105372 396808 105787 396810
rect 105372 396752 105726 396808
rect 105782 396752 105787 396808
rect 105372 396750 105787 396752
rect 105998 396750 106044 396810
rect 106108 396808 106155 396812
rect 107510 396810 107516 396812
rect 106150 396752 106155 396808
rect 105372 396748 105378 396750
rect 105721 396747 105787 396750
rect 106038 396748 106044 396750
rect 106108 396748 106155 396752
rect 107470 396750 107516 396810
rect 107580 396808 107627 396812
rect 107622 396752 107627 396808
rect 107510 396748 107516 396750
rect 107580 396748 107627 396752
rect 108798 396748 108804 396812
rect 108868 396810 108874 396812
rect 108941 396810 109007 396813
rect 108868 396808 109007 396810
rect 108868 396752 108946 396808
rect 109002 396752 109007 396808
rect 108868 396750 109007 396752
rect 108868 396748 108874 396750
rect 106089 396747 106155 396748
rect 107561 396747 107627 396748
rect 108941 396747 109007 396750
rect 111006 396748 111012 396812
rect 111076 396810 111082 396812
rect 111701 396810 111767 396813
rect 111076 396808 111767 396810
rect 111076 396752 111706 396808
rect 111762 396752 111767 396808
rect 111076 396750 111767 396752
rect 111076 396748 111082 396750
rect 111701 396747 111767 396750
rect 115974 396748 115980 396812
rect 116044 396810 116050 396812
rect 117037 396810 117103 396813
rect 116044 396808 117103 396810
rect 116044 396752 117042 396808
rect 117098 396752 117103 396808
rect 116044 396750 117103 396752
rect 116044 396748 116050 396750
rect 117037 396747 117103 396750
rect 119102 396748 119108 396812
rect 119172 396810 119178 396812
rect 119889 396810 119955 396813
rect 119172 396808 119955 396810
rect 119172 396752 119894 396808
rect 119950 396752 119955 396808
rect 119172 396750 119955 396752
rect 119172 396748 119178 396750
rect 119889 396747 119955 396750
rect 120073 396810 120139 396813
rect 120758 396810 120764 396812
rect 120073 396808 120764 396810
rect 120073 396752 120078 396808
rect 120134 396752 120764 396808
rect 120073 396750 120764 396752
rect 120073 396747 120139 396750
rect 120758 396748 120764 396750
rect 120828 396748 120834 396812
rect 129733 396810 129799 396813
rect 130878 396810 130884 396812
rect 129733 396808 130884 396810
rect 129733 396752 129738 396808
rect 129794 396752 130884 396808
rect 129733 396750 130884 396752
rect 129733 396747 129799 396750
rect 130878 396748 130884 396750
rect 130948 396748 130954 396812
rect 133454 396748 133460 396812
rect 133524 396810 133530 396812
rect 133781 396810 133847 396813
rect 133524 396808 133847 396810
rect 133524 396752 133786 396808
rect 133842 396752 133847 396808
rect 133524 396750 133847 396752
rect 133524 396748 133530 396750
rect 133781 396747 133847 396750
rect 140773 396812 140839 396813
rect 140773 396808 140820 396812
rect 140884 396810 140890 396812
rect 140773 396752 140778 396808
rect 140773 396748 140820 396752
rect 140884 396750 140930 396810
rect 140884 396748 140890 396750
rect 143574 396748 143580 396812
rect 143644 396810 143650 396812
rect 144821 396810 144887 396813
rect 143644 396808 144887 396810
rect 143644 396752 144826 396808
rect 144882 396752 144887 396808
rect 143644 396750 144887 396752
rect 143644 396748 143650 396750
rect 140773 396747 140839 396748
rect 144821 396747 144887 396750
rect 147673 396810 147739 396813
rect 148542 396810 148548 396812
rect 147673 396808 148548 396810
rect 147673 396752 147678 396808
rect 147734 396752 148548 396808
rect 147673 396750 148548 396752
rect 147673 396747 147739 396750
rect 148542 396748 148548 396750
rect 148612 396748 148618 396812
rect 150934 396748 150940 396812
rect 151004 396810 151010 396812
rect 151721 396810 151787 396813
rect 151004 396808 151787 396810
rect 151004 396752 151726 396808
rect 151782 396752 151787 396808
rect 151004 396750 151787 396752
rect 151004 396748 151010 396750
rect 151721 396747 151787 396750
rect 154062 396748 154068 396812
rect 154132 396810 154138 396812
rect 154481 396810 154547 396813
rect 154132 396808 154547 396810
rect 154132 396752 154486 396808
rect 154542 396752 154547 396808
rect 154132 396750 154547 396752
rect 154132 396748 154138 396750
rect 154481 396747 154547 396750
rect 158478 396748 158484 396812
rect 158548 396810 158554 396812
rect 158621 396810 158687 396813
rect 158548 396808 158687 396810
rect 158548 396752 158626 396808
rect 158682 396752 158687 396808
rect 158548 396750 158687 396752
rect 158548 396748 158554 396750
rect 158621 396747 158687 396750
rect 160870 396748 160876 396812
rect 160940 396810 160946 396812
rect 161381 396810 161447 396813
rect 160940 396808 161447 396810
rect 160940 396752 161386 396808
rect 161442 396752 161447 396808
rect 160940 396750 161447 396752
rect 160940 396748 160946 396750
rect 161381 396747 161447 396750
rect 165613 396810 165679 396813
rect 165838 396810 165844 396812
rect 165613 396808 165844 396810
rect 165613 396752 165618 396808
rect 165674 396752 165844 396808
rect 165613 396750 165844 396752
rect 165613 396747 165679 396750
rect 165838 396748 165844 396750
rect 165908 396748 165914 396812
rect 182173 396810 182239 396813
rect 183461 396812 183527 396813
rect 242893 396812 242959 396813
rect 183134 396810 183140 396812
rect 182173 396808 183140 396810
rect 182173 396752 182178 396808
rect 182234 396752 183140 396808
rect 182173 396750 183140 396752
rect 182173 396747 182239 396750
rect 183134 396748 183140 396750
rect 183204 396748 183210 396812
rect 183461 396808 183508 396812
rect 183572 396810 183578 396812
rect 183461 396752 183466 396808
rect 183461 396748 183508 396752
rect 183572 396750 183618 396810
rect 242893 396808 242940 396812
rect 243004 396810 243010 396812
rect 242893 396752 242898 396808
rect 183572 396748 183578 396750
rect 242893 396748 242940 396752
rect 243004 396750 243050 396810
rect 243004 396748 243010 396750
rect 244222 396748 244228 396812
rect 244292 396810 244298 396812
rect 244365 396810 244431 396813
rect 244292 396808 244431 396810
rect 244292 396752 244370 396808
rect 244426 396752 244431 396808
rect 244292 396750 244431 396752
rect 244292 396748 244298 396750
rect 183461 396747 183527 396748
rect 242893 396747 242959 396748
rect 244365 396747 244431 396750
rect 245653 396810 245719 396813
rect 246430 396810 246436 396812
rect 245653 396808 246436 396810
rect 245653 396752 245658 396808
rect 245714 396752 246436 396808
rect 245653 396750 246436 396752
rect 245653 396747 245719 396750
rect 246430 396748 246436 396750
rect 246500 396748 246506 396812
rect 247585 396810 247651 396813
rect 248270 396810 248276 396812
rect 247585 396808 248276 396810
rect 247585 396752 247590 396808
rect 247646 396752 248276 396808
rect 247585 396750 248276 396752
rect 247585 396747 247651 396750
rect 248270 396748 248276 396750
rect 248340 396748 248346 396812
rect 248413 396810 248479 396813
rect 248638 396810 248644 396812
rect 248413 396808 248644 396810
rect 248413 396752 248418 396808
rect 248474 396752 248644 396808
rect 248413 396750 248644 396752
rect 248413 396747 248479 396750
rect 248638 396748 248644 396750
rect 248708 396748 248714 396812
rect 249793 396810 249859 396813
rect 250110 396810 250116 396812
rect 249793 396808 250116 396810
rect 249793 396752 249798 396808
rect 249854 396752 250116 396808
rect 249793 396750 250116 396752
rect 249793 396747 249859 396750
rect 250110 396748 250116 396750
rect 250180 396748 250186 396812
rect 252645 396810 252711 396813
rect 254485 396812 254551 396813
rect 253606 396810 253612 396812
rect 252645 396808 253612 396810
rect 252645 396752 252650 396808
rect 252706 396752 253612 396808
rect 252645 396750 253612 396752
rect 252645 396747 252711 396750
rect 253606 396748 253612 396750
rect 253676 396748 253682 396812
rect 254485 396808 254532 396812
rect 254596 396810 254602 396812
rect 255405 396810 255471 396813
rect 256877 396812 256943 396813
rect 255814 396810 255820 396812
rect 254485 396752 254490 396808
rect 254485 396748 254532 396752
rect 254596 396750 254642 396810
rect 255405 396808 255820 396810
rect 255405 396752 255410 396808
rect 255466 396752 255820 396808
rect 255405 396750 255820 396752
rect 254596 396748 254602 396750
rect 254485 396747 254551 396748
rect 255405 396747 255471 396750
rect 255814 396748 255820 396750
rect 255884 396748 255890 396812
rect 256877 396808 256924 396812
rect 256988 396810 256994 396812
rect 258165 396810 258231 396813
rect 259545 396812 259611 396813
rect 258390 396810 258396 396812
rect 256877 396752 256882 396808
rect 256877 396748 256924 396752
rect 256988 396750 257034 396810
rect 258165 396808 258396 396810
rect 258165 396752 258170 396808
rect 258226 396752 258396 396808
rect 258165 396750 258396 396752
rect 256988 396748 256994 396750
rect 256877 396747 256943 396748
rect 258165 396747 258231 396750
rect 258390 396748 258396 396750
rect 258460 396748 258466 396812
rect 259494 396810 259500 396812
rect 259454 396750 259500 396810
rect 259564 396808 259611 396812
rect 259606 396752 259611 396808
rect 259494 396748 259500 396750
rect 259564 396748 259611 396752
rect 259545 396747 259611 396748
rect 260925 396812 260991 396813
rect 260925 396808 260972 396812
rect 261036 396810 261042 396812
rect 262213 396810 262279 396813
rect 263593 396812 263659 396813
rect 266353 396812 266419 396813
rect 262806 396810 262812 396812
rect 260925 396752 260930 396808
rect 260925 396748 260972 396752
rect 261036 396750 261082 396810
rect 262213 396808 262812 396810
rect 262213 396752 262218 396808
rect 262274 396752 262812 396808
rect 262213 396750 262812 396752
rect 261036 396748 261042 396750
rect 260925 396747 260991 396748
rect 262213 396747 262279 396750
rect 262806 396748 262812 396750
rect 262876 396748 262882 396812
rect 263542 396810 263548 396812
rect 263502 396750 263548 396810
rect 263612 396808 263659 396812
rect 266302 396810 266308 396812
rect 263654 396752 263659 396808
rect 263542 396748 263548 396750
rect 263612 396748 263659 396752
rect 266262 396750 266308 396810
rect 266372 396808 266419 396812
rect 266414 396752 266419 396808
rect 266302 396748 266308 396750
rect 266372 396748 266419 396752
rect 263593 396747 263659 396748
rect 266353 396747 266419 396748
rect 267825 396810 267891 396813
rect 268694 396810 268700 396812
rect 267825 396808 268700 396810
rect 267825 396752 267830 396808
rect 267886 396752 268700 396808
rect 267825 396750 268700 396752
rect 267825 396747 267891 396750
rect 268694 396748 268700 396750
rect 268764 396748 268770 396812
rect 269113 396810 269179 396813
rect 269798 396810 269804 396812
rect 269113 396808 269804 396810
rect 269113 396752 269118 396808
rect 269174 396752 269804 396808
rect 269113 396750 269804 396752
rect 269113 396747 269179 396750
rect 269798 396748 269804 396750
rect 269868 396748 269874 396812
rect 270585 396810 270651 396813
rect 273253 396812 273319 396813
rect 271270 396810 271276 396812
rect 270585 396808 271276 396810
rect 270585 396752 270590 396808
rect 270646 396752 271276 396808
rect 270585 396750 271276 396752
rect 270585 396747 270651 396750
rect 271270 396748 271276 396750
rect 271340 396748 271346 396812
rect 273253 396808 273300 396812
rect 273364 396810 273370 396812
rect 274633 396810 274699 396813
rect 275318 396810 275324 396812
rect 273253 396752 273258 396808
rect 273253 396748 273300 396752
rect 273364 396750 273410 396810
rect 274633 396808 275324 396810
rect 274633 396752 274638 396808
rect 274694 396752 275324 396808
rect 274633 396750 275324 396752
rect 273364 396748 273370 396750
rect 273253 396747 273319 396748
rect 274633 396747 274699 396750
rect 275318 396748 275324 396750
rect 275388 396748 275394 396812
rect 277485 396810 277551 396813
rect 278446 396810 278452 396812
rect 277485 396808 278452 396810
rect 277485 396752 277490 396808
rect 277546 396752 278452 396808
rect 277485 396750 278452 396752
rect 277485 396747 277551 396750
rect 278446 396748 278452 396750
rect 278516 396748 278522 396812
rect 280153 396810 280219 396813
rect 280838 396810 280844 396812
rect 280153 396808 280844 396810
rect 280153 396752 280158 396808
rect 280214 396752 280844 396808
rect 280153 396750 280844 396752
rect 280153 396747 280219 396750
rect 280838 396748 280844 396750
rect 280908 396748 280914 396812
rect 285673 396810 285739 396813
rect 285990 396810 285996 396812
rect 285673 396808 285996 396810
rect 285673 396752 285678 396808
rect 285734 396752 285996 396808
rect 285673 396750 285996 396752
rect 285673 396747 285739 396750
rect 285990 396748 285996 396750
rect 286060 396748 286066 396812
rect 287053 396810 287119 396813
rect 288198 396810 288204 396812
rect 287053 396808 288204 396810
rect 287053 396752 287058 396808
rect 287114 396752 288204 396808
rect 287053 396750 288204 396752
rect 287053 396747 287119 396750
rect 288198 396748 288204 396750
rect 288268 396748 288274 396812
rect 292941 396810 293007 396813
rect 295885 396812 295951 396813
rect 293350 396810 293356 396812
rect 292941 396808 293356 396810
rect 292941 396752 292946 396808
rect 293002 396752 293356 396808
rect 292941 396750 293356 396752
rect 292941 396747 293007 396750
rect 293350 396748 293356 396750
rect 293420 396748 293426 396812
rect 295885 396808 295932 396812
rect 295996 396810 296002 396812
rect 302233 396810 302299 396813
rect 303470 396810 303476 396812
rect 295885 396752 295890 396808
rect 295885 396748 295932 396752
rect 295996 396750 296042 396810
rect 302233 396808 303476 396810
rect 302233 396752 302238 396808
rect 302294 396752 303476 396808
rect 302233 396750 303476 396752
rect 295996 396748 296002 396750
rect 295885 396747 295951 396748
rect 302233 396747 302299 396750
rect 303470 396748 303476 396750
rect 303540 396748 303546 396812
rect 305269 396810 305335 396813
rect 305862 396810 305868 396812
rect 305269 396808 305868 396810
rect 305269 396752 305274 396808
rect 305330 396752 305868 396808
rect 305269 396750 305868 396752
rect 305269 396747 305335 396750
rect 305862 396748 305868 396750
rect 305932 396748 305938 396812
rect 307845 396810 307911 396813
rect 308622 396810 308628 396812
rect 307845 396808 308628 396810
rect 307845 396752 307850 396808
rect 307906 396752 308628 396808
rect 307845 396750 308628 396752
rect 307845 396747 307911 396750
rect 308622 396748 308628 396750
rect 308692 396748 308698 396812
rect 310513 396810 310579 396813
rect 311014 396810 311020 396812
rect 310513 396808 311020 396810
rect 310513 396752 310518 396808
rect 310574 396752 311020 396808
rect 310513 396750 311020 396752
rect 310513 396747 310579 396750
rect 311014 396748 311020 396750
rect 311084 396748 311090 396812
rect 313273 396810 313339 396813
rect 313406 396810 313412 396812
rect 313273 396808 313412 396810
rect 313273 396752 313278 396808
rect 313334 396752 313412 396808
rect 313273 396750 313412 396752
rect 313273 396747 313339 396750
rect 313406 396748 313412 396750
rect 313476 396748 313482 396812
rect 317413 396810 317479 396813
rect 318374 396810 318380 396812
rect 317413 396808 318380 396810
rect 317413 396752 317418 396808
rect 317474 396752 318380 396808
rect 317413 396750 318380 396752
rect 317413 396747 317479 396750
rect 318374 396748 318380 396750
rect 318444 396748 318450 396812
rect 320173 396810 320239 396813
rect 320950 396810 320956 396812
rect 320173 396808 320956 396810
rect 320173 396752 320178 396808
rect 320234 396752 320956 396808
rect 320173 396750 320956 396752
rect 320173 396747 320239 396750
rect 320950 396748 320956 396750
rect 321020 396748 321026 396812
rect 323117 396810 323183 396813
rect 323342 396810 323348 396812
rect 323117 396808 323348 396810
rect 323117 396752 323122 396808
rect 323178 396752 323348 396808
rect 323117 396750 323348 396752
rect 323117 396747 323183 396750
rect 323342 396748 323348 396750
rect 323412 396748 323418 396812
rect 342345 396810 342411 396813
rect 343214 396810 343220 396812
rect 342345 396808 343220 396810
rect 342345 396752 342350 396808
rect 342406 396752 343220 396808
rect 342345 396750 343220 396752
rect 342345 396747 342411 396750
rect 343214 396748 343220 396750
rect 343284 396748 343290 396812
rect 76046 396612 76052 396676
rect 76116 396674 76122 396676
rect 77109 396674 77175 396677
rect 76116 396672 77175 396674
rect 76116 396616 77114 396672
rect 77170 396616 77175 396672
rect 76116 396614 77175 396616
rect 76116 396612 76122 396614
rect 77109 396611 77175 396614
rect 93342 396612 93348 396676
rect 93412 396674 93418 396676
rect 93761 396674 93827 396677
rect 93412 396672 93827 396674
rect 93412 396616 93766 396672
rect 93822 396616 93827 396672
rect 93412 396614 93827 396616
rect 93412 396612 93418 396614
rect 93761 396611 93827 396614
rect 98126 396612 98132 396676
rect 98196 396674 98202 396676
rect 99281 396674 99347 396677
rect 98196 396672 99347 396674
rect 98196 396616 99286 396672
rect 99342 396616 99347 396672
rect 98196 396614 99347 396616
rect 98196 396612 98202 396614
rect 99281 396611 99347 396614
rect 108246 396612 108252 396676
rect 108316 396674 108322 396676
rect 108849 396674 108915 396677
rect 108316 396672 108915 396674
rect 108316 396616 108854 396672
rect 108910 396616 108915 396672
rect 108316 396614 108915 396616
rect 108316 396612 108322 396614
rect 108849 396611 108915 396614
rect 244273 396674 244339 396677
rect 245326 396674 245332 396676
rect 244273 396672 245332 396674
rect 244273 396616 244278 396672
rect 244334 396616 245332 396672
rect 244273 396614 245332 396616
rect 244273 396611 244339 396614
rect 245326 396612 245332 396614
rect 245396 396612 245402 396676
rect 255313 396674 255379 396677
rect 256182 396674 256188 396676
rect 255313 396672 256188 396674
rect 255313 396616 255318 396672
rect 255374 396616 256188 396672
rect 255313 396614 256188 396616
rect 255313 396611 255379 396614
rect 256182 396612 256188 396614
rect 256252 396612 256258 396676
rect 263685 396674 263751 396677
rect 263910 396674 263916 396676
rect 263685 396672 263916 396674
rect 263685 396616 263690 396672
rect 263746 396616 263916 396672
rect 263685 396614 263916 396616
rect 263685 396611 263751 396614
rect 263910 396612 263916 396614
rect 263980 396612 263986 396676
rect 266445 396674 266511 396677
rect 267590 396674 267596 396676
rect 266445 396672 267596 396674
rect 266445 396616 266450 396672
rect 266506 396616 267596 396672
rect 266445 396614 267596 396616
rect 266445 396611 266511 396614
rect 267590 396612 267596 396614
rect 267660 396612 267666 396676
rect 128670 396068 128676 396132
rect 128740 396130 128746 396132
rect 129641 396130 129707 396133
rect 128740 396128 129707 396130
rect 128740 396072 129646 396128
rect 129702 396072 129707 396128
rect 128740 396070 129707 396072
rect 128740 396068 128746 396070
rect 129641 396067 129707 396070
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 580165 378450 580231 378453
rect 583520 378450 584960 378540
rect 580165 378448 584960 378450
rect 580165 378392 580170 378448
rect 580226 378392 584960 378448
rect 580165 378390 584960 378392
rect 580165 378387 580231 378390
rect 583520 378300 584960 378390
rect -960 371378 480 371468
rect 3417 371378 3483 371381
rect -960 371376 3483 371378
rect -960 371320 3422 371376
rect 3478 371320 3483 371376
rect -960 371318 3483 371320
rect -960 371228 480 371318
rect 3417 371315 3483 371318
rect 579613 365122 579679 365125
rect 583520 365122 584960 365212
rect 579613 365120 584960 365122
rect 579613 365064 579618 365120
rect 579674 365064 584960 365120
rect 579613 365062 584960 365064
rect 579613 365059 579679 365062
rect 583520 364972 584960 365062
rect -960 358458 480 358548
rect 3141 358458 3207 358461
rect -960 358456 3207 358458
rect -960 358400 3146 358456
rect 3202 358400 3207 358456
rect -960 358398 3207 358400
rect -960 358308 480 358398
rect 3141 358395 3207 358398
rect 580165 351930 580231 351933
rect 583520 351930 584960 352020
rect 580165 351928 584960 351930
rect 580165 351872 580170 351928
rect 580226 351872 584960 351928
rect 580165 351870 584960 351872
rect 580165 351867 580231 351870
rect 583520 351780 584960 351870
rect -960 345402 480 345492
rect 3325 345402 3391 345405
rect -960 345400 3391 345402
rect -960 345344 3330 345400
rect 3386 345344 3391 345400
rect -960 345342 3391 345344
rect -960 345252 480 345342
rect 3325 345339 3391 345342
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 580165 325274 580231 325277
rect 583520 325274 584960 325364
rect 580165 325272 584960 325274
rect 580165 325216 580170 325272
rect 580226 325216 584960 325272
rect 580165 325214 584960 325216
rect 580165 325211 580231 325214
rect 583520 325124 584960 325214
rect -960 319290 480 319380
rect 3417 319290 3483 319293
rect -960 319288 3483 319290
rect -960 319232 3422 319288
rect 3478 319232 3483 319288
rect -960 319230 3483 319232
rect -960 319140 480 319230
rect 3417 319227 3483 319230
rect 579981 312082 580047 312085
rect 583520 312082 584960 312172
rect 579981 312080 584960 312082
rect 579981 312024 579986 312080
rect 580042 312024 584960 312080
rect 579981 312022 584960 312024
rect 579981 312019 580047 312022
rect 583520 311932 584960 312022
rect -960 306234 480 306324
rect 3233 306234 3299 306237
rect -960 306232 3299 306234
rect -960 306176 3238 306232
rect 3294 306176 3299 306232
rect -960 306174 3299 306176
rect -960 306084 480 306174
rect 3233 306171 3299 306174
rect 580165 298754 580231 298757
rect 583520 298754 584960 298844
rect 580165 298752 584960 298754
rect 580165 298696 580170 298752
rect 580226 298696 584960 298752
rect 580165 298694 584960 298696
rect 580165 298691 580231 298694
rect 583520 298604 584960 298694
rect -960 293178 480 293268
rect 3417 293178 3483 293181
rect -960 293176 3483 293178
rect -960 293120 3422 293176
rect 3478 293120 3483 293176
rect -960 293118 3483 293120
rect -960 293028 480 293118
rect 3417 293115 3483 293118
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 580165 272234 580231 272237
rect 583520 272234 584960 272324
rect 580165 272232 584960 272234
rect 580165 272176 580170 272232
rect 580226 272176 584960 272232
rect 580165 272174 584960 272176
rect 580165 272171 580231 272174
rect 583520 272084 584960 272174
rect -960 267202 480 267292
rect 3049 267202 3115 267205
rect -960 267200 3115 267202
rect -960 267144 3054 267200
rect 3110 267144 3115 267200
rect -960 267142 3115 267144
rect -960 267052 480 267142
rect 3049 267139 3115 267142
rect 580165 258906 580231 258909
rect 583520 258906 584960 258996
rect 580165 258904 584960 258906
rect 580165 258848 580170 258904
rect 580226 258848 584960 258904
rect 580165 258846 584960 258848
rect 580165 258843 580231 258846
rect 583520 258756 584960 258846
rect -960 254146 480 254236
rect 3417 254146 3483 254149
rect -960 254144 3483 254146
rect -960 254088 3422 254144
rect 3478 254088 3483 254144
rect -960 254086 3483 254088
rect -960 253996 480 254086
rect 3417 254083 3483 254086
rect 579797 245578 579863 245581
rect 583520 245578 584960 245668
rect 579797 245576 584960 245578
rect 579797 245520 579802 245576
rect 579858 245520 584960 245576
rect 579797 245518 584960 245520
rect 579797 245515 579863 245518
rect 583520 245428 584960 245518
rect 57237 242178 57303 242181
rect 226742 242178 226748 242180
rect 57237 242176 226748 242178
rect 57237 242120 57242 242176
rect 57298 242120 226748 242176
rect 57237 242118 226748 242120
rect 57237 242115 57303 242118
rect 226742 242116 226748 242118
rect 226812 242116 226818 242180
rect -960 241090 480 241180
rect 3417 241090 3483 241093
rect -960 241088 3483 241090
rect -960 241032 3422 241088
rect 3478 241032 3483 241088
rect -960 241030 3483 241032
rect -960 240940 480 241030
rect 3417 241027 3483 241030
rect 121269 237962 121335 237965
rect 135897 237962 135963 237965
rect 121269 237960 135963 237962
rect 121269 237904 121274 237960
rect 121330 237904 135902 237960
rect 135958 237904 135963 237960
rect 121269 237902 135963 237904
rect 121269 237899 121335 237902
rect 135897 237899 135963 237902
rect 76925 236058 76991 236061
rect 228398 236058 228404 236060
rect 76925 236056 228404 236058
rect 76925 236000 76930 236056
rect 76986 236000 228404 236056
rect 76925 235998 228404 236000
rect 76925 235995 76991 235998
rect 228398 235996 228404 235998
rect 228468 235996 228474 236060
rect 215569 235242 215635 235245
rect 227069 235242 227135 235245
rect 215569 235240 227135 235242
rect 215569 235184 215574 235240
rect 215630 235184 227074 235240
rect 227130 235184 227135 235240
rect 215569 235182 227135 235184
rect 215569 235179 215635 235182
rect 227069 235179 227135 235182
rect 33777 234834 33843 234837
rect 167361 234834 167427 234837
rect 33777 234832 167427 234834
rect 33777 234776 33782 234832
rect 33838 234776 167366 234832
rect 167422 234776 167427 234832
rect 33777 234774 167427 234776
rect 33777 234771 33843 234774
rect 167361 234771 167427 234774
rect 74165 234698 74231 234701
rect 231209 234698 231275 234701
rect 74165 234696 231275 234698
rect 74165 234640 74170 234696
rect 74226 234640 231214 234696
rect 231270 234640 231275 234696
rect 74165 234638 231275 234640
rect 74165 234635 74231 234638
rect 231209 234635 231275 234638
rect 129733 234018 129799 234021
rect 130377 234018 130443 234021
rect 129733 234016 130443 234018
rect 129733 233960 129738 234016
rect 129794 233960 130382 234016
rect 130438 233960 130443 234016
rect 129733 233958 130443 233960
rect 129733 233955 129799 233958
rect 130377 233955 130443 233958
rect 132493 234018 132559 234021
rect 133137 234018 133203 234021
rect 132493 234016 133203 234018
rect 132493 233960 132498 234016
rect 132554 233960 133142 234016
rect 133198 233960 133203 234016
rect 132493 233958 133203 233960
rect 132493 233955 132559 233958
rect 133137 233955 133203 233958
rect 106917 233882 106983 233885
rect 152273 233882 152339 233885
rect 106917 233880 152339 233882
rect 106917 233824 106922 233880
rect 106978 233824 152278 233880
rect 152334 233824 152339 233880
rect 106917 233822 152339 233824
rect 106917 233819 106983 233822
rect 152273 233819 152339 233822
rect 70301 233474 70367 233477
rect 229921 233474 229987 233477
rect 70301 233472 229987 233474
rect 70301 233416 70306 233472
rect 70362 233416 229926 233472
rect 229982 233416 229987 233472
rect 70301 233414 229987 233416
rect 70301 233411 70367 233414
rect 229921 233411 229987 233414
rect 67541 233338 67607 233341
rect 228214 233338 228220 233340
rect 67541 233336 228220 233338
rect 67541 233280 67546 233336
rect 67602 233280 228220 233336
rect 67541 233278 228220 233280
rect 67541 233275 67607 233278
rect 228214 233276 228220 233278
rect 228284 233276 228290 233340
rect 218973 233202 219039 233205
rect 227529 233202 227595 233205
rect 218973 233200 227595 233202
rect 218973 233144 218978 233200
rect 219034 233144 227534 233200
rect 227590 233144 227595 233200
rect 218973 233142 227595 233144
rect 218973 233139 219039 233142
rect 227529 233139 227595 233142
rect 215661 233066 215727 233069
rect 224902 233066 224908 233068
rect 215661 233064 224908 233066
rect 215661 233008 215666 233064
rect 215722 233008 224908 233064
rect 215661 233006 224908 233008
rect 215661 233003 215727 233006
rect 224902 233004 224908 233006
rect 224972 233004 224978 233068
rect 215293 232930 215359 232933
rect 224585 232930 224651 232933
rect 215293 232928 224651 232930
rect 215293 232872 215298 232928
rect 215354 232872 224590 232928
rect 224646 232872 224651 232928
rect 215293 232870 224651 232872
rect 215293 232867 215359 232870
rect 224585 232867 224651 232870
rect 215845 232794 215911 232797
rect 225321 232794 225387 232797
rect 215845 232792 225387 232794
rect 215845 232736 215850 232792
rect 215906 232736 225326 232792
rect 225382 232736 225387 232792
rect 215845 232734 225387 232736
rect 215845 232731 215911 232734
rect 225321 232731 225387 232734
rect 215753 232658 215819 232661
rect 227437 232658 227503 232661
rect 215753 232656 227503 232658
rect 215753 232600 215758 232656
rect 215814 232600 227442 232656
rect 227498 232600 227503 232656
rect 215753 232598 227503 232600
rect 215753 232595 215819 232598
rect 227437 232595 227503 232598
rect 59997 232522 60063 232525
rect 125041 232522 125107 232525
rect 59997 232520 125107 232522
rect 59997 232464 60002 232520
rect 60058 232464 125046 232520
rect 125102 232464 125107 232520
rect 59997 232462 125107 232464
rect 59997 232459 60063 232462
rect 125041 232459 125107 232462
rect 215477 232522 215543 232525
rect 226926 232522 226932 232524
rect 215477 232520 226932 232522
rect 215477 232464 215482 232520
rect 215538 232464 226932 232520
rect 215477 232462 226932 232464
rect 215477 232459 215543 232462
rect 226926 232460 226932 232462
rect 226996 232460 227002 232524
rect 15837 232386 15903 232389
rect 157977 232386 158043 232389
rect 583520 232386 584960 232476
rect 15837 232384 158043 232386
rect 15837 232328 15842 232384
rect 15898 232328 157982 232384
rect 158038 232328 158043 232384
rect 15837 232326 158043 232328
rect 15837 232323 15903 232326
rect 157977 232323 158043 232326
rect 583342 232326 584960 232386
rect 17217 232250 17283 232253
rect 160737 232250 160803 232253
rect 17217 232248 160803 232250
rect 17217 232192 17222 232248
rect 17278 232192 160742 232248
rect 160798 232192 160803 232248
rect 17217 232190 160803 232192
rect 583342 232250 583402 232326
rect 583520 232250 584960 232326
rect 583342 232236 584960 232250
rect 583342 232190 583586 232236
rect 17217 232187 17283 232190
rect 160737 232187 160803 232190
rect 64597 232114 64663 232117
rect 232589 232114 232655 232117
rect 64597 232112 232655 232114
rect 64597 232056 64602 232112
rect 64658 232056 232594 232112
rect 232650 232056 232655 232112
rect 64597 232054 232655 232056
rect 64597 232051 64663 232054
rect 232589 232051 232655 232054
rect 75729 231978 75795 231981
rect 583526 231978 583586 232190
rect 75729 231976 583586 231978
rect 75729 231920 75734 231976
rect 75790 231920 583586 231976
rect 75729 231918 583586 231920
rect 75729 231915 75795 231918
rect 108757 231162 108823 231165
rect 108941 231162 109007 231165
rect 108757 231160 109007 231162
rect 108757 231104 108762 231160
rect 108818 231104 108946 231160
rect 109002 231104 109007 231160
rect 108757 231102 109007 231104
rect 108757 231099 108823 231102
rect 108941 231099 109007 231102
rect 22737 231026 22803 231029
rect 165981 231026 166047 231029
rect 22737 231024 166047 231026
rect 22737 230968 22742 231024
rect 22798 230968 165986 231024
rect 166042 230968 166047 231024
rect 22737 230966 166047 230968
rect 22737 230963 22803 230966
rect 165981 230963 166047 230966
rect 14457 230890 14523 230893
rect 160277 230890 160343 230893
rect 14457 230888 160343 230890
rect 14457 230832 14462 230888
rect 14518 230832 160282 230888
rect 160338 230832 160343 230888
rect 14457 230830 160343 230832
rect 14457 230827 14523 230830
rect 160277 230827 160343 230830
rect 217317 230890 217383 230893
rect 220077 230890 220143 230893
rect 217317 230888 220143 230890
rect 217317 230832 217322 230888
rect 217378 230832 220082 230888
rect 220138 230832 220143 230888
rect 217317 230830 220143 230832
rect 217317 230827 217383 230830
rect 220077 230827 220143 230830
rect 72785 230754 72851 230757
rect 278037 230754 278103 230757
rect 72785 230752 278103 230754
rect 72785 230696 72790 230752
rect 72846 230696 278042 230752
rect 278098 230696 278103 230752
rect 72785 230694 278103 230696
rect 72785 230691 72851 230694
rect 278037 230691 278103 230694
rect 63309 230618 63375 230621
rect 287697 230618 287763 230621
rect 63309 230616 287763 230618
rect 63309 230560 63314 230616
rect 63370 230560 287702 230616
rect 287758 230560 287763 230616
rect 63309 230558 287763 230560
rect 63309 230555 63375 230558
rect 287697 230555 287763 230558
rect 219893 230482 219959 230485
rect 225505 230482 225571 230485
rect 219893 230480 225571 230482
rect 219893 230424 219898 230480
rect 219954 230424 225510 230480
rect 225566 230424 225571 230480
rect 219893 230422 225571 230424
rect 219893 230419 219959 230422
rect 225505 230419 225571 230422
rect 95969 230346 96035 230349
rect 96521 230346 96587 230349
rect 95969 230344 96587 230346
rect 95969 230288 95974 230344
rect 96030 230288 96526 230344
rect 96582 230288 96587 230344
rect 95969 230286 96587 230288
rect 95969 230283 96035 230286
rect 96521 230283 96587 230286
rect 99649 230346 99715 230349
rect 100661 230346 100727 230349
rect 99649 230344 100727 230346
rect 99649 230288 99654 230344
rect 99710 230288 100666 230344
rect 100722 230288 100727 230344
rect 99649 230286 100727 230288
rect 99649 230283 99715 230286
rect 100661 230283 100727 230286
rect 105353 230346 105419 230349
rect 106181 230346 106247 230349
rect 105353 230344 106247 230346
rect 105353 230288 105358 230344
rect 105414 230288 106186 230344
rect 106242 230288 106247 230344
rect 105353 230286 106247 230288
rect 105353 230283 105419 230286
rect 106181 230283 106247 230286
rect 126973 230346 127039 230349
rect 127525 230346 127591 230349
rect 126973 230344 127591 230346
rect 126973 230288 126978 230344
rect 127034 230288 127530 230344
rect 127586 230288 127591 230344
rect 126973 230286 127591 230288
rect 126973 230283 127039 230286
rect 127525 230283 127591 230286
rect 203425 230346 203491 230349
rect 204161 230346 204227 230349
rect 203425 230344 204227 230346
rect 203425 230288 203430 230344
rect 203486 230288 204166 230344
rect 204222 230288 204227 230344
rect 203425 230286 204227 230288
rect 203425 230283 203491 230286
rect 204161 230283 204227 230286
rect 212533 230346 212599 230349
rect 213085 230346 213151 230349
rect 212533 230344 213151 230346
rect 212533 230288 212538 230344
rect 212594 230288 213090 230344
rect 213146 230288 213151 230344
rect 212533 230286 213151 230288
rect 212533 230283 212599 230286
rect 213085 230283 213151 230286
rect 218646 230284 218652 230348
rect 218716 230346 218722 230348
rect 224902 230346 224908 230348
rect 218716 230286 224908 230346
rect 218716 230284 218722 230286
rect 224902 230284 224908 230286
rect 224972 230284 224978 230348
rect 218789 230210 218855 230213
rect 226241 230210 226307 230213
rect 218789 230208 226307 230210
rect 218789 230152 218794 230208
rect 218850 230152 226246 230208
rect 226302 230152 226307 230208
rect 218789 230150 226307 230152
rect 218789 230147 218855 230150
rect 226241 230147 226307 230150
rect 216121 230074 216187 230077
rect 224677 230074 224743 230077
rect 216121 230072 224743 230074
rect 216121 230016 216126 230072
rect 216182 230016 224682 230072
rect 224738 230016 224743 230072
rect 216121 230014 224743 230016
rect 216121 230011 216187 230014
rect 224677 230011 224743 230014
rect 216489 229938 216555 229941
rect 225597 229938 225663 229941
rect 216489 229936 225663 229938
rect 216489 229880 216494 229936
rect 216550 229880 225602 229936
rect 225658 229880 225663 229936
rect 216489 229878 225663 229880
rect 216489 229875 216555 229878
rect 225597 229875 225663 229878
rect 216305 229802 216371 229805
rect 225689 229802 225755 229805
rect 216305 229800 225755 229802
rect 216305 229744 216310 229800
rect 216366 229744 225694 229800
rect 225750 229744 225755 229800
rect 216305 229742 225755 229744
rect 216305 229739 216371 229742
rect 225689 229739 225755 229742
rect 21357 229666 21423 229669
rect 163129 229666 163195 229669
rect 21357 229664 163195 229666
rect 21357 229608 21362 229664
rect 21418 229608 163134 229664
rect 163190 229608 163195 229664
rect 21357 229606 163195 229608
rect 21357 229603 21423 229606
rect 163129 229603 163195 229606
rect 11697 229530 11763 229533
rect 157425 229530 157491 229533
rect 11697 229528 157491 229530
rect 11697 229472 11702 229528
rect 11758 229472 157430 229528
rect 157486 229472 157491 229528
rect 11697 229470 157491 229472
rect 11697 229467 11763 229470
rect 157425 229467 157491 229470
rect 7557 229394 7623 229397
rect 154573 229394 154639 229397
rect 7557 229392 154639 229394
rect 7557 229336 7562 229392
rect 7618 229336 154578 229392
rect 154634 229336 154639 229392
rect 7557 229334 154639 229336
rect 7557 229331 7623 229334
rect 154573 229331 154639 229334
rect 69013 229258 69079 229261
rect 271137 229258 271203 229261
rect 69013 229256 271203 229258
rect 69013 229200 69018 229256
rect 69074 229200 271142 229256
rect 271198 229200 271203 229256
rect 69013 229198 271203 229200
rect 69013 229195 69079 229198
rect 271137 229195 271203 229198
rect 66161 229122 66227 229125
rect 580257 229122 580323 229125
rect 66161 229120 580323 229122
rect 66161 229064 66166 229120
rect 66222 229064 580262 229120
rect 580318 229064 580323 229120
rect 66161 229062 580323 229064
rect 66161 229059 66227 229062
rect 580257 229059 580323 229062
rect 102225 228986 102291 228989
rect 103329 228986 103395 228989
rect 102225 228984 103395 228986
rect 102225 228928 102230 228984
rect 102286 228928 103334 228984
rect 103390 228928 103395 228984
rect 102225 228926 103395 228928
rect 102225 228923 102291 228926
rect 103329 228923 103395 228926
rect 107929 228986 107995 228989
rect 108849 228986 108915 228989
rect 107929 228984 108915 228986
rect 107929 228928 107934 228984
rect 107990 228928 108854 228984
rect 108910 228928 108915 228984
rect 107929 228926 108915 228928
rect 107929 228923 107995 228926
rect 108849 228923 108915 228926
rect 216397 228850 216463 228853
rect 220169 228850 220235 228853
rect 216397 228848 220235 228850
rect 216397 228792 216402 228848
rect 216458 228792 220174 228848
rect 220230 228792 220235 228848
rect 216397 228790 220235 228792
rect 216397 228787 216463 228790
rect 220169 228787 220235 228790
rect 184933 228714 184999 228717
rect 200757 228714 200823 228717
rect 184933 228712 200823 228714
rect 184933 228656 184938 228712
rect 184994 228656 200762 228712
rect 200818 228656 200823 228712
rect 184933 228654 200823 228656
rect 184933 228651 184999 228654
rect 200757 228651 200823 228654
rect 216213 228714 216279 228717
rect 222009 228714 222075 228717
rect 216213 228712 222075 228714
rect 216213 228656 216218 228712
rect 216274 228656 222014 228712
rect 222070 228656 222075 228712
rect 216213 228654 222075 228656
rect 216213 228651 216279 228654
rect 222009 228651 222075 228654
rect 18597 228578 18663 228581
rect 159265 228578 159331 228581
rect 18597 228576 159331 228578
rect 18597 228520 18602 228576
rect 18658 228520 159270 228576
rect 159326 228520 159331 228576
rect 18597 228518 159331 228520
rect 18597 228515 18663 228518
rect 159265 228515 159331 228518
rect 179229 228578 179295 228581
rect 197353 228578 197419 228581
rect 179229 228576 197419 228578
rect 179229 228520 179234 228576
rect 179290 228520 197358 228576
rect 197414 228520 197419 228576
rect 179229 228518 197419 228520
rect 179229 228515 179295 228518
rect 197353 228515 197419 228518
rect 58341 228442 58407 228445
rect 123201 228442 123267 228445
rect 58341 228440 123267 228442
rect 58341 228384 58346 228440
rect 58402 228384 123206 228440
rect 123262 228384 123267 228440
rect 58341 228382 123267 228384
rect 58341 228379 58407 228382
rect 123201 228379 123267 228382
rect 174537 228442 174603 228445
rect 196709 228442 196775 228445
rect 174537 228440 196775 228442
rect 174537 228384 174542 228440
rect 174598 228384 196714 228440
rect 196770 228384 196775 228440
rect 174537 228382 196775 228384
rect 174537 228379 174603 228382
rect 196709 228379 196775 228382
rect 40677 228306 40743 228309
rect 164049 228306 164115 228309
rect 40677 228304 164115 228306
rect 40677 228248 40682 228304
rect 40738 228248 164054 228304
rect 164110 228248 164115 228304
rect 40677 228246 164115 228248
rect 40677 228243 40743 228246
rect 164049 228243 164115 228246
rect 170673 228306 170739 228309
rect 206461 228306 206527 228309
rect 170673 228304 206527 228306
rect 170673 228248 170678 228304
rect 170734 228248 206466 228304
rect 206522 228248 206527 228304
rect 170673 228246 206527 228248
rect 170673 228243 170739 228246
rect 206461 228243 206527 228246
rect 217961 228306 218027 228309
rect 227621 228306 227687 228309
rect 217961 228304 227687 228306
rect 217961 228248 217966 228304
rect 218022 228248 227626 228304
rect 227682 228248 227687 228304
rect 217961 228246 227687 228248
rect 217961 228243 218027 228246
rect 227621 228243 227687 228246
rect 36537 228170 36603 228173
rect 164969 228170 165035 228173
rect 36537 228168 165035 228170
rect -960 227884 480 228124
rect 36537 228112 36542 228168
rect 36598 228112 164974 228168
rect 165030 228112 165035 228168
rect 36537 228110 165035 228112
rect 36537 228107 36603 228110
rect 164969 228107 165035 228110
rect 25497 228034 25563 228037
rect 162117 228034 162183 228037
rect 25497 228032 162183 228034
rect 25497 227976 25502 228032
rect 25558 227976 162122 228032
rect 162178 227976 162183 228032
rect 25497 227974 162183 227976
rect 25497 227971 25563 227974
rect 162117 227971 162183 227974
rect 156597 227898 156663 227901
rect 166901 227898 166967 227901
rect 156597 227896 166967 227898
rect 156597 227840 156602 227896
rect 156658 227840 166906 227896
rect 166962 227840 166967 227896
rect 156597 227838 166967 227840
rect 156597 227835 156663 227838
rect 166901 227835 166967 227838
rect 183093 227898 183159 227901
rect 184197 227898 184263 227901
rect 183093 227896 184263 227898
rect 183093 227840 183098 227896
rect 183154 227840 184202 227896
rect 184258 227840 184263 227896
rect 183093 227838 184263 227840
rect 183093 227835 183159 227838
rect 184197 227835 184263 227838
rect 191649 227898 191715 227901
rect 197445 227898 197511 227901
rect 191649 227896 197511 227898
rect 191649 227840 191654 227896
rect 191710 227840 197450 227896
rect 197506 227840 197511 227896
rect 191649 227838 197511 227840
rect 191649 227835 191715 227838
rect 197445 227835 197511 227838
rect 222837 227898 222903 227901
rect 226558 227898 226564 227900
rect 222837 227896 226564 227898
rect 222837 227840 222842 227896
rect 222898 227840 226564 227896
rect 222837 227838 226564 227840
rect 222837 227835 222903 227838
rect 226558 227836 226564 227838
rect 226628 227836 226634 227900
rect 68001 227762 68067 227765
rect 302877 227762 302943 227765
rect 68001 227760 302943 227762
rect 68001 227704 68006 227760
rect 68062 227704 302882 227760
rect 302938 227704 302943 227760
rect 68001 227702 302943 227704
rect 68001 227699 68067 227702
rect 302877 227699 302943 227702
rect 74993 227490 75059 227493
rect 75821 227490 75887 227493
rect 74993 227488 75887 227490
rect 74993 227432 74998 227488
rect 75054 227432 75826 227488
rect 75882 227432 75887 227488
rect 74993 227430 75887 227432
rect 74993 227427 75059 227430
rect 75821 227427 75887 227430
rect 84561 227490 84627 227493
rect 85481 227490 85547 227493
rect 84561 227488 85547 227490
rect 84561 227432 84566 227488
rect 84622 227432 85486 227488
rect 85542 227432 85547 227488
rect 84561 227430 85547 227432
rect 84561 227427 84627 227430
rect 85481 227427 85547 227430
rect 138013 227490 138079 227493
rect 138933 227490 138999 227493
rect 138013 227488 138999 227490
rect 138013 227432 138018 227488
rect 138074 227432 138938 227488
rect 138994 227432 138999 227488
rect 138013 227430 138999 227432
rect 138013 227427 138079 227430
rect 138933 227427 138999 227430
rect 144913 227490 144979 227493
rect 145741 227490 145807 227493
rect 144913 227488 145807 227490
rect 144913 227432 144918 227488
rect 144974 227432 145746 227488
rect 145802 227432 145807 227488
rect 144913 227430 145807 227432
rect 144913 227427 144979 227430
rect 145741 227427 145807 227430
rect 175825 227490 175891 227493
rect 176561 227490 176627 227493
rect 175825 227488 176627 227490
rect 175825 227432 175830 227488
rect 175886 227432 176566 227488
rect 176622 227432 176627 227488
rect 175825 227430 176627 227432
rect 175825 227427 175891 227430
rect 176561 227427 176627 227430
rect 215753 227490 215819 227493
rect 216581 227490 216647 227493
rect 215753 227488 216647 227490
rect 215753 227432 215758 227488
rect 215814 227432 216586 227488
rect 216642 227432 216647 227488
rect 215753 227430 216647 227432
rect 215753 227427 215819 227430
rect 216581 227427 216647 227430
rect 218881 227490 218947 227493
rect 226006 227490 226012 227492
rect 218881 227488 226012 227490
rect 218881 227432 218886 227488
rect 218942 227432 226012 227488
rect 218881 227430 226012 227432
rect 218881 227427 218947 227430
rect 226006 227428 226012 227430
rect 226076 227428 226082 227492
rect 218697 227354 218763 227357
rect 225873 227354 225939 227357
rect 218697 227352 225939 227354
rect 218697 227296 218702 227352
rect 218758 227296 225878 227352
rect 225934 227296 225939 227352
rect 218697 227294 225939 227296
rect 218697 227291 218763 227294
rect 225873 227291 225939 227294
rect 219249 227218 219315 227221
rect 227345 227218 227411 227221
rect 219249 227216 227411 227218
rect 219249 227160 219254 227216
rect 219310 227160 227350 227216
rect 227406 227160 227411 227216
rect 219249 227158 227411 227160
rect 219249 227155 219315 227158
rect 227345 227155 227411 227158
rect 219065 227082 219131 227085
rect 227253 227082 227319 227085
rect 219065 227080 227319 227082
rect 219065 227024 219070 227080
rect 219126 227024 227258 227080
rect 227314 227024 227319 227080
rect 219065 227022 227319 227024
rect 219065 227019 219131 227022
rect 227253 227019 227319 227022
rect 3417 226946 3483 226949
rect 156597 226946 156663 226949
rect 3417 226944 156663 226946
rect 3417 226888 3422 226944
rect 3478 226888 156602 226944
rect 156658 226888 156663 226944
rect 3417 226886 156663 226888
rect 3417 226883 3483 226886
rect 156597 226883 156663 226886
rect 216029 226946 216095 226949
rect 229553 226946 229619 226949
rect 216029 226944 229619 226946
rect 216029 226888 216034 226944
rect 216090 226888 229558 226944
rect 229614 226888 229619 226944
rect 216029 226886 229619 226888
rect 216029 226883 216095 226886
rect 229553 226883 229619 226886
rect 29637 226810 29703 226813
rect 156413 226810 156479 226813
rect 29637 226808 156479 226810
rect 29637 226752 29642 226808
rect 29698 226752 156418 226808
rect 156474 226752 156479 226808
rect 29637 226750 156479 226752
rect 29637 226747 29703 226750
rect 156413 226747 156479 226750
rect 219985 226810 220051 226813
rect 225781 226810 225847 226813
rect 219985 226808 225847 226810
rect 219985 226752 219990 226808
rect 220046 226752 225786 226808
rect 225842 226752 225847 226808
rect 219985 226750 225847 226752
rect 219985 226747 220051 226750
rect 225781 226747 225847 226750
rect 4797 226674 4863 226677
rect 155125 226674 155191 226677
rect 4797 226672 155191 226674
rect 4797 226616 4802 226672
rect 4858 226616 155130 226672
rect 155186 226616 155191 226672
rect 4797 226614 155191 226616
rect 4797 226611 4863 226614
rect 155125 226611 155191 226614
rect 172881 226674 172947 226677
rect 173801 226674 173867 226677
rect 172881 226672 173867 226674
rect 172881 226616 172886 226672
rect 172942 226616 173806 226672
rect 173862 226616 173867 226672
rect 172881 226614 173867 226616
rect 172881 226611 172947 226614
rect 173801 226611 173867 226614
rect 180885 226674 180951 226677
rect 181805 226674 181871 226677
rect 180885 226672 181871 226674
rect 180885 226616 180890 226672
rect 180946 226616 181810 226672
rect 181866 226616 181871 226672
rect 180885 226614 181871 226616
rect 180885 226611 180951 226614
rect 181805 226611 181871 226614
rect 224217 226674 224283 226677
rect 224861 226674 224927 226677
rect 224217 226672 224927 226674
rect 224217 226616 224222 226672
rect 224278 226616 224866 226672
rect 224922 226616 224927 226672
rect 224217 226614 224927 226616
rect 224217 226611 224283 226614
rect 224861 226611 224927 226614
rect 65425 226538 65491 226541
rect 295977 226538 296043 226541
rect 65425 226536 296043 226538
rect 65425 226480 65430 226536
rect 65486 226480 295982 226536
rect 296038 226480 296043 226536
rect 65425 226478 296043 226480
rect 65425 226475 65491 226478
rect 295977 226475 296043 226478
rect 55673 226402 55739 226405
rect 62113 226402 62179 226405
rect 55673 226400 62179 226402
rect 55673 226344 55678 226400
rect 55734 226344 62118 226400
rect 62174 226344 62179 226400
rect 55673 226342 62179 226344
rect 55673 226339 55739 226342
rect 62113 226339 62179 226342
rect 71129 226402 71195 226405
rect 410517 226402 410583 226405
rect 71129 226400 410583 226402
rect 71129 226344 71134 226400
rect 71190 226344 410522 226400
rect 410578 226344 410583 226400
rect 71129 226342 410583 226344
rect 71129 226339 71195 226342
rect 410517 226339 410583 226342
rect 55765 226130 55831 226133
rect 61101 226130 61167 226133
rect 55765 226128 61167 226130
rect 55765 226072 55770 226128
rect 55826 226072 61106 226128
rect 61162 226072 61167 226128
rect 55765 226070 61167 226072
rect 55765 226067 55831 226070
rect 61101 226067 61167 226070
rect 57881 225994 57947 225997
rect 61745 225994 61811 225997
rect 78857 225994 78923 225997
rect 57881 225992 61811 225994
rect 57881 225936 57886 225992
rect 57942 225936 61750 225992
rect 61806 225936 61811 225992
rect 57881 225934 61811 225936
rect 57881 225931 57947 225934
rect 61745 225931 61811 225934
rect 64830 225992 78923 225994
rect 64830 225936 78862 225992
rect 78918 225936 78923 225992
rect 64830 225934 78923 225936
rect 58341 225586 58407 225589
rect 64830 225586 64890 225934
rect 78857 225931 78923 225934
rect 223665 225994 223731 225997
rect 223665 225992 223866 225994
rect 223665 225936 223670 225992
rect 223726 225936 223866 225992
rect 223665 225934 223866 225936
rect 223665 225931 223731 225934
rect 58341 225584 64890 225586
rect 58341 225528 58346 225584
rect 58402 225528 64890 225584
rect 58341 225526 64890 225528
rect 58341 225523 58407 225526
rect 56409 225314 56475 225317
rect 56409 225312 60076 225314
rect 56409 225256 56414 225312
rect 56470 225256 60076 225312
rect 223806 225284 223866 225934
rect 56409 225254 60076 225256
rect 56409 225251 56475 225254
rect 224769 225042 224835 225045
rect 227161 225042 227227 225045
rect 224769 225040 227227 225042
rect 224769 224984 224774 225040
rect 224830 224984 227166 225040
rect 227222 224984 227227 225040
rect 224769 224982 227227 224984
rect 224769 224979 224835 224982
rect 227161 224979 227227 224982
rect 56317 222594 56383 222597
rect 225413 222594 225479 222597
rect 56317 222592 60076 222594
rect 56317 222536 56322 222592
rect 56378 222536 60076 222592
rect 56317 222534 60076 222536
rect 224388 222592 225479 222594
rect 224388 222536 225418 222592
rect 225474 222536 225479 222592
rect 224388 222534 225479 222536
rect 56317 222531 56383 222534
rect 225413 222531 225479 222534
rect 227161 220962 227227 220965
rect 227294 220962 227300 220964
rect 227161 220960 227300 220962
rect 227161 220904 227166 220960
rect 227222 220904 227300 220960
rect 227161 220902 227300 220904
rect 227161 220899 227227 220902
rect 227294 220900 227300 220902
rect 227364 220900 227370 220964
rect 227161 220826 227227 220829
rect 282177 220826 282243 220829
rect 227161 220824 282243 220826
rect 227161 220768 227166 220824
rect 227222 220768 282182 220824
rect 282238 220768 282243 220824
rect 227161 220766 282243 220768
rect 227161 220763 227227 220766
rect 282177 220763 282243 220766
rect 57881 219874 57947 219877
rect 227161 219874 227227 219877
rect 57881 219872 60076 219874
rect 57881 219816 57886 219872
rect 57942 219816 60076 219872
rect 57881 219814 60076 219816
rect 224388 219872 227227 219874
rect 224388 219816 227166 219872
rect 227222 219816 227227 219872
rect 224388 219814 227227 219816
rect 57881 219811 57947 219814
rect 227161 219811 227227 219814
rect 227161 219738 227227 219741
rect 227621 219738 227687 219741
rect 227161 219736 227687 219738
rect 227161 219680 227166 219736
rect 227222 219680 227626 219736
rect 227682 219680 227687 219736
rect 227161 219678 227687 219680
rect 227161 219675 227227 219678
rect 227621 219675 227687 219678
rect 227294 219540 227300 219604
rect 227364 219602 227370 219604
rect 227621 219602 227687 219605
rect 227364 219600 227687 219602
rect 227364 219544 227626 219600
rect 227682 219544 227687 219600
rect 227364 219542 227687 219544
rect 227364 219540 227370 219542
rect 227621 219539 227687 219542
rect 583520 219058 584960 219148
rect 583342 218998 584960 219058
rect 583342 218922 583402 218998
rect 583520 218922 584960 218998
rect 583342 218908 584960 218922
rect 583342 218862 583586 218908
rect 228398 218044 228404 218108
rect 228468 218106 228474 218108
rect 583526 218106 583586 218862
rect 228468 218046 583586 218106
rect 228468 218044 228474 218046
rect 57513 217154 57579 217157
rect 227529 217154 227595 217157
rect 57513 217152 60076 217154
rect 57513 217096 57518 217152
rect 57574 217096 60076 217152
rect 57513 217094 60076 217096
rect 224388 217152 227595 217154
rect 224388 217096 227534 217152
rect 227590 217096 227595 217152
rect 224388 217094 227595 217096
rect 57513 217091 57579 217094
rect 227529 217091 227595 217094
rect -960 214978 480 215068
rect 3509 214978 3575 214981
rect -960 214976 3575 214978
rect -960 214920 3514 214976
rect 3570 214920 3575 214976
rect -960 214918 3575 214920
rect -960 214828 480 214918
rect 3509 214915 3575 214918
rect 59629 214570 59695 214573
rect 227621 214570 227687 214573
rect 59629 214568 60076 214570
rect 59629 214512 59634 214568
rect 59690 214512 60076 214568
rect 59629 214510 60076 214512
rect 224388 214568 227687 214570
rect 224388 214512 227626 214568
rect 227682 214512 227687 214568
rect 224388 214510 227687 214512
rect 59629 214507 59695 214510
rect 227621 214507 227687 214510
rect 227529 212530 227595 212533
rect 232681 212530 232747 212533
rect 227529 212528 232747 212530
rect 227529 212472 227534 212528
rect 227590 212472 232686 212528
rect 232742 212472 232747 212528
rect 227529 212470 232747 212472
rect 227529 212467 227595 212470
rect 232681 212467 232747 212470
rect 57605 211850 57671 211853
rect 227529 211850 227595 211853
rect 57605 211848 60076 211850
rect 57605 211792 57610 211848
rect 57666 211792 60076 211848
rect 57605 211790 60076 211792
rect 224388 211848 227595 211850
rect 224388 211792 227534 211848
rect 227590 211792 227595 211848
rect 224388 211790 227595 211792
rect 57605 211787 57671 211790
rect 227529 211787 227595 211790
rect 58433 209130 58499 209133
rect 228633 209130 228699 209133
rect 58433 209128 60076 209130
rect 58433 209072 58438 209128
rect 58494 209072 60076 209128
rect 58433 209070 60076 209072
rect 224388 209128 228699 209130
rect 224388 209072 228638 209128
rect 228694 209072 228699 209128
rect 224388 209070 228699 209072
rect 58433 209067 58499 209070
rect 228633 209067 228699 209070
rect 58525 206410 58591 206413
rect 228909 206410 228975 206413
rect 58525 206408 60076 206410
rect 58525 206352 58530 206408
rect 58586 206352 60076 206408
rect 58525 206350 60076 206352
rect 224388 206408 228975 206410
rect 224388 206352 228914 206408
rect 228970 206352 228975 206408
rect 224388 206350 228975 206352
rect 58525 206347 58591 206350
rect 228909 206347 228975 206350
rect 580165 205730 580231 205733
rect 583520 205730 584960 205820
rect 580165 205728 584960 205730
rect 580165 205672 580170 205728
rect 580226 205672 584960 205728
rect 580165 205670 584960 205672
rect 580165 205667 580231 205670
rect 583520 205580 584960 205670
rect 56501 203826 56567 203829
rect 235349 203826 235415 203829
rect 56501 203824 60076 203826
rect 56501 203768 56506 203824
rect 56562 203768 60076 203824
rect 56501 203766 60076 203768
rect 224388 203824 235415 203826
rect 224388 203768 235354 203824
rect 235410 203768 235415 203824
rect 224388 203766 235415 203768
rect 56501 203763 56567 203766
rect 235349 203763 235415 203766
rect -960 201922 480 202012
rect 3049 201922 3115 201925
rect -960 201920 3115 201922
rect -960 201864 3054 201920
rect 3110 201864 3115 201920
rect -960 201862 3115 201864
rect -960 201772 480 201862
rect 3049 201859 3115 201862
rect 307017 201378 307083 201381
rect 229050 201376 307083 201378
rect 229050 201320 307022 201376
rect 307078 201320 307083 201376
rect 229050 201318 307083 201320
rect 58709 201106 58775 201109
rect 229050 201106 229110 201318
rect 307017 201315 307083 201318
rect 58709 201104 60076 201106
rect 58709 201048 58714 201104
rect 58770 201048 60076 201104
rect 58709 201046 60076 201048
rect 224388 201046 229110 201106
rect 58709 201043 58775 201046
rect 57605 198386 57671 198389
rect 227437 198386 227503 198389
rect 57605 198384 60076 198386
rect 57605 198328 57610 198384
rect 57666 198328 60076 198384
rect 57605 198326 60076 198328
rect 224388 198384 227503 198386
rect 224388 198328 227442 198384
rect 227498 198328 227503 198384
rect 224388 198326 227503 198328
rect 57605 198323 57671 198326
rect 227437 198323 227503 198326
rect 57605 195666 57671 195669
rect 226149 195666 226215 195669
rect 57605 195664 60076 195666
rect 57605 195608 57610 195664
rect 57666 195608 60076 195664
rect 57605 195606 60076 195608
rect 224388 195664 226215 195666
rect 224388 195608 226154 195664
rect 226210 195608 226215 195664
rect 224388 195606 226215 195608
rect 57605 195603 57671 195606
rect 226149 195603 226215 195606
rect 233877 193898 233943 193901
rect 267825 193898 267891 193901
rect 233877 193896 267891 193898
rect 233877 193840 233882 193896
rect 233938 193840 267830 193896
rect 267886 193840 267891 193896
rect 233877 193838 267891 193840
rect 233877 193835 233943 193838
rect 267825 193835 267891 193838
rect 55857 192946 55923 192949
rect 233877 192946 233943 192949
rect 55857 192944 60076 192946
rect 55857 192888 55862 192944
rect 55918 192888 60076 192944
rect 55857 192886 60076 192888
rect 224388 192944 233943 192946
rect 224388 192888 233882 192944
rect 233938 192888 233943 192944
rect 224388 192886 233943 192888
rect 55857 192883 55923 192886
rect 233877 192883 233943 192886
rect 580165 192538 580231 192541
rect 583520 192538 584960 192628
rect 580165 192536 584960 192538
rect 580165 192480 580170 192536
rect 580226 192480 584960 192536
rect 580165 192478 584960 192480
rect 580165 192475 580231 192478
rect 583520 192388 584960 192478
rect 57605 190362 57671 190365
rect 230749 190362 230815 190365
rect 57605 190360 60076 190362
rect 57605 190304 57610 190360
rect 57666 190304 60076 190360
rect 57605 190302 60076 190304
rect 224388 190360 230815 190362
rect 224388 190304 230754 190360
rect 230810 190304 230815 190360
rect 224388 190302 230815 190304
rect 57605 190299 57671 190302
rect 230749 190299 230815 190302
rect -960 188866 480 188956
rect 2773 188866 2839 188869
rect -960 188864 2839 188866
rect -960 188808 2778 188864
rect 2834 188808 2839 188864
rect -960 188806 2839 188808
rect -960 188716 480 188806
rect 2773 188803 2839 188806
rect 58801 187642 58867 187645
rect 300117 187642 300183 187645
rect 58801 187640 60076 187642
rect 58801 187584 58806 187640
rect 58862 187584 60076 187640
rect 58801 187582 60076 187584
rect 224388 187640 300183 187642
rect 224388 187584 300122 187640
rect 300178 187584 300183 187640
rect 224388 187582 300183 187584
rect 58801 187579 58867 187582
rect 300117 187579 300183 187582
rect 57605 184922 57671 184925
rect 228449 184922 228515 184925
rect 57605 184920 60076 184922
rect 57605 184864 57610 184920
rect 57666 184864 60076 184920
rect 57605 184862 60076 184864
rect 224388 184920 228515 184922
rect 224388 184864 228454 184920
rect 228510 184864 228515 184920
rect 224388 184862 228515 184864
rect 57605 184859 57671 184862
rect 228449 184859 228515 184862
rect 57605 182202 57671 182205
rect 226701 182202 226767 182205
rect 57605 182200 60076 182202
rect 57605 182144 57610 182200
rect 57666 182144 60076 182200
rect 57605 182142 60076 182144
rect 224388 182200 226767 182202
rect 224388 182144 226706 182200
rect 226762 182144 226767 182200
rect 224388 182142 226767 182144
rect 57605 182139 57671 182142
rect 226701 182139 226767 182142
rect 56869 179618 56935 179621
rect 228357 179618 228423 179621
rect 56869 179616 60076 179618
rect 56869 179560 56874 179616
rect 56930 179560 60076 179616
rect 56869 179558 60076 179560
rect 224388 179616 228423 179618
rect 224388 179560 228362 179616
rect 228418 179560 228423 179616
rect 224388 179558 228423 179560
rect 56869 179555 56935 179558
rect 228357 179555 228423 179558
rect 583520 179210 584960 179300
rect 583342 179150 584960 179210
rect 583342 179074 583402 179150
rect 583520 179074 584960 179150
rect 583342 179060 584960 179074
rect 583342 179014 583586 179060
rect 231209 178122 231275 178125
rect 583526 178122 583586 179014
rect 231209 178120 583586 178122
rect 231209 178064 231214 178120
rect 231270 178064 583586 178120
rect 231209 178062 583586 178064
rect 231209 178059 231275 178062
rect 55949 176898 56015 176901
rect 229001 176898 229067 176901
rect 55949 176896 60076 176898
rect 55949 176840 55954 176896
rect 56010 176840 60076 176896
rect 55949 176838 60076 176840
rect 224388 176896 229067 176898
rect 224388 176840 229006 176896
rect 229062 176840 229067 176896
rect 224388 176838 229067 176840
rect 55949 176835 56015 176838
rect 229001 176835 229067 176838
rect -960 175796 480 176036
rect 226701 175266 226767 175269
rect 262213 175266 262279 175269
rect 226701 175264 262279 175266
rect 226701 175208 226706 175264
rect 226762 175208 262218 175264
rect 262274 175208 262279 175264
rect 226701 175206 262279 175208
rect 226701 175203 226767 175206
rect 262213 175203 262279 175206
rect 58157 174178 58223 174181
rect 226701 174178 226767 174181
rect 58157 174176 60076 174178
rect 58157 174120 58162 174176
rect 58218 174120 60076 174176
rect 58157 174118 60076 174120
rect 224388 174176 226767 174178
rect 224388 174120 226706 174176
rect 226762 174120 226767 174176
rect 224388 174118 226767 174120
rect 58157 174115 58223 174118
rect 226701 174115 226767 174118
rect 57605 171458 57671 171461
rect 228265 171458 228331 171461
rect 57605 171456 60076 171458
rect 57605 171400 57610 171456
rect 57666 171400 60076 171456
rect 57605 171398 60076 171400
rect 224388 171456 228331 171458
rect 224388 171400 228270 171456
rect 228326 171400 228331 171456
rect 224388 171398 228331 171400
rect 57605 171395 57671 171398
rect 228265 171395 228331 171398
rect 226701 169690 226767 169693
rect 246297 169690 246363 169693
rect 226701 169688 246363 169690
rect 226701 169632 226706 169688
rect 226762 169632 246302 169688
rect 246358 169632 246363 169688
rect 226701 169630 246363 169632
rect 226701 169627 226767 169630
rect 246297 169627 246363 169630
rect 57605 168738 57671 168741
rect 226701 168738 226767 168741
rect 57605 168736 60076 168738
rect 57605 168680 57610 168736
rect 57666 168680 60076 168736
rect 57605 168678 60076 168680
rect 224388 168736 226767 168738
rect 224388 168680 226706 168736
rect 226762 168680 226767 168736
rect 224388 168678 226767 168680
rect 57605 168675 57671 168678
rect 226701 168675 226767 168678
rect 57605 166154 57671 166157
rect 227345 166154 227411 166157
rect 57605 166152 60076 166154
rect 57605 166096 57610 166152
rect 57666 166096 60076 166152
rect 57605 166094 60076 166096
rect 224388 166152 227411 166154
rect 224388 166096 227350 166152
rect 227406 166096 227411 166152
rect 224388 166094 227411 166096
rect 57605 166091 57671 166094
rect 227345 166091 227411 166094
rect 580165 165882 580231 165885
rect 583520 165882 584960 165972
rect 580165 165880 584960 165882
rect 580165 165824 580170 165880
rect 580226 165824 584960 165880
rect 580165 165822 584960 165824
rect 580165 165819 580231 165822
rect 583520 165732 584960 165822
rect 57605 163434 57671 163437
rect 228081 163434 228147 163437
rect 57605 163432 60076 163434
rect 57605 163376 57610 163432
rect 57666 163376 60076 163432
rect 57605 163374 60076 163376
rect 224388 163432 228147 163434
rect 224388 163376 228086 163432
rect 228142 163376 228147 163432
rect 224388 163374 228147 163376
rect 57605 163371 57671 163374
rect 228081 163371 228147 163374
rect -960 162890 480 162980
rect 3233 162890 3299 162893
rect -960 162888 3299 162890
rect -960 162832 3238 162888
rect 3294 162832 3299 162888
rect -960 162830 3299 162832
rect -960 162740 480 162830
rect 3233 162827 3299 162830
rect 57237 160714 57303 160717
rect 228173 160714 228239 160717
rect 57237 160712 60076 160714
rect 57237 160656 57242 160712
rect 57298 160656 60076 160712
rect 57237 160654 60076 160656
rect 224388 160712 228239 160714
rect 224388 160656 228178 160712
rect 228234 160656 228239 160712
rect 224388 160654 228239 160656
rect 57237 160651 57303 160654
rect 228173 160651 228239 160654
rect 57605 157994 57671 157997
rect 226609 157994 226675 157997
rect 57605 157992 60076 157994
rect 57605 157936 57610 157992
rect 57666 157936 60076 157992
rect 57605 157934 60076 157936
rect 224388 157992 226675 157994
rect 224388 157936 226614 157992
rect 226670 157936 226675 157992
rect 224388 157934 226675 157936
rect 57605 157931 57671 157934
rect 226609 157931 226675 157934
rect 240869 155954 240935 155957
rect 229050 155952 240935 155954
rect 229050 155896 240874 155952
rect 240930 155896 240935 155952
rect 229050 155894 240935 155896
rect 58893 155410 58959 155413
rect 229050 155410 229110 155894
rect 240869 155891 240935 155894
rect 58893 155408 60076 155410
rect 58893 155352 58898 155408
rect 58954 155352 60076 155408
rect 58893 155350 60076 155352
rect 224388 155350 229110 155410
rect 58893 155347 58959 155350
rect 57605 152690 57671 152693
rect 230657 152690 230723 152693
rect 583520 152690 584960 152780
rect 57605 152688 60076 152690
rect 57605 152632 57610 152688
rect 57666 152632 60076 152688
rect 57605 152630 60076 152632
rect 224388 152688 230723 152690
rect 224388 152632 230662 152688
rect 230718 152632 230723 152688
rect 224388 152630 230723 152632
rect 57605 152627 57671 152630
rect 230657 152627 230723 152630
rect 583342 152630 584960 152690
rect 583342 152554 583402 152630
rect 583520 152554 584960 152630
rect 583342 152540 584960 152554
rect 583342 152494 583586 152540
rect 229921 151874 229987 151877
rect 583526 151874 583586 152494
rect 229921 151872 583586 151874
rect 229921 151816 229926 151872
rect 229982 151816 583586 151872
rect 229921 151814 583586 151816
rect 229921 151811 229987 151814
rect 57605 149970 57671 149973
rect 226517 149970 226583 149973
rect 57605 149968 60076 149970
rect -960 149834 480 149924
rect 57605 149912 57610 149968
rect 57666 149912 60076 149968
rect 57605 149910 60076 149912
rect 224388 149968 226583 149970
rect 224388 149912 226522 149968
rect 226578 149912 226583 149968
rect 224388 149910 226583 149912
rect 57605 149907 57671 149910
rect 226517 149907 226583 149910
rect 3509 149834 3575 149837
rect -960 149832 3575 149834
rect -960 149776 3514 149832
rect 3570 149776 3575 149832
rect -960 149774 3575 149776
rect -960 149684 480 149774
rect 3509 149771 3575 149774
rect 244917 147658 244983 147661
rect 229050 147656 244983 147658
rect 229050 147600 244922 147656
rect 244978 147600 244983 147656
rect 229050 147598 244983 147600
rect 58985 147250 59051 147253
rect 229050 147250 229110 147598
rect 244917 147595 244983 147598
rect 58985 147248 60076 147250
rect 58985 147192 58990 147248
rect 59046 147192 60076 147248
rect 58985 147190 60076 147192
rect 224388 147190 229110 147250
rect 58985 147187 59051 147190
rect 57605 144666 57671 144669
rect 227253 144666 227319 144669
rect 57605 144664 60076 144666
rect 57605 144608 57610 144664
rect 57666 144608 60076 144664
rect 57605 144606 60076 144608
rect 224388 144664 227319 144666
rect 224388 144608 227258 144664
rect 227314 144608 227319 144664
rect 224388 144606 227319 144608
rect 57605 144603 57671 144606
rect 227253 144603 227319 144606
rect 57605 141946 57671 141949
rect 226057 141946 226123 141949
rect 57605 141944 60076 141946
rect 57605 141888 57610 141944
rect 57666 141888 60076 141944
rect 57605 141886 60076 141888
rect 224388 141944 226123 141946
rect 224388 141888 226062 141944
rect 226118 141888 226123 141944
rect 224388 141886 226123 141888
rect 57605 141883 57671 141886
rect 226057 141883 226123 141886
rect 580165 139362 580231 139365
rect 583520 139362 584960 139452
rect 580165 139360 584960 139362
rect 580165 139304 580170 139360
rect 580226 139304 584960 139360
rect 580165 139302 584960 139304
rect 580165 139299 580231 139302
rect 56041 139226 56107 139229
rect 226425 139226 226491 139229
rect 56041 139224 60076 139226
rect 56041 139168 56046 139224
rect 56102 139168 60076 139224
rect 56041 139166 60076 139168
rect 224388 139224 226491 139226
rect 224388 139168 226430 139224
rect 226486 139168 226491 139224
rect 583520 139212 584960 139302
rect 224388 139166 226491 139168
rect 56041 139163 56107 139166
rect 226425 139163 226491 139166
rect -960 136778 480 136868
rect 3509 136778 3575 136781
rect -960 136776 3575 136778
rect -960 136720 3514 136776
rect 3570 136720 3575 136776
rect -960 136718 3575 136720
rect -960 136628 480 136718
rect 3509 136715 3575 136718
rect 253197 136642 253263 136645
rect 229050 136640 253263 136642
rect 229050 136584 253202 136640
rect 253258 136584 253263 136640
rect 229050 136582 253263 136584
rect 57605 136506 57671 136509
rect 229050 136506 229110 136582
rect 253197 136579 253263 136582
rect 57605 136504 60076 136506
rect 57605 136448 57610 136504
rect 57666 136448 60076 136504
rect 57605 136446 60076 136448
rect 224388 136446 229110 136506
rect 57605 136443 57671 136446
rect 57605 133786 57671 133789
rect 238109 133786 238175 133789
rect 57605 133784 60076 133786
rect 57605 133728 57610 133784
rect 57666 133728 60076 133784
rect 57605 133726 60076 133728
rect 224388 133784 238175 133786
rect 224388 133728 238114 133784
rect 238170 133728 238175 133784
rect 224388 133726 238175 133728
rect 57605 133723 57671 133726
rect 238109 133723 238175 133726
rect 57605 131202 57671 131205
rect 225965 131202 226031 131205
rect 57605 131200 60076 131202
rect 57605 131144 57610 131200
rect 57666 131144 60076 131200
rect 57605 131142 60076 131144
rect 224388 131200 226031 131202
rect 224388 131144 225970 131200
rect 226026 131144 226031 131200
rect 224388 131142 226031 131144
rect 57605 131139 57671 131142
rect 225965 131139 226031 131142
rect 59077 128482 59143 128485
rect 227069 128482 227135 128485
rect 59077 128480 60076 128482
rect 59077 128424 59082 128480
rect 59138 128424 60076 128480
rect 59077 128422 60076 128424
rect 224388 128480 227135 128482
rect 224388 128424 227074 128480
rect 227130 128424 227135 128480
rect 224388 128422 227135 128424
rect 59077 128419 59143 128422
rect 227069 128419 227135 128422
rect 226425 126986 226491 126989
rect 232497 126986 232563 126989
rect 226425 126984 232563 126986
rect 226425 126928 226430 126984
rect 226486 126928 232502 126984
rect 232558 126928 232563 126984
rect 226425 126926 232563 126928
rect 226425 126923 226491 126926
rect 232497 126923 232563 126926
rect 580165 126034 580231 126037
rect 583520 126034 584960 126124
rect 580165 126032 584960 126034
rect 580165 125976 580170 126032
rect 580226 125976 584960 126032
rect 580165 125974 584960 125976
rect 580165 125971 580231 125974
rect 583520 125884 584960 125974
rect 59537 125762 59603 125765
rect 226425 125762 226491 125765
rect 59537 125760 60076 125762
rect 59537 125704 59542 125760
rect 59598 125704 60076 125760
rect 59537 125702 60076 125704
rect 224388 125760 226491 125762
rect 224388 125704 226430 125760
rect 226486 125704 226491 125760
rect 224388 125702 226491 125704
rect 59537 125699 59603 125702
rect 226425 125699 226491 125702
rect -960 123572 480 123812
rect 57789 123042 57855 123045
rect 227161 123042 227227 123045
rect 57789 123040 60076 123042
rect 57789 122984 57794 123040
rect 57850 122984 60076 123040
rect 57789 122982 60076 122984
rect 224388 123040 227227 123042
rect 224388 122984 227166 123040
rect 227222 122984 227227 123040
rect 224388 122982 227227 122984
rect 57789 122979 57855 122982
rect 227161 122979 227227 122982
rect 57697 120458 57763 120461
rect 232313 120458 232379 120461
rect 57697 120456 60076 120458
rect 57697 120400 57702 120456
rect 57758 120400 60076 120456
rect 57697 120398 60076 120400
rect 224388 120456 232379 120458
rect 224388 120400 232318 120456
rect 232374 120400 232379 120456
rect 224388 120398 232379 120400
rect 57697 120395 57763 120398
rect 232313 120395 232379 120398
rect 57605 117738 57671 117741
rect 229829 117738 229895 117741
rect 57605 117736 60076 117738
rect 57605 117680 57610 117736
rect 57666 117680 60076 117736
rect 57605 117678 60076 117680
rect 224388 117736 229895 117738
rect 224388 117680 229834 117736
rect 229890 117680 229895 117736
rect 224388 117678 229895 117680
rect 57605 117675 57671 117678
rect 229829 117675 229895 117678
rect 57605 115018 57671 115021
rect 226742 115018 226748 115020
rect 57605 115016 60076 115018
rect 57605 114960 57610 115016
rect 57666 114960 60076 115016
rect 57605 114958 60076 114960
rect 224388 114958 226748 115018
rect 57605 114955 57671 114958
rect 226742 114956 226748 114958
rect 226812 114956 226818 115020
rect 583520 112842 584960 112932
rect 583342 112782 584960 112842
rect 583342 112706 583402 112782
rect 583520 112706 584960 112782
rect 583342 112692 584960 112706
rect 583342 112646 583586 112692
rect 58249 112298 58315 112301
rect 231117 112298 231183 112301
rect 58249 112296 60076 112298
rect 58249 112240 58254 112296
rect 58310 112240 60076 112296
rect 58249 112238 60076 112240
rect 224388 112296 231183 112298
rect 224388 112240 231122 112296
rect 231178 112240 231183 112296
rect 224388 112238 231183 112240
rect 58249 112235 58315 112238
rect 231117 112235 231183 112238
rect 228214 111828 228220 111892
rect 228284 111890 228290 111892
rect 583526 111890 583586 112646
rect 228284 111830 583586 111890
rect 228284 111828 228290 111830
rect -960 110666 480 110756
rect 3141 110666 3207 110669
rect -960 110664 3207 110666
rect -960 110608 3146 110664
rect 3202 110608 3207 110664
rect -960 110606 3207 110608
rect -960 110516 480 110606
rect 3141 110603 3207 110606
rect 57605 109578 57671 109581
rect 226333 109578 226399 109581
rect 57605 109576 60076 109578
rect 57605 109520 57610 109576
rect 57666 109520 60076 109576
rect 57605 109518 60076 109520
rect 224388 109576 226399 109578
rect 224388 109520 226338 109576
rect 226394 109520 226399 109576
rect 224388 109518 226399 109520
rect 57605 109515 57671 109518
rect 226333 109515 226399 109518
rect 57605 106994 57671 106997
rect 226926 106994 226932 106996
rect 57605 106992 60076 106994
rect 57605 106936 57610 106992
rect 57666 106936 60076 106992
rect 57605 106934 60076 106936
rect 224388 106934 226932 106994
rect 57605 106931 57671 106934
rect 226926 106932 226932 106934
rect 226996 106932 227002 106996
rect 57605 104274 57671 104277
rect 229645 104274 229711 104277
rect 57605 104272 60076 104274
rect 57605 104216 57610 104272
rect 57666 104216 60076 104272
rect 57605 104214 60076 104216
rect 224388 104272 229711 104274
rect 224388 104216 229650 104272
rect 229706 104216 229711 104272
rect 224388 104214 229711 104216
rect 57605 104211 57671 104214
rect 229645 104211 229711 104214
rect 57605 101554 57671 101557
rect 232221 101554 232287 101557
rect 57605 101552 60076 101554
rect 57605 101496 57610 101552
rect 57666 101496 60076 101552
rect 57605 101494 60076 101496
rect 224388 101552 232287 101554
rect 224388 101496 232226 101552
rect 232282 101496 232287 101552
rect 224388 101494 232287 101496
rect 57605 101491 57671 101494
rect 232221 101491 232287 101494
rect 580165 99514 580231 99517
rect 583520 99514 584960 99604
rect 580165 99512 584960 99514
rect 580165 99456 580170 99512
rect 580226 99456 584960 99512
rect 580165 99454 584960 99456
rect 580165 99451 580231 99454
rect 583520 99364 584960 99454
rect 58525 98834 58591 98837
rect 229737 98834 229803 98837
rect 58525 98832 60076 98834
rect 58525 98776 58530 98832
rect 58586 98776 60076 98832
rect 58525 98774 60076 98776
rect 224388 98832 229803 98834
rect 224388 98776 229742 98832
rect 229798 98776 229803 98832
rect 224388 98774 229803 98776
rect 58525 98771 58591 98774
rect 229737 98771 229803 98774
rect -960 97610 480 97700
rect 3509 97610 3575 97613
rect -960 97608 3575 97610
rect -960 97552 3514 97608
rect 3570 97552 3575 97608
rect -960 97550 3575 97552
rect -960 97460 480 97550
rect 3509 97547 3575 97550
rect 57145 96250 57211 96253
rect 232037 96250 232103 96253
rect 57145 96248 60076 96250
rect 57145 96192 57150 96248
rect 57206 96192 60076 96248
rect 57145 96190 60076 96192
rect 224388 96248 232103 96250
rect 224388 96192 232042 96248
rect 232098 96192 232103 96248
rect 224388 96190 232103 96192
rect 57145 96187 57211 96190
rect 232037 96187 232103 96190
rect 59261 93530 59327 93533
rect 232129 93530 232195 93533
rect 59261 93528 60076 93530
rect 59261 93472 59266 93528
rect 59322 93472 60076 93528
rect 59261 93470 60076 93472
rect 224388 93528 232195 93530
rect 224388 93472 232134 93528
rect 232190 93472 232195 93528
rect 224388 93470 232195 93472
rect 59261 93467 59327 93470
rect 232129 93467 232195 93470
rect 228081 91762 228147 91765
rect 255313 91762 255379 91765
rect 228081 91760 255379 91762
rect 228081 91704 228086 91760
rect 228142 91704 255318 91760
rect 255374 91704 255379 91760
rect 228081 91702 255379 91704
rect 228081 91699 228147 91702
rect 255313 91699 255379 91702
rect 57605 90810 57671 90813
rect 228081 90810 228147 90813
rect 57605 90808 60076 90810
rect 57605 90752 57610 90808
rect 57666 90752 60076 90808
rect 57605 90750 60076 90752
rect 224388 90808 228147 90810
rect 224388 90752 228086 90808
rect 228142 90752 228147 90808
rect 224388 90750 228147 90752
rect 57605 90747 57671 90750
rect 228081 90747 228147 90750
rect 57605 88090 57671 88093
rect 226885 88090 226951 88093
rect 57605 88088 60076 88090
rect 57605 88032 57610 88088
rect 57666 88032 60076 88088
rect 57605 88030 60076 88032
rect 224388 88088 226951 88090
rect 224388 88032 226890 88088
rect 226946 88032 226951 88088
rect 224388 88030 226951 88032
rect 57605 88027 57671 88030
rect 226885 88027 226951 88030
rect 580257 86186 580323 86189
rect 583520 86186 584960 86276
rect 580257 86184 584960 86186
rect 580257 86128 580262 86184
rect 580318 86128 584960 86184
rect 580257 86126 584960 86128
rect 580257 86123 580323 86126
rect 583520 86036 584960 86126
rect 57605 85370 57671 85373
rect 226374 85370 226380 85372
rect 57605 85368 60076 85370
rect 57605 85312 57610 85368
rect 57666 85312 60076 85368
rect 57605 85310 60076 85312
rect 224388 85310 226380 85370
rect 57605 85307 57671 85310
rect 226374 85308 226380 85310
rect 226444 85308 226450 85372
rect -960 84690 480 84780
rect 3509 84690 3575 84693
rect -960 84688 3575 84690
rect -960 84632 3514 84688
rect 3570 84632 3575 84688
rect -960 84630 3575 84632
rect -960 84540 480 84630
rect 3509 84627 3575 84630
rect 59445 82786 59511 82789
rect 244273 82786 244339 82789
rect 59445 82784 60076 82786
rect 59445 82728 59450 82784
rect 59506 82728 60076 82784
rect 59445 82726 60076 82728
rect 224388 82784 244339 82786
rect 224388 82728 244278 82784
rect 244334 82728 244339 82784
rect 224388 82726 244339 82728
rect 59445 82723 59511 82726
rect 244273 82723 244339 82726
rect 57605 80066 57671 80069
rect 226977 80066 227043 80069
rect 57605 80064 60076 80066
rect 57605 80008 57610 80064
rect 57666 80008 60076 80064
rect 57605 80006 60076 80008
rect 224388 80064 227043 80066
rect 224388 80008 226982 80064
rect 227038 80008 227043 80064
rect 224388 80006 227043 80008
rect 57605 80003 57671 80006
rect 226977 80003 227043 80006
rect 57605 77346 57671 77349
rect 233509 77346 233575 77349
rect 57605 77344 60076 77346
rect 57605 77288 57610 77344
rect 57666 77288 60076 77344
rect 57605 77286 60076 77288
rect 224388 77344 233575 77346
rect 224388 77288 233514 77344
rect 233570 77288 233575 77344
rect 224388 77286 233575 77288
rect 57605 77283 57671 77286
rect 233509 77283 233575 77286
rect 57605 74626 57671 74629
rect 228817 74626 228883 74629
rect 57605 74624 60076 74626
rect 57605 74568 57610 74624
rect 57666 74568 60076 74624
rect 57605 74566 60076 74568
rect 224388 74624 228883 74626
rect 224388 74568 228822 74624
rect 228878 74568 228883 74624
rect 224388 74566 228883 74568
rect 57605 74563 57671 74566
rect 228817 74563 228883 74566
rect 226425 73130 226491 73133
rect 235257 73130 235323 73133
rect 226425 73128 235323 73130
rect 226425 73072 226430 73128
rect 226486 73072 235262 73128
rect 235318 73072 235323 73128
rect 226425 73070 235323 73072
rect 226425 73067 226491 73070
rect 235257 73067 235323 73070
rect 583520 72994 584960 73084
rect 583342 72934 584960 72994
rect 583342 72858 583402 72934
rect 583520 72858 584960 72934
rect 583342 72844 584960 72858
rect 583342 72798 583586 72844
rect 59721 72042 59787 72045
rect 226425 72042 226491 72045
rect 59721 72040 60076 72042
rect 59721 71984 59726 72040
rect 59782 71984 60076 72040
rect 59721 71982 60076 71984
rect 224388 72040 226491 72042
rect 224388 71984 226430 72040
rect 226486 71984 226491 72040
rect 224388 71982 226491 71984
rect 59721 71979 59787 71982
rect 226425 71979 226491 71982
rect 232589 71906 232655 71909
rect 583526 71906 583586 72798
rect 232589 71904 583586 71906
rect 232589 71848 232594 71904
rect 232650 71848 583586 71904
rect 232589 71846 583586 71848
rect 232589 71843 232655 71846
rect -960 71634 480 71724
rect 3509 71634 3575 71637
rect -960 71632 3575 71634
rect -960 71576 3514 71632
rect 3570 71576 3575 71632
rect -960 71574 3575 71576
rect -960 71484 480 71574
rect 3509 71571 3575 71574
rect 57605 69322 57671 69325
rect 226558 69322 226564 69324
rect 57605 69320 60076 69322
rect 57605 69264 57610 69320
rect 57666 69264 60076 69320
rect 57605 69262 60076 69264
rect 224388 69262 226564 69322
rect 57605 69259 57671 69262
rect 226558 69260 226564 69262
rect 226628 69260 226634 69324
rect 56225 66602 56291 66605
rect 233693 66602 233759 66605
rect 56225 66600 60076 66602
rect 56225 66544 56230 66600
rect 56286 66544 60076 66600
rect 56225 66542 60076 66544
rect 224388 66600 233759 66602
rect 224388 66544 233698 66600
rect 233754 66544 233759 66600
rect 224388 66542 233759 66544
rect 56225 66539 56291 66542
rect 233693 66539 233759 66542
rect 226793 63882 226859 63885
rect 224388 63880 226859 63882
rect 60598 63612 60658 63852
rect 224388 63824 226798 63880
rect 226854 63824 226859 63880
rect 224388 63822 226859 63824
rect 226793 63819 226859 63822
rect 60590 63548 60596 63612
rect 60660 63548 60666 63612
rect 59169 61298 59235 61301
rect 231945 61298 232011 61301
rect 59169 61296 60076 61298
rect 59169 61240 59174 61296
rect 59230 61240 60076 61296
rect 59169 61238 60076 61240
rect 224388 61296 232011 61298
rect 224388 61240 231950 61296
rect 232006 61240 232011 61296
rect 224388 61238 232011 61240
rect 59169 61235 59235 61238
rect 231945 61235 232011 61238
rect 60590 60284 60596 60348
rect 60660 60346 60666 60348
rect 357433 60346 357499 60349
rect 60660 60344 357499 60346
rect 60660 60288 357438 60344
rect 357494 60288 357499 60344
rect 60660 60286 357499 60288
rect 60660 60284 60666 60286
rect 357433 60283 357499 60286
rect 221733 60210 221799 60213
rect 224585 60210 224651 60213
rect 221733 60208 224651 60210
rect 221733 60152 221738 60208
rect 221794 60152 224590 60208
rect 224646 60152 224651 60208
rect 221733 60150 224651 60152
rect 221733 60147 221799 60150
rect 224585 60147 224651 60150
rect 222929 60074 222995 60077
rect 225505 60074 225571 60077
rect 222929 60072 225571 60074
rect 222929 60016 222934 60072
rect 222990 60016 225510 60072
rect 225566 60016 225571 60072
rect 222929 60014 225571 60016
rect 222929 60011 222995 60014
rect 225505 60011 225571 60014
rect 223297 59938 223363 59941
rect 225781 59938 225847 59941
rect 223297 59936 225847 59938
rect 223297 59880 223302 59936
rect 223358 59880 225786 59936
rect 225842 59880 225847 59936
rect 223297 59878 225847 59880
rect 223297 59875 223363 59878
rect 225781 59875 225847 59878
rect 580165 59666 580231 59669
rect 583520 59666 584960 59756
rect 580165 59664 584960 59666
rect 580165 59608 580170 59664
rect 580226 59608 584960 59664
rect 580165 59606 584960 59608
rect 580165 59603 580231 59606
rect 583520 59516 584960 59606
rect 212349 59394 212415 59397
rect 224953 59394 225019 59397
rect 212349 59392 225019 59394
rect 212349 59336 212354 59392
rect 212410 59336 224958 59392
rect 225014 59336 225019 59392
rect 212349 59334 225019 59336
rect 212349 59331 212415 59334
rect 224953 59331 225019 59334
rect 210233 59258 210299 59261
rect 358813 59258 358879 59261
rect 210233 59256 358879 59258
rect 210233 59200 210238 59256
rect 210294 59200 358818 59256
rect 358874 59200 358879 59256
rect 210233 59198 358879 59200
rect 210233 59195 210299 59198
rect 358813 59195 358879 59198
rect -960 58578 480 58668
rect 3049 58578 3115 58581
rect -960 58576 3115 58578
rect -960 58520 3054 58576
rect 3110 58520 3115 58576
rect -960 58518 3115 58520
rect -960 58428 480 58518
rect 3049 58515 3115 58518
rect 58709 57898 58775 57901
rect 214741 57898 214807 57901
rect 58709 57896 214807 57898
rect 58709 57840 58714 57896
rect 58770 57840 214746 57896
rect 214802 57840 214807 57896
rect 58709 57838 214807 57840
rect 58709 57835 58775 57838
rect 214741 57835 214807 57838
rect 218237 57898 218303 57901
rect 219525 57898 219591 57901
rect 218237 57896 219591 57898
rect 218237 57840 218242 57896
rect 218298 57840 219530 57896
rect 219586 57840 219591 57896
rect 218237 57838 219591 57840
rect 218237 57835 218303 57838
rect 219525 57835 219591 57838
rect 219709 57898 219775 57901
rect 225597 57898 225663 57901
rect 219709 57896 225663 57898
rect 219709 57840 219714 57896
rect 219770 57840 225602 57896
rect 225658 57840 225663 57896
rect 219709 57838 225663 57840
rect 219709 57835 219775 57838
rect 225597 57835 225663 57838
rect 216489 57762 216555 57765
rect 225873 57762 225939 57765
rect 216489 57760 225939 57762
rect 216489 57704 216494 57760
rect 216550 57704 225878 57760
rect 225934 57704 225939 57760
rect 216489 57702 225939 57704
rect 216489 57699 216555 57702
rect 225873 57699 225939 57702
rect 219525 57626 219591 57629
rect 226241 57626 226307 57629
rect 219525 57624 226307 57626
rect 219525 57568 219530 57624
rect 219586 57568 226246 57624
rect 226302 57568 226307 57624
rect 219525 57566 226307 57568
rect 219525 57563 219591 57566
rect 226241 57563 226307 57566
rect 211153 57490 211219 57493
rect 224902 57490 224908 57492
rect 211153 57488 224908 57490
rect 211153 57432 211158 57488
rect 211214 57432 224908 57488
rect 211153 57430 224908 57432
rect 211153 57427 211219 57430
rect 224902 57428 224908 57430
rect 224972 57428 224978 57492
rect 207289 57354 207355 57357
rect 226006 57354 226012 57356
rect 207289 57352 226012 57354
rect 207289 57296 207294 57352
rect 207350 57296 226012 57352
rect 207289 57294 226012 57296
rect 207289 57291 207355 57294
rect 226006 57292 226012 57294
rect 226076 57292 226082 57356
rect 208761 57218 208827 57221
rect 356513 57218 356579 57221
rect 208761 57216 356579 57218
rect 208761 57160 208766 57216
rect 208822 57160 356518 57216
rect 356574 57160 356579 57216
rect 208761 57158 356579 57160
rect 208761 57155 208827 57158
rect 356513 57155 356579 57158
rect 213821 57082 213887 57085
rect 225321 57082 225387 57085
rect 213821 57080 225387 57082
rect 213821 57024 213826 57080
rect 213882 57024 225326 57080
rect 225382 57024 225387 57080
rect 213821 57022 225387 57024
rect 213821 57019 213887 57022
rect 225321 57019 225387 57022
rect 208485 56946 208551 56949
rect 224902 56946 224908 56948
rect 208485 56944 224908 56946
rect 208485 56888 208490 56944
rect 208546 56888 224908 56944
rect 208485 56886 224908 56888
rect 208485 56883 208551 56886
rect 224902 56884 224908 56886
rect 224972 56884 224978 56948
rect 580165 46338 580231 46341
rect 583520 46338 584960 46428
rect 580165 46336 584960 46338
rect 580165 46280 580170 46336
rect 580226 46280 584960 46336
rect 580165 46278 584960 46280
rect 580165 46275 580231 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3509 45522 3575 45525
rect -960 45520 3575 45522
rect -960 45464 3514 45520
rect 3570 45464 3575 45520
rect -960 45462 3575 45464
rect -960 45372 480 45462
rect 3509 45459 3575 45462
rect 580165 33146 580231 33149
rect 583520 33146 584960 33236
rect 580165 33144 584960 33146
rect 580165 33088 580170 33144
rect 580226 33088 584960 33144
rect 580165 33086 584960 33088
rect 580165 33083 580231 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 3509 32466 3575 32469
rect -960 32464 3575 32466
rect -960 32408 3514 32464
rect 3570 32408 3575 32464
rect -960 32406 3575 32408
rect -960 32316 480 32406
rect 3509 32403 3575 32406
rect 580165 19818 580231 19821
rect 583520 19818 584960 19908
rect 580165 19816 584960 19818
rect 580165 19760 580170 19816
rect 580226 19760 584960 19816
rect 580165 19758 584960 19760
rect 580165 19755 580231 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3509 19410 3575 19413
rect -960 19408 3575 19410
rect -960 19352 3514 19408
rect 3570 19352 3575 19408
rect -960 19350 3575 19352
rect -960 19260 480 19350
rect 3509 19347 3575 19350
rect 580257 6626 580323 6629
rect 583520 6626 584960 6716
rect 580257 6624 584960 6626
rect -960 6490 480 6580
rect 580257 6568 580262 6624
rect 580318 6568 584960 6624
rect 580257 6566 584960 6568
rect 580257 6563 580323 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect 583520 6476 584960 6566
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
<< via3 >>
rect 218652 505140 218716 505204
rect 128676 504324 128740 504388
rect 248460 504188 248524 504252
rect 258396 503916 258460 503980
rect 256188 503780 256252 503844
rect 116164 503644 116228 503708
rect 134932 503644 134996 503708
rect 151124 503644 151188 503708
rect 178540 503644 178604 503708
rect 278452 503644 278516 503708
rect 288572 503644 288636 503708
rect 88748 503508 88812 503572
rect 96476 503568 96540 503572
rect 96476 503512 96526 503568
rect 96526 503512 96540 503568
rect 96476 503508 96540 503512
rect 98500 503568 98564 503572
rect 98500 503512 98550 503568
rect 98550 503512 98564 503568
rect 98500 503508 98564 503512
rect 101260 503568 101324 503572
rect 101260 503512 101310 503568
rect 101310 503512 101324 503568
rect 101260 503508 101324 503512
rect 103836 503568 103900 503572
rect 103836 503512 103886 503568
rect 103886 503512 103900 503568
rect 103836 503508 103900 503512
rect 106044 503508 106108 503572
rect 118188 503508 118252 503572
rect 123524 503568 123588 503572
rect 123524 503512 123574 503568
rect 123574 503512 123588 503568
rect 123524 503508 123588 503512
rect 123892 503508 123956 503572
rect 129780 503568 129844 503572
rect 129780 503512 129794 503568
rect 129794 503512 129844 503568
rect 129780 503508 129844 503512
rect 143212 503508 143276 503572
rect 144868 503508 144932 503572
rect 146524 503568 146588 503572
rect 146524 503512 146574 503568
rect 146574 503512 146588 503568
rect 146524 503508 146588 503512
rect 148364 503508 148428 503572
rect 155908 503508 155972 503572
rect 158668 503568 158732 503572
rect 158668 503512 158682 503568
rect 158682 503512 158732 503568
rect 158668 503508 158732 503512
rect 160140 503568 160204 503572
rect 160140 503512 160154 503568
rect 160154 503512 160204 503568
rect 160140 503508 160204 503512
rect 163452 503508 163516 503572
rect 165660 503568 165724 503572
rect 165660 503512 165674 503568
rect 165674 503512 165724 503568
rect 165660 503508 165724 503512
rect 251036 503508 251100 503572
rect 260972 503508 261036 503572
rect 266124 503508 266188 503572
rect 267780 503568 267844 503572
rect 267780 503512 267794 503568
rect 267794 503512 267844 503568
rect 267780 503508 267844 503512
rect 270540 503568 270604 503572
rect 270540 503512 270554 503568
rect 270554 503512 270604 503568
rect 270540 503508 270604 503512
rect 273300 503568 273364 503572
rect 273300 503512 273314 503568
rect 273314 503512 273364 503568
rect 273300 503508 273364 503512
rect 276244 503508 276308 503572
rect 280108 503568 280172 503572
rect 280108 503512 280158 503568
rect 280158 503512 280172 503568
rect 280108 503508 280172 503512
rect 285628 503568 285692 503572
rect 285628 503512 285678 503568
rect 285678 503512 285692 503568
rect 285628 503508 285692 503512
rect 290964 503508 291028 503572
rect 292620 503568 292684 503572
rect 292620 503512 292634 503568
rect 292634 503512 292684 503568
rect 292620 503508 292684 503512
rect 295380 503568 295444 503572
rect 295380 503512 295394 503568
rect 295394 503512 295444 503568
rect 295380 503508 295444 503512
rect 323348 503508 323412 503572
rect 298140 492688 298204 492692
rect 298140 492632 298154 492688
rect 298154 492632 298204 492688
rect 298140 492628 298204 492632
rect 300900 492688 300964 492692
rect 300900 492632 300914 492688
rect 300914 492632 300964 492688
rect 300900 492628 300964 492632
rect 302188 492688 302252 492692
rect 302188 492632 302238 492688
rect 302238 492632 302252 492688
rect 302188 492628 302252 492632
rect 304948 492688 305012 492692
rect 304948 492632 304998 492688
rect 304998 492632 305012 492688
rect 304948 492628 305012 492632
rect 307708 492688 307772 492692
rect 307708 492632 307758 492688
rect 307758 492632 307772 492688
rect 307708 492628 307772 492632
rect 310468 492688 310532 492692
rect 310468 492632 310518 492688
rect 310518 492632 310532 492688
rect 310468 492628 310532 492632
rect 313228 492688 313292 492692
rect 313228 492632 313278 492688
rect 313278 492632 313292 492688
rect 313228 492628 313292 492632
rect 316022 492688 316086 492692
rect 316022 492632 316038 492688
rect 316038 492632 316086 492688
rect 316022 492628 316086 492632
rect 317460 492688 317524 492692
rect 317460 492632 317474 492688
rect 317474 492632 317524 492688
rect 317460 492628 317524 492632
rect 320220 492688 320284 492692
rect 320220 492632 320234 492688
rect 320234 492632 320284 492688
rect 320220 492628 320284 492632
rect 339356 492688 339420 492692
rect 339540 492688 339604 492692
rect 339356 492632 339406 492688
rect 339406 492632 339420 492688
rect 339540 492632 339554 492688
rect 339554 492632 339604 492688
rect 339356 492628 339420 492632
rect 339540 492628 339604 492632
rect 133598 491872 133662 491876
rect 133598 491816 133602 491872
rect 133602 491816 133658 491872
rect 133658 491816 133662 491872
rect 133598 491812 133662 491816
rect 153010 491736 153074 491740
rect 153010 491680 153014 491736
rect 153014 491680 153070 491736
rect 153070 491680 153074 491736
rect 153010 491676 153074 491680
rect 108298 491056 108362 491060
rect 108298 491000 108302 491056
rect 108302 491000 108358 491056
rect 108358 491000 108362 491056
rect 108298 490996 108362 491000
rect 89530 490376 89594 490380
rect 89530 490320 89534 490376
rect 89534 490320 89590 490376
rect 89590 490320 89594 490376
rect 89530 490316 89594 490320
rect 91554 490376 91618 490380
rect 91554 490320 91558 490376
rect 91558 490320 91614 490376
rect 91614 490320 91618 490376
rect 91554 490316 91618 490320
rect 111978 488336 112042 488340
rect 111978 488280 111982 488336
rect 111982 488280 112038 488336
rect 112038 488280 112042 488336
rect 111978 488276 112042 488280
rect 326614 488336 326678 488340
rect 326614 488280 326618 488336
rect 326618 488280 326674 488336
rect 326674 488280 326678 488336
rect 326614 488276 326678 488280
rect 253290 487656 253354 487660
rect 253290 487600 253294 487656
rect 253294 487600 253350 487656
rect 253350 487600 253354 487656
rect 253290 487596 253354 487600
rect 263686 487656 263750 487660
rect 263686 487600 263690 487656
rect 263690 487600 263746 487656
rect 263746 487600 263750 487656
rect 263686 487596 263750 487600
rect 284386 487656 284450 487660
rect 284386 487600 284390 487656
rect 284390 487600 284446 487656
rect 284446 487600 284450 487656
rect 284386 487596 284450 487600
rect 196756 486296 196820 486300
rect 196756 486240 196770 486296
rect 196770 486240 196820 486296
rect 196756 486236 196820 486240
rect 219756 486024 219820 486028
rect 219756 485968 219806 486024
rect 219806 485968 219820 486024
rect 219756 485964 219820 485968
rect 356836 485480 356900 485484
rect 356836 485424 356850 485480
rect 356850 485424 356900 485480
rect 356836 485420 356900 485424
rect 118510 485208 118574 485212
rect 118510 485152 118514 485208
rect 118514 485152 118570 485208
rect 118570 485152 118574 485208
rect 118510 485148 118574 485152
rect 143028 484120 143092 484124
rect 143028 484064 143078 484120
rect 143078 484064 143092 484120
rect 143028 484060 143092 484064
rect 180196 484120 180260 484124
rect 180196 484064 180246 484120
rect 180246 484064 180260 484120
rect 180196 484060 180260 484064
rect 111380 483712 111444 483716
rect 111380 483656 111430 483712
rect 111430 483656 111444 483712
rect 111380 483652 111444 483656
rect 219756 480992 219820 480996
rect 219756 480936 219806 480992
rect 219806 480936 219820 480992
rect 219756 480932 219820 480936
rect 85436 398168 85500 398172
rect 85436 398112 85486 398168
rect 85486 398112 85500 398168
rect 85436 398108 85500 398112
rect 92428 398168 92492 398172
rect 92428 398112 92442 398168
rect 92442 398112 92492 398168
rect 92428 398108 92492 398112
rect 95924 398168 95988 398172
rect 95924 398112 95974 398168
rect 95974 398112 95988 398168
rect 95924 398108 95988 398112
rect 99420 398168 99484 398172
rect 99420 398112 99434 398168
rect 99434 398112 99484 398168
rect 99420 398108 99484 398112
rect 113588 398168 113652 398172
rect 113588 398112 113638 398168
rect 113638 398112 113652 398168
rect 113588 398108 113652 398112
rect 145972 398168 146036 398172
rect 145972 398112 146022 398168
rect 146022 398112 146036 398168
rect 145972 398108 146036 398112
rect 235948 398168 236012 398172
rect 235948 398112 235998 398168
rect 235998 398112 236012 398168
rect 235948 398108 236012 398112
rect 265204 398108 265268 398172
rect 300900 398108 300964 398172
rect 315804 398168 315868 398172
rect 315804 398112 315818 398168
rect 315818 398112 315868 398168
rect 315804 398108 315868 398112
rect 325924 398168 325988 398172
rect 325924 398112 325938 398168
rect 325938 398112 325988 398168
rect 325924 398108 325988 398112
rect 226380 397972 226444 398036
rect 78260 397352 78324 397356
rect 78260 397296 78310 397352
rect 78310 397296 78324 397352
rect 78260 397292 78324 397296
rect 80652 397292 80716 397356
rect 81940 397352 82004 397356
rect 81940 397296 81990 397352
rect 81990 397296 82004 397352
rect 81940 397292 82004 397296
rect 83228 397292 83292 397356
rect 84332 397292 84396 397356
rect 87644 397352 87708 397356
rect 87644 397296 87658 397352
rect 87658 397296 87708 397352
rect 87644 397292 87708 397296
rect 88748 397352 88812 397356
rect 88748 397296 88798 397352
rect 88798 397296 88812 397352
rect 88748 397292 88812 397296
rect 90036 397292 90100 397356
rect 91324 397352 91388 397356
rect 91324 397296 91338 397352
rect 91338 397296 91388 397352
rect 91324 397292 91388 397296
rect 94452 397292 94516 397356
rect 97028 397292 97092 397356
rect 100708 397352 100772 397356
rect 100708 397296 100758 397352
rect 100758 397296 100772 397352
rect 100708 397292 100772 397296
rect 101812 397292 101876 397356
rect 104020 397352 104084 397356
rect 104020 397296 104070 397352
rect 104070 397296 104084 397352
rect 104020 397292 104084 397296
rect 106412 397352 106476 397356
rect 106412 397296 106462 397352
rect 106462 397296 106476 397352
rect 106412 397292 106476 397296
rect 109540 397352 109604 397356
rect 109540 397296 109554 397352
rect 109554 397296 109604 397352
rect 109540 397292 109604 397296
rect 111196 397352 111260 397356
rect 111196 397296 111246 397352
rect 111246 397296 111260 397352
rect 111196 397292 111260 397296
rect 112116 397352 112180 397356
rect 112116 397296 112130 397352
rect 112130 397296 112180 397352
rect 112116 397292 112180 397296
rect 113220 397352 113284 397356
rect 113220 397296 113234 397352
rect 113234 397296 113284 397352
rect 113220 397292 113284 397296
rect 114324 397292 114388 397356
rect 115796 397352 115860 397356
rect 115796 397296 115846 397352
rect 115846 397296 115860 397352
rect 115796 397292 115860 397296
rect 117084 397352 117148 397356
rect 117084 397296 117134 397352
rect 117134 397296 117148 397352
rect 117084 397292 117148 397296
rect 118188 397292 118252 397356
rect 118556 397352 118620 397356
rect 118556 397296 118606 397352
rect 118606 397296 118620 397352
rect 118556 397292 118620 397296
rect 123524 397352 123588 397356
rect 123524 397296 123538 397352
rect 123538 397296 123588 397352
rect 123524 397292 123588 397296
rect 125916 397352 125980 397356
rect 125916 397296 125966 397352
rect 125966 397296 125980 397352
rect 125916 397292 125980 397296
rect 136036 397292 136100 397356
rect 138428 397352 138492 397356
rect 138428 397296 138442 397352
rect 138442 397296 138492 397352
rect 138428 397292 138492 397296
rect 155908 397292 155972 397356
rect 163452 397292 163516 397356
rect 237052 397352 237116 397356
rect 237052 397296 237066 397352
rect 237066 397296 237116 397352
rect 237052 397292 237116 397296
rect 238156 397352 238220 397356
rect 238156 397296 238170 397352
rect 238170 397296 238220 397352
rect 238156 397292 238220 397296
rect 239260 397352 239324 397356
rect 239260 397296 239274 397352
rect 239274 397296 239324 397352
rect 239260 397292 239324 397296
rect 240548 397352 240612 397356
rect 240548 397296 240562 397352
rect 240562 397296 240612 397352
rect 240548 397292 240612 397296
rect 241652 397352 241716 397356
rect 241652 397296 241666 397352
rect 241666 397296 241716 397352
rect 241652 397292 241716 397296
rect 247724 397352 247788 397356
rect 247724 397296 247738 397352
rect 247738 397296 247788 397352
rect 247724 397292 247788 397296
rect 250668 397292 250732 397356
rect 252324 397292 252388 397356
rect 253428 397292 253492 397356
rect 260604 397292 260668 397356
rect 262076 397352 262140 397356
rect 262076 397296 262090 397352
rect 262090 397296 262140 397352
rect 262076 397292 262140 397296
rect 265940 397352 266004 397356
rect 265940 397296 265954 397352
rect 265954 397296 266004 397352
rect 265940 397292 266004 397296
rect 268332 397352 268396 397356
rect 268332 397296 268346 397352
rect 268346 397296 268396 397352
rect 268332 397292 268396 397296
rect 270908 397352 270972 397356
rect 270908 397296 270922 397352
rect 270922 397296 270972 397352
rect 270908 397292 270972 397296
rect 272564 397292 272628 397356
rect 274404 397292 274468 397356
rect 276244 397352 276308 397356
rect 276244 397296 276258 397352
rect 276258 397296 276308 397352
rect 276244 397292 276308 397296
rect 276980 397292 277044 397356
rect 278084 397352 278148 397356
rect 278084 397296 278098 397352
rect 278098 397296 278148 397352
rect 278084 397292 278148 397296
rect 279004 397352 279068 397356
rect 279004 397296 279018 397352
rect 279018 397296 279068 397352
rect 279004 397292 279068 397296
rect 283788 397292 283852 397356
rect 290964 397292 291028 397356
rect 298508 397352 298572 397356
rect 298508 397296 298522 397352
rect 298522 397296 298572 397352
rect 298508 397292 298572 397296
rect 343404 397352 343468 397356
rect 343404 397296 343418 397352
rect 343418 397296 343468 397352
rect 343404 397292 343468 397296
rect 251220 397216 251284 397220
rect 251220 397160 251270 397216
rect 251270 397160 251284 397216
rect 251220 397156 251284 397160
rect 273484 397156 273548 397220
rect 258396 396884 258460 396948
rect 77156 396808 77220 396812
rect 77156 396752 77206 396808
rect 77206 396752 77220 396808
rect 77156 396748 77220 396752
rect 79548 396748 79612 396812
rect 86540 396748 86604 396812
rect 88380 396808 88444 396812
rect 88380 396752 88394 396808
rect 88394 396752 88444 396808
rect 88380 396748 88444 396752
rect 90772 396748 90836 396812
rect 93716 396808 93780 396812
rect 93716 396752 93730 396808
rect 93730 396752 93780 396808
rect 93716 396748 93780 396752
rect 96292 396808 96356 396812
rect 96292 396752 96342 396808
rect 96342 396752 96356 396808
rect 96292 396748 96356 396752
rect 98500 396748 98564 396812
rect 101076 396748 101140 396812
rect 102732 396748 102796 396812
rect 103836 396748 103900 396812
rect 105308 396748 105372 396812
rect 106044 396808 106108 396812
rect 106044 396752 106094 396808
rect 106094 396752 106108 396808
rect 106044 396748 106108 396752
rect 107516 396808 107580 396812
rect 107516 396752 107566 396808
rect 107566 396752 107580 396808
rect 107516 396748 107580 396752
rect 108804 396748 108868 396812
rect 111012 396748 111076 396812
rect 115980 396748 116044 396812
rect 119108 396748 119172 396812
rect 120764 396748 120828 396812
rect 130884 396748 130948 396812
rect 133460 396748 133524 396812
rect 140820 396808 140884 396812
rect 140820 396752 140834 396808
rect 140834 396752 140884 396808
rect 140820 396748 140884 396752
rect 143580 396748 143644 396812
rect 148548 396748 148612 396812
rect 150940 396748 151004 396812
rect 154068 396748 154132 396812
rect 158484 396748 158548 396812
rect 160876 396748 160940 396812
rect 165844 396748 165908 396812
rect 183140 396748 183204 396812
rect 183508 396808 183572 396812
rect 183508 396752 183522 396808
rect 183522 396752 183572 396808
rect 183508 396748 183572 396752
rect 242940 396808 243004 396812
rect 242940 396752 242954 396808
rect 242954 396752 243004 396808
rect 242940 396748 243004 396752
rect 244228 396748 244292 396812
rect 246436 396748 246500 396812
rect 248276 396748 248340 396812
rect 248644 396748 248708 396812
rect 250116 396748 250180 396812
rect 253612 396748 253676 396812
rect 254532 396808 254596 396812
rect 254532 396752 254546 396808
rect 254546 396752 254596 396808
rect 254532 396748 254596 396752
rect 255820 396748 255884 396812
rect 256924 396808 256988 396812
rect 256924 396752 256938 396808
rect 256938 396752 256988 396808
rect 256924 396748 256988 396752
rect 258396 396748 258460 396812
rect 259500 396808 259564 396812
rect 259500 396752 259550 396808
rect 259550 396752 259564 396808
rect 259500 396748 259564 396752
rect 260972 396808 261036 396812
rect 260972 396752 260986 396808
rect 260986 396752 261036 396808
rect 260972 396748 261036 396752
rect 262812 396748 262876 396812
rect 263548 396808 263612 396812
rect 263548 396752 263598 396808
rect 263598 396752 263612 396808
rect 263548 396748 263612 396752
rect 266308 396808 266372 396812
rect 266308 396752 266358 396808
rect 266358 396752 266372 396808
rect 266308 396748 266372 396752
rect 268700 396748 268764 396812
rect 269804 396748 269868 396812
rect 271276 396748 271340 396812
rect 273300 396808 273364 396812
rect 273300 396752 273314 396808
rect 273314 396752 273364 396808
rect 273300 396748 273364 396752
rect 275324 396748 275388 396812
rect 278452 396748 278516 396812
rect 280844 396748 280908 396812
rect 285996 396748 286060 396812
rect 288204 396748 288268 396812
rect 293356 396748 293420 396812
rect 295932 396808 295996 396812
rect 295932 396752 295946 396808
rect 295946 396752 295996 396808
rect 295932 396748 295996 396752
rect 303476 396748 303540 396812
rect 305868 396748 305932 396812
rect 308628 396748 308692 396812
rect 311020 396748 311084 396812
rect 313412 396748 313476 396812
rect 318380 396748 318444 396812
rect 320956 396748 321020 396812
rect 323348 396748 323412 396812
rect 343220 396748 343284 396812
rect 76052 396612 76116 396676
rect 93348 396612 93412 396676
rect 98132 396612 98196 396676
rect 108252 396612 108316 396676
rect 245332 396612 245396 396676
rect 256188 396612 256252 396676
rect 263916 396612 263980 396676
rect 267596 396612 267660 396676
rect 128676 396068 128740 396132
rect 226748 242116 226812 242180
rect 228404 235996 228468 236060
rect 228220 233276 228284 233340
rect 224908 233004 224972 233068
rect 226932 232460 226996 232524
rect 218652 230284 218716 230348
rect 224908 230284 224972 230348
rect 226564 227836 226628 227900
rect 226012 227428 226076 227492
rect 227300 220900 227364 220964
rect 227300 219540 227364 219604
rect 228404 218044 228468 218108
rect 226748 114956 226812 115020
rect 228220 111828 228284 111892
rect 226932 106932 226996 106996
rect 226380 85308 226444 85372
rect 226564 69260 226628 69324
rect 60596 63548 60660 63612
rect 60596 60284 60660 60348
rect 224908 57428 224972 57492
rect 226012 57292 226076 57356
rect 224908 56884 224972 56948
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 680614 -8106 711002
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 -8106 680614
rect -8726 680294 -8106 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 -8106 680294
rect -8726 644614 -8106 680058
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 -8106 644614
rect -8726 644294 -8106 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 -8106 644294
rect -8726 608614 -8106 644058
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 -8106 608614
rect -8726 608294 -8106 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 -8106 608294
rect -8726 572614 -8106 608058
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 -8106 572614
rect -8726 572294 -8106 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 -8106 572294
rect -8726 536614 -8106 572058
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 -8106 536614
rect -8726 536294 -8106 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 -8106 536294
rect -8726 500614 -8106 536058
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 -8106 500614
rect -8726 500294 -8106 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 -8106 500294
rect -8726 464614 -8106 500058
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 -8106 464614
rect -8726 464294 -8106 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 -8106 464294
rect -8726 428614 -8106 464058
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 -8106 428614
rect -8726 428294 -8106 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 -8106 428294
rect -8726 392614 -8106 428058
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 -8106 392614
rect -8726 392294 -8106 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 -8106 392294
rect -8726 356614 -8106 392058
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 -8106 356614
rect -8726 356294 -8106 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 -8106 356294
rect -8726 320614 -8106 356058
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 -8106 320614
rect -8726 320294 -8106 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 -8106 320294
rect -8726 284614 -8106 320058
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 -8106 284614
rect -8726 284294 -8106 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 -8106 284294
rect -8726 248614 -8106 284058
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 -8106 248614
rect -8726 248294 -8106 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 -8106 248294
rect -8726 212614 -8106 248058
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 -8106 212614
rect -8726 212294 -8106 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 -8106 212294
rect -8726 176614 -8106 212058
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 -8106 176614
rect -8726 176294 -8106 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 -8106 176294
rect -8726 140614 -8106 176058
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 -8106 140614
rect -8726 140294 -8106 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 -8106 140294
rect -8726 104614 -8106 140058
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 -8106 104614
rect -8726 104294 -8106 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 -8106 104294
rect -8726 68614 -8106 104058
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 -8106 68614
rect -8726 68294 -8106 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 -8106 68294
rect -8726 32614 -8106 68058
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 -8106 32614
rect -8726 32294 -8106 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 -8106 32294
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 13574 710598
rect 12954 710278 13574 710362
rect 12954 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 13574 710278
rect -7766 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 -7146 698614
rect -7766 698294 -7146 698378
rect -7766 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 -7146 698294
rect -7766 662614 -7146 698058
rect -7766 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 -7146 662614
rect -7766 662294 -7146 662378
rect -7766 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 -7146 662294
rect -7766 626614 -7146 662058
rect -7766 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 -7146 626614
rect -7766 626294 -7146 626378
rect -7766 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 -7146 626294
rect -7766 590614 -7146 626058
rect -7766 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 -7146 590614
rect -7766 590294 -7146 590378
rect -7766 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 -7146 590294
rect -7766 554614 -7146 590058
rect -7766 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 -7146 554614
rect -7766 554294 -7146 554378
rect -7766 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 -7146 554294
rect -7766 518614 -7146 554058
rect -7766 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 -7146 518614
rect -7766 518294 -7146 518378
rect -7766 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 -7146 518294
rect -7766 482614 -7146 518058
rect -7766 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 -7146 482614
rect -7766 482294 -7146 482378
rect -7766 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 -7146 482294
rect -7766 446614 -7146 482058
rect -7766 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 -7146 446614
rect -7766 446294 -7146 446378
rect -7766 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 -7146 446294
rect -7766 410614 -7146 446058
rect -7766 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 -7146 410614
rect -7766 410294 -7146 410378
rect -7766 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 -7146 410294
rect -7766 374614 -7146 410058
rect -7766 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 -7146 374614
rect -7766 374294 -7146 374378
rect -7766 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 -7146 374294
rect -7766 338614 -7146 374058
rect -7766 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 -7146 338614
rect -7766 338294 -7146 338378
rect -7766 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 -7146 338294
rect -7766 302614 -7146 338058
rect -7766 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 -7146 302614
rect -7766 302294 -7146 302378
rect -7766 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 -7146 302294
rect -7766 266614 -7146 302058
rect -7766 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 -7146 266614
rect -7766 266294 -7146 266378
rect -7766 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 -7146 266294
rect -7766 230614 -7146 266058
rect -7766 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 -7146 230614
rect -7766 230294 -7146 230378
rect -7766 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 -7146 230294
rect -7766 194614 -7146 230058
rect -7766 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 -7146 194614
rect -7766 194294 -7146 194378
rect -7766 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 -7146 194294
rect -7766 158614 -7146 194058
rect -7766 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 -7146 158614
rect -7766 158294 -7146 158378
rect -7766 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 -7146 158294
rect -7766 122614 -7146 158058
rect -7766 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 -7146 122614
rect -7766 122294 -7146 122378
rect -7766 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 -7146 122294
rect -7766 86614 -7146 122058
rect -7766 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 -7146 86614
rect -7766 86294 -7146 86378
rect -7766 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 -7146 86294
rect -7766 50614 -7146 86058
rect -7766 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 -7146 50614
rect -7766 50294 -7146 50378
rect -7766 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 -7146 50294
rect -7766 14614 -7146 50058
rect -7766 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 -7146 14614
rect -7766 14294 -7146 14378
rect -7766 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 -7146 14294
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 676894 -6186 709082
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 -6186 676894
rect -6806 676574 -6186 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 -6186 676574
rect -6806 640894 -6186 676338
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 -6186 640894
rect -6806 640574 -6186 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 -6186 640574
rect -6806 604894 -6186 640338
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 -6186 604894
rect -6806 604574 -6186 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 -6186 604574
rect -6806 568894 -6186 604338
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 -6186 568894
rect -6806 568574 -6186 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 -6186 568574
rect -6806 532894 -6186 568338
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 -6186 532894
rect -6806 532574 -6186 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 -6186 532574
rect -6806 496894 -6186 532338
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 -6186 496894
rect -6806 496574 -6186 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 -6186 496574
rect -6806 460894 -6186 496338
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 -6186 460894
rect -6806 460574 -6186 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 -6186 460574
rect -6806 424894 -6186 460338
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 -6186 424894
rect -6806 424574 -6186 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 -6186 424574
rect -6806 388894 -6186 424338
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 -6186 388894
rect -6806 388574 -6186 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 -6186 388574
rect -6806 352894 -6186 388338
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 -6186 352894
rect -6806 352574 -6186 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 -6186 352574
rect -6806 316894 -6186 352338
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 -6186 316894
rect -6806 316574 -6186 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 -6186 316574
rect -6806 280894 -6186 316338
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 -6186 280894
rect -6806 280574 -6186 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 -6186 280574
rect -6806 244894 -6186 280338
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 -6186 244894
rect -6806 244574 -6186 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 -6186 244574
rect -6806 208894 -6186 244338
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 -6186 208894
rect -6806 208574 -6186 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 -6186 208574
rect -6806 172894 -6186 208338
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 -6186 172894
rect -6806 172574 -6186 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 -6186 172574
rect -6806 136894 -6186 172338
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 -6186 136894
rect -6806 136574 -6186 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 -6186 136574
rect -6806 100894 -6186 136338
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 -6186 100894
rect -6806 100574 -6186 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 -6186 100574
rect -6806 64894 -6186 100338
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 -6186 64894
rect -6806 64574 -6186 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 -6186 64574
rect -6806 28894 -6186 64338
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 -6186 28894
rect -6806 28574 -6186 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 -6186 28574
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 9854 708678
rect 9234 708358 9854 708442
rect 9234 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 9854 708358
rect -5846 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 -5226 694894
rect -5846 694574 -5226 694658
rect -5846 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 -5226 694574
rect -5846 658894 -5226 694338
rect -5846 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 -5226 658894
rect -5846 658574 -5226 658658
rect -5846 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 -5226 658574
rect -5846 622894 -5226 658338
rect -5846 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 -5226 622894
rect -5846 622574 -5226 622658
rect -5846 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 -5226 622574
rect -5846 586894 -5226 622338
rect -5846 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 -5226 586894
rect -5846 586574 -5226 586658
rect -5846 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 -5226 586574
rect -5846 550894 -5226 586338
rect -5846 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 -5226 550894
rect -5846 550574 -5226 550658
rect -5846 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 -5226 550574
rect -5846 514894 -5226 550338
rect -5846 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 -5226 514894
rect -5846 514574 -5226 514658
rect -5846 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 -5226 514574
rect -5846 478894 -5226 514338
rect -5846 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 -5226 478894
rect -5846 478574 -5226 478658
rect -5846 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 -5226 478574
rect -5846 442894 -5226 478338
rect -5846 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 -5226 442894
rect -5846 442574 -5226 442658
rect -5846 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 -5226 442574
rect -5846 406894 -5226 442338
rect -5846 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 -5226 406894
rect -5846 406574 -5226 406658
rect -5846 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 -5226 406574
rect -5846 370894 -5226 406338
rect -5846 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 -5226 370894
rect -5846 370574 -5226 370658
rect -5846 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 -5226 370574
rect -5846 334894 -5226 370338
rect -5846 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 -5226 334894
rect -5846 334574 -5226 334658
rect -5846 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 -5226 334574
rect -5846 298894 -5226 334338
rect -5846 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 -5226 298894
rect -5846 298574 -5226 298658
rect -5846 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 -5226 298574
rect -5846 262894 -5226 298338
rect -5846 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 -5226 262894
rect -5846 262574 -5226 262658
rect -5846 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 -5226 262574
rect -5846 226894 -5226 262338
rect -5846 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 -5226 226894
rect -5846 226574 -5226 226658
rect -5846 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 -5226 226574
rect -5846 190894 -5226 226338
rect -5846 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 -5226 190894
rect -5846 190574 -5226 190658
rect -5846 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 -5226 190574
rect -5846 154894 -5226 190338
rect -5846 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 -5226 154894
rect -5846 154574 -5226 154658
rect -5846 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 -5226 154574
rect -5846 118894 -5226 154338
rect -5846 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 -5226 118894
rect -5846 118574 -5226 118658
rect -5846 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 -5226 118574
rect -5846 82894 -5226 118338
rect -5846 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 -5226 82894
rect -5846 82574 -5226 82658
rect -5846 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 -5226 82574
rect -5846 46894 -5226 82338
rect -5846 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 -5226 46894
rect -5846 46574 -5226 46658
rect -5846 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 -5226 46574
rect -5846 10894 -5226 46338
rect -5846 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 -5226 10894
rect -5846 10574 -5226 10658
rect -5846 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 -5226 10574
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 673174 -4266 707162
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 -4266 673174
rect -4886 672854 -4266 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 -4266 672854
rect -4886 637174 -4266 672618
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 -4266 637174
rect -4886 636854 -4266 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 -4266 636854
rect -4886 601174 -4266 636618
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 -4266 601174
rect -4886 600854 -4266 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 -4266 600854
rect -4886 565174 -4266 600618
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 -4266 565174
rect -4886 564854 -4266 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 -4266 564854
rect -4886 529174 -4266 564618
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 -4266 529174
rect -4886 528854 -4266 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 -4266 528854
rect -4886 493174 -4266 528618
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 -4266 493174
rect -4886 492854 -4266 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 -4266 492854
rect -4886 457174 -4266 492618
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 -4266 457174
rect -4886 456854 -4266 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 -4266 456854
rect -4886 421174 -4266 456618
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 -4266 421174
rect -4886 420854 -4266 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 -4266 420854
rect -4886 385174 -4266 420618
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 -4266 385174
rect -4886 384854 -4266 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 -4266 384854
rect -4886 349174 -4266 384618
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 -4266 349174
rect -4886 348854 -4266 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 -4266 348854
rect -4886 313174 -4266 348618
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 -4266 313174
rect -4886 312854 -4266 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 -4266 312854
rect -4886 277174 -4266 312618
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 -4266 277174
rect -4886 276854 -4266 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 -4266 276854
rect -4886 241174 -4266 276618
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 -4266 241174
rect -4886 240854 -4266 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 -4266 240854
rect -4886 205174 -4266 240618
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 -4266 205174
rect -4886 204854 -4266 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 -4266 204854
rect -4886 169174 -4266 204618
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 -4266 169174
rect -4886 168854 -4266 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 -4266 168854
rect -4886 133174 -4266 168618
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 -4266 133174
rect -4886 132854 -4266 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 -4266 132854
rect -4886 97174 -4266 132618
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 -4266 97174
rect -4886 96854 -4266 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 -4266 96854
rect -4886 61174 -4266 96618
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 -4266 61174
rect -4886 60854 -4266 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 -4266 60854
rect -4886 25174 -4266 60618
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 -4266 25174
rect -4886 24854 -4266 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 -4266 24854
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 6134 706758
rect 5514 706438 6134 706522
rect 5514 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 6134 706438
rect -3926 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 -3306 691174
rect -3926 690854 -3306 690938
rect -3926 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 -3306 690854
rect -3926 655174 -3306 690618
rect -3926 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 -3306 655174
rect -3926 654854 -3306 654938
rect -3926 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 -3306 654854
rect -3926 619174 -3306 654618
rect -3926 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 -3306 619174
rect -3926 618854 -3306 618938
rect -3926 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 -3306 618854
rect -3926 583174 -3306 618618
rect -3926 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 -3306 583174
rect -3926 582854 -3306 582938
rect -3926 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 -3306 582854
rect -3926 547174 -3306 582618
rect -3926 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 -3306 547174
rect -3926 546854 -3306 546938
rect -3926 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 -3306 546854
rect -3926 511174 -3306 546618
rect -3926 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 -3306 511174
rect -3926 510854 -3306 510938
rect -3926 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 -3306 510854
rect -3926 475174 -3306 510618
rect -3926 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 -3306 475174
rect -3926 474854 -3306 474938
rect -3926 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 -3306 474854
rect -3926 439174 -3306 474618
rect -3926 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 -3306 439174
rect -3926 438854 -3306 438938
rect -3926 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 -3306 438854
rect -3926 403174 -3306 438618
rect -3926 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 -3306 403174
rect -3926 402854 -3306 402938
rect -3926 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 -3306 402854
rect -3926 367174 -3306 402618
rect -3926 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 -3306 367174
rect -3926 366854 -3306 366938
rect -3926 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 -3306 366854
rect -3926 331174 -3306 366618
rect -3926 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 -3306 331174
rect -3926 330854 -3306 330938
rect -3926 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 -3306 330854
rect -3926 295174 -3306 330618
rect -3926 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 -3306 295174
rect -3926 294854 -3306 294938
rect -3926 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 -3306 294854
rect -3926 259174 -3306 294618
rect -3926 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 -3306 259174
rect -3926 258854 -3306 258938
rect -3926 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 -3306 258854
rect -3926 223174 -3306 258618
rect -3926 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 -3306 223174
rect -3926 222854 -3306 222938
rect -3926 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 -3306 222854
rect -3926 187174 -3306 222618
rect -3926 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 -3306 187174
rect -3926 186854 -3306 186938
rect -3926 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 -3306 186854
rect -3926 151174 -3306 186618
rect -3926 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 -3306 151174
rect -3926 150854 -3306 150938
rect -3926 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 -3306 150854
rect -3926 115174 -3306 150618
rect -3926 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 -3306 115174
rect -3926 114854 -3306 114938
rect -3926 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 -3306 114854
rect -3926 79174 -3306 114618
rect -3926 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 -3306 79174
rect -3926 78854 -3306 78938
rect -3926 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 -3306 78854
rect -3926 43174 -3306 78618
rect -3926 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 -3306 43174
rect -3926 42854 -3306 42938
rect -3926 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 -3306 42854
rect -3926 7174 -3306 42618
rect -3926 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 -3306 7174
rect -3926 6854 -3306 6938
rect -3926 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 -3306 6854
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 5514 691174 6134 706202
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 6618
rect 5514 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 6134 -2266
rect 5514 -2586 6134 -2502
rect 5514 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 6134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect 9234 694894 9854 708122
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 10338
rect 9234 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 9854 -4186
rect 9234 -4506 9854 -4422
rect 9234 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 9854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect 12954 698614 13574 710042
rect 30954 711558 31574 711590
rect 30954 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 31574 711558
rect 30954 711238 31574 711322
rect 30954 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 31574 711238
rect 27234 709638 27854 709670
rect 27234 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 27854 709638
rect 27234 709318 27854 709402
rect 27234 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 27854 709318
rect 23514 707718 24134 707750
rect 23514 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 24134 707718
rect 23514 707398 24134 707482
rect 23514 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 24134 707398
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 14058
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 19794 669454 20414 705242
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -1306 20414 20898
rect 19794 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 20414 -1306
rect 19794 -1626 20414 -1542
rect 19794 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 20414 -1626
rect 19794 -1894 20414 -1862
rect 23514 673174 24134 707162
rect 23514 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 24134 673174
rect 23514 672854 24134 672938
rect 23514 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 24134 672854
rect 23514 637174 24134 672618
rect 23514 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 24134 637174
rect 23514 636854 24134 636938
rect 23514 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 24134 636854
rect 23514 601174 24134 636618
rect 23514 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 24134 601174
rect 23514 600854 24134 600938
rect 23514 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 24134 600854
rect 23514 565174 24134 600618
rect 23514 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 24134 565174
rect 23514 564854 24134 564938
rect 23514 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 24134 564854
rect 23514 529174 24134 564618
rect 23514 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 24134 529174
rect 23514 528854 24134 528938
rect 23514 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 24134 528854
rect 23514 493174 24134 528618
rect 23514 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 24134 493174
rect 23514 492854 24134 492938
rect 23514 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 24134 492854
rect 23514 457174 24134 492618
rect 23514 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 24134 457174
rect 23514 456854 24134 456938
rect 23514 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 24134 456854
rect 23514 421174 24134 456618
rect 23514 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 24134 421174
rect 23514 420854 24134 420938
rect 23514 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 24134 420854
rect 23514 385174 24134 420618
rect 23514 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 24134 385174
rect 23514 384854 24134 384938
rect 23514 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 24134 384854
rect 23514 349174 24134 384618
rect 23514 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 24134 349174
rect 23514 348854 24134 348938
rect 23514 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 24134 348854
rect 23514 313174 24134 348618
rect 23514 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 24134 313174
rect 23514 312854 24134 312938
rect 23514 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 24134 312854
rect 23514 277174 24134 312618
rect 23514 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 24134 277174
rect 23514 276854 24134 276938
rect 23514 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 24134 276854
rect 23514 241174 24134 276618
rect 23514 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 24134 241174
rect 23514 240854 24134 240938
rect 23514 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 24134 240854
rect 23514 205174 24134 240618
rect 23514 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 24134 205174
rect 23514 204854 24134 204938
rect 23514 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 24134 204854
rect 23514 169174 24134 204618
rect 23514 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 24134 169174
rect 23514 168854 24134 168938
rect 23514 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 24134 168854
rect 23514 133174 24134 168618
rect 23514 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 24134 133174
rect 23514 132854 24134 132938
rect 23514 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 24134 132854
rect 23514 97174 24134 132618
rect 23514 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 24134 97174
rect 23514 96854 24134 96938
rect 23514 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 24134 96854
rect 23514 61174 24134 96618
rect 23514 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 24134 61174
rect 23514 60854 24134 60938
rect 23514 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 24134 60854
rect 23514 25174 24134 60618
rect 23514 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 24134 25174
rect 23514 24854 24134 24938
rect 23514 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 24134 24854
rect 23514 -3226 24134 24618
rect 23514 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 24134 -3226
rect 23514 -3546 24134 -3462
rect 23514 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 24134 -3546
rect 23514 -3814 24134 -3782
rect 27234 676894 27854 709082
rect 27234 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 27854 676894
rect 27234 676574 27854 676658
rect 27234 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 27854 676574
rect 27234 640894 27854 676338
rect 27234 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 27854 640894
rect 27234 640574 27854 640658
rect 27234 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 27854 640574
rect 27234 604894 27854 640338
rect 27234 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 27854 604894
rect 27234 604574 27854 604658
rect 27234 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 27854 604574
rect 27234 568894 27854 604338
rect 27234 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 27854 568894
rect 27234 568574 27854 568658
rect 27234 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 27854 568574
rect 27234 532894 27854 568338
rect 27234 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 27854 532894
rect 27234 532574 27854 532658
rect 27234 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 27854 532574
rect 27234 496894 27854 532338
rect 27234 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 27854 496894
rect 27234 496574 27854 496658
rect 27234 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 27854 496574
rect 27234 460894 27854 496338
rect 27234 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 27854 460894
rect 27234 460574 27854 460658
rect 27234 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 27854 460574
rect 27234 424894 27854 460338
rect 27234 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 27854 424894
rect 27234 424574 27854 424658
rect 27234 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 27854 424574
rect 27234 388894 27854 424338
rect 27234 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 27854 388894
rect 27234 388574 27854 388658
rect 27234 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 27854 388574
rect 27234 352894 27854 388338
rect 27234 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 27854 352894
rect 27234 352574 27854 352658
rect 27234 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 27854 352574
rect 27234 316894 27854 352338
rect 27234 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 27854 316894
rect 27234 316574 27854 316658
rect 27234 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 27854 316574
rect 27234 280894 27854 316338
rect 27234 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 27854 280894
rect 27234 280574 27854 280658
rect 27234 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 27854 280574
rect 27234 244894 27854 280338
rect 27234 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 27854 244894
rect 27234 244574 27854 244658
rect 27234 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 27854 244574
rect 27234 208894 27854 244338
rect 27234 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 27854 208894
rect 27234 208574 27854 208658
rect 27234 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 27854 208574
rect 27234 172894 27854 208338
rect 27234 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 27854 172894
rect 27234 172574 27854 172658
rect 27234 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 27854 172574
rect 27234 136894 27854 172338
rect 27234 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 27854 136894
rect 27234 136574 27854 136658
rect 27234 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 27854 136574
rect 27234 100894 27854 136338
rect 27234 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 27854 100894
rect 27234 100574 27854 100658
rect 27234 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 27854 100574
rect 27234 64894 27854 100338
rect 27234 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 27854 64894
rect 27234 64574 27854 64658
rect 27234 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 27854 64574
rect 27234 28894 27854 64338
rect 27234 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 27854 28894
rect 27234 28574 27854 28658
rect 27234 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 27854 28574
rect 27234 -5146 27854 28338
rect 27234 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 27854 -5146
rect 27234 -5466 27854 -5382
rect 27234 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 27854 -5466
rect 27234 -5734 27854 -5702
rect 30954 680614 31574 711002
rect 48954 710598 49574 711590
rect 48954 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 49574 710598
rect 48954 710278 49574 710362
rect 48954 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 49574 710278
rect 45234 708678 45854 709670
rect 45234 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 45854 708678
rect 45234 708358 45854 708442
rect 45234 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 45854 708358
rect 41514 706758 42134 707750
rect 41514 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 42134 706758
rect 41514 706438 42134 706522
rect 41514 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 42134 706438
rect 30954 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 31574 680614
rect 30954 680294 31574 680378
rect 30954 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 31574 680294
rect 30954 644614 31574 680058
rect 30954 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 31574 644614
rect 30954 644294 31574 644378
rect 30954 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 31574 644294
rect 30954 608614 31574 644058
rect 30954 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 31574 608614
rect 30954 608294 31574 608378
rect 30954 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 31574 608294
rect 30954 572614 31574 608058
rect 30954 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 31574 572614
rect 30954 572294 31574 572378
rect 30954 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 31574 572294
rect 30954 536614 31574 572058
rect 30954 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 31574 536614
rect 30954 536294 31574 536378
rect 30954 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 31574 536294
rect 30954 500614 31574 536058
rect 30954 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 31574 500614
rect 30954 500294 31574 500378
rect 30954 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 31574 500294
rect 30954 464614 31574 500058
rect 30954 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 31574 464614
rect 30954 464294 31574 464378
rect 30954 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 31574 464294
rect 30954 428614 31574 464058
rect 30954 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 31574 428614
rect 30954 428294 31574 428378
rect 30954 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 31574 428294
rect 30954 392614 31574 428058
rect 30954 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 31574 392614
rect 30954 392294 31574 392378
rect 30954 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 31574 392294
rect 30954 356614 31574 392058
rect 30954 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 31574 356614
rect 30954 356294 31574 356378
rect 30954 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 31574 356294
rect 30954 320614 31574 356058
rect 30954 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 31574 320614
rect 30954 320294 31574 320378
rect 30954 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 31574 320294
rect 30954 284614 31574 320058
rect 30954 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 31574 284614
rect 30954 284294 31574 284378
rect 30954 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 31574 284294
rect 30954 248614 31574 284058
rect 30954 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 31574 248614
rect 30954 248294 31574 248378
rect 30954 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 31574 248294
rect 30954 212614 31574 248058
rect 30954 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 31574 212614
rect 30954 212294 31574 212378
rect 30954 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 31574 212294
rect 30954 176614 31574 212058
rect 30954 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 31574 176614
rect 30954 176294 31574 176378
rect 30954 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 31574 176294
rect 30954 140614 31574 176058
rect 30954 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 31574 140614
rect 30954 140294 31574 140378
rect 30954 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 31574 140294
rect 30954 104614 31574 140058
rect 30954 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 31574 104614
rect 30954 104294 31574 104378
rect 30954 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 31574 104294
rect 30954 68614 31574 104058
rect 30954 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 31574 68614
rect 30954 68294 31574 68378
rect 30954 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 31574 68294
rect 30954 32614 31574 68058
rect 30954 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 31574 32614
rect 30954 32294 31574 32378
rect 30954 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 31574 32294
rect 12954 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 13574 -6106
rect 12954 -6426 13574 -6342
rect 12954 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 13574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 32058
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 41514 691174 42134 706202
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 655174 42134 690618
rect 41514 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 42134 655174
rect 41514 654854 42134 654938
rect 41514 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 42134 654854
rect 41514 619174 42134 654618
rect 41514 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 42134 619174
rect 41514 618854 42134 618938
rect 41514 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 42134 618854
rect 41514 583174 42134 618618
rect 41514 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 42134 583174
rect 41514 582854 42134 582938
rect 41514 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 42134 582854
rect 41514 547174 42134 582618
rect 41514 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 42134 547174
rect 41514 546854 42134 546938
rect 41514 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 42134 546854
rect 41514 511174 42134 546618
rect 41514 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 42134 511174
rect 41514 510854 42134 510938
rect 41514 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 42134 510854
rect 41514 475174 42134 510618
rect 41514 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 42134 475174
rect 41514 474854 42134 474938
rect 41514 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 42134 474854
rect 41514 439174 42134 474618
rect 41514 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 42134 439174
rect 41514 438854 42134 438938
rect 41514 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 42134 438854
rect 41514 403174 42134 438618
rect 41514 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 42134 403174
rect 41514 402854 42134 402938
rect 41514 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 42134 402854
rect 41514 367174 42134 402618
rect 41514 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 42134 367174
rect 41514 366854 42134 366938
rect 41514 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 42134 366854
rect 41514 331174 42134 366618
rect 41514 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 42134 331174
rect 41514 330854 42134 330938
rect 41514 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 42134 330854
rect 41514 295174 42134 330618
rect 41514 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 42134 295174
rect 41514 294854 42134 294938
rect 41514 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 42134 294854
rect 41514 259174 42134 294618
rect 41514 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 42134 259174
rect 41514 258854 42134 258938
rect 41514 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 42134 258854
rect 41514 223174 42134 258618
rect 41514 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 42134 223174
rect 41514 222854 42134 222938
rect 41514 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 42134 222854
rect 41514 187174 42134 222618
rect 41514 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 42134 187174
rect 41514 186854 42134 186938
rect 41514 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 42134 186854
rect 41514 151174 42134 186618
rect 41514 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 42134 151174
rect 41514 150854 42134 150938
rect 41514 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 42134 150854
rect 41514 115174 42134 150618
rect 41514 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 42134 115174
rect 41514 114854 42134 114938
rect 41514 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 42134 114854
rect 41514 79174 42134 114618
rect 41514 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 42134 79174
rect 41514 78854 42134 78938
rect 41514 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 42134 78854
rect 41514 43174 42134 78618
rect 41514 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 42134 43174
rect 41514 42854 42134 42938
rect 41514 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 42134 42854
rect 41514 7174 42134 42618
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -2266 42134 6618
rect 41514 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 42134 -2266
rect 41514 -2586 42134 -2502
rect 41514 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 42134 -2586
rect 41514 -3814 42134 -2822
rect 45234 694894 45854 708122
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 658894 45854 694338
rect 45234 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 45854 658894
rect 45234 658574 45854 658658
rect 45234 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 45854 658574
rect 45234 622894 45854 658338
rect 45234 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 45854 622894
rect 45234 622574 45854 622658
rect 45234 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 45854 622574
rect 45234 586894 45854 622338
rect 45234 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 45854 586894
rect 45234 586574 45854 586658
rect 45234 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 45854 586574
rect 45234 550894 45854 586338
rect 45234 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 45854 550894
rect 45234 550574 45854 550658
rect 45234 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 45854 550574
rect 45234 514894 45854 550338
rect 45234 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 45854 514894
rect 45234 514574 45854 514658
rect 45234 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 45854 514574
rect 45234 478894 45854 514338
rect 45234 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 45854 478894
rect 45234 478574 45854 478658
rect 45234 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 45854 478574
rect 45234 442894 45854 478338
rect 45234 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 45854 442894
rect 45234 442574 45854 442658
rect 45234 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 45854 442574
rect 45234 406894 45854 442338
rect 45234 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 45854 406894
rect 45234 406574 45854 406658
rect 45234 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 45854 406574
rect 45234 370894 45854 406338
rect 45234 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 45854 370894
rect 45234 370574 45854 370658
rect 45234 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 45854 370574
rect 45234 334894 45854 370338
rect 45234 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 45854 334894
rect 45234 334574 45854 334658
rect 45234 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 45854 334574
rect 45234 298894 45854 334338
rect 45234 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 45854 298894
rect 45234 298574 45854 298658
rect 45234 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 45854 298574
rect 45234 262894 45854 298338
rect 45234 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 45854 262894
rect 45234 262574 45854 262658
rect 45234 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 45854 262574
rect 45234 226894 45854 262338
rect 45234 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 45854 226894
rect 45234 226574 45854 226658
rect 45234 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 45854 226574
rect 45234 190894 45854 226338
rect 45234 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 45854 190894
rect 45234 190574 45854 190658
rect 45234 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 45854 190574
rect 45234 154894 45854 190338
rect 45234 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 45854 154894
rect 45234 154574 45854 154658
rect 45234 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 45854 154574
rect 45234 118894 45854 154338
rect 45234 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 45854 118894
rect 45234 118574 45854 118658
rect 45234 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 45854 118574
rect 45234 82894 45854 118338
rect 45234 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 45854 82894
rect 45234 82574 45854 82658
rect 45234 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 45854 82574
rect 45234 46894 45854 82338
rect 45234 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 45854 46894
rect 45234 46574 45854 46658
rect 45234 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 45854 46574
rect 45234 10894 45854 46338
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -4186 45854 10338
rect 45234 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 45854 -4186
rect 45234 -4506 45854 -4422
rect 45234 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 45854 -4506
rect 45234 -5734 45854 -4742
rect 48954 698614 49574 710042
rect 66954 711558 67574 711590
rect 66954 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 67574 711558
rect 66954 711238 67574 711322
rect 66954 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 67574 711238
rect 63234 709638 63854 709670
rect 63234 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 63854 709638
rect 63234 709318 63854 709402
rect 63234 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 63854 709318
rect 59514 707718 60134 707750
rect 59514 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 60134 707718
rect 59514 707398 60134 707482
rect 59514 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 60134 707398
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 662614 49574 698058
rect 48954 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 49574 662614
rect 48954 662294 49574 662378
rect 48954 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 49574 662294
rect 48954 626614 49574 662058
rect 48954 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 49574 626614
rect 48954 626294 49574 626378
rect 48954 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 49574 626294
rect 48954 590614 49574 626058
rect 48954 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 49574 590614
rect 48954 590294 49574 590378
rect 48954 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 49574 590294
rect 48954 554614 49574 590058
rect 48954 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 49574 554614
rect 48954 554294 49574 554378
rect 48954 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 49574 554294
rect 48954 518614 49574 554058
rect 48954 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 49574 518614
rect 48954 518294 49574 518378
rect 48954 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 49574 518294
rect 48954 482614 49574 518058
rect 48954 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 49574 482614
rect 48954 482294 49574 482378
rect 48954 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 49574 482294
rect 48954 446614 49574 482058
rect 48954 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 49574 446614
rect 48954 446294 49574 446378
rect 48954 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 49574 446294
rect 48954 410614 49574 446058
rect 48954 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 49574 410614
rect 48954 410294 49574 410378
rect 48954 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 49574 410294
rect 48954 374614 49574 410058
rect 48954 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 49574 374614
rect 48954 374294 49574 374378
rect 48954 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 49574 374294
rect 48954 338614 49574 374058
rect 48954 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 49574 338614
rect 48954 338294 49574 338378
rect 48954 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 49574 338294
rect 48954 302614 49574 338058
rect 48954 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 49574 302614
rect 48954 302294 49574 302378
rect 48954 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 49574 302294
rect 48954 266614 49574 302058
rect 48954 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 49574 266614
rect 48954 266294 49574 266378
rect 48954 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 49574 266294
rect 48954 230614 49574 266058
rect 48954 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 49574 230614
rect 48954 230294 49574 230378
rect 48954 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 49574 230294
rect 48954 194614 49574 230058
rect 48954 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 49574 194614
rect 48954 194294 49574 194378
rect 48954 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 49574 194294
rect 48954 158614 49574 194058
rect 48954 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 49574 158614
rect 48954 158294 49574 158378
rect 48954 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 49574 158294
rect 48954 122614 49574 158058
rect 48954 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 49574 122614
rect 48954 122294 49574 122378
rect 48954 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 49574 122294
rect 48954 86614 49574 122058
rect 48954 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 49574 86614
rect 48954 86294 49574 86378
rect 48954 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 49574 86294
rect 48954 50614 49574 86058
rect 48954 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 49574 50614
rect 48954 50294 49574 50378
rect 48954 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 49574 50294
rect 48954 14614 49574 50058
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 30954 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 31574 -7066
rect 30954 -7386 31574 -7302
rect 30954 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 31574 -7386
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 14058
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 669454 56414 705242
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 59514 673174 60134 707162
rect 59514 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 60134 673174
rect 59514 672854 60134 672938
rect 59514 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 60134 672854
rect 59514 637174 60134 672618
rect 59514 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 60134 637174
rect 59514 636854 60134 636938
rect 59514 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 60134 636854
rect 59514 601174 60134 636618
rect 59514 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 60134 601174
rect 59514 600854 60134 600938
rect 59514 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 60134 600854
rect 59514 565174 60134 600618
rect 59514 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 60134 565174
rect 59514 564854 60134 564938
rect 59514 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 60134 564854
rect 59514 529174 60134 564618
rect 59514 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 60134 529174
rect 59514 528854 60134 528938
rect 59514 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 60134 528854
rect 59514 493174 60134 528618
rect 59514 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 60134 493174
rect 59514 492854 60134 492938
rect 59514 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 60134 492854
rect 59514 485308 60134 492618
rect 63234 676894 63854 709082
rect 63234 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 63854 676894
rect 63234 676574 63854 676658
rect 63234 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 63854 676574
rect 63234 640894 63854 676338
rect 63234 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 63854 640894
rect 63234 640574 63854 640658
rect 63234 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 63854 640574
rect 63234 604894 63854 640338
rect 63234 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 63854 604894
rect 63234 604574 63854 604658
rect 63234 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 63854 604574
rect 63234 568894 63854 604338
rect 63234 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 63854 568894
rect 63234 568574 63854 568658
rect 63234 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 63854 568574
rect 63234 532894 63854 568338
rect 63234 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 63854 532894
rect 63234 532574 63854 532658
rect 63234 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 63854 532574
rect 63234 496894 63854 532338
rect 63234 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 63854 496894
rect 63234 496574 63854 496658
rect 63234 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 63854 496574
rect 63234 485308 63854 496338
rect 66954 680614 67574 711002
rect 84954 710598 85574 711590
rect 84954 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 85574 710598
rect 84954 710278 85574 710362
rect 84954 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 85574 710278
rect 81234 708678 81854 709670
rect 81234 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 81854 708678
rect 81234 708358 81854 708442
rect 81234 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 81854 708358
rect 77514 706758 78134 707750
rect 77514 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 78134 706758
rect 77514 706438 78134 706522
rect 77514 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 78134 706438
rect 66954 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 67574 680614
rect 66954 680294 67574 680378
rect 66954 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 67574 680294
rect 66954 644614 67574 680058
rect 66954 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 67574 644614
rect 66954 644294 67574 644378
rect 66954 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 67574 644294
rect 66954 608614 67574 644058
rect 66954 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 67574 608614
rect 66954 608294 67574 608378
rect 66954 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 67574 608294
rect 66954 572614 67574 608058
rect 66954 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 67574 572614
rect 66954 572294 67574 572378
rect 66954 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 67574 572294
rect 66954 536614 67574 572058
rect 66954 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 67574 536614
rect 66954 536294 67574 536378
rect 66954 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 67574 536294
rect 66954 500614 67574 536058
rect 66954 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 67574 500614
rect 66954 500294 67574 500378
rect 66954 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 67574 500294
rect 66954 485308 67574 500058
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 543454 74414 578898
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 507454 74414 542898
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 485308 74414 506898
rect 77514 691174 78134 706202
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 655174 78134 690618
rect 77514 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 78134 655174
rect 77514 654854 78134 654938
rect 77514 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 78134 654854
rect 77514 619174 78134 654618
rect 77514 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 78134 619174
rect 77514 618854 78134 618938
rect 77514 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 78134 618854
rect 77514 583174 78134 618618
rect 77514 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 78134 583174
rect 77514 582854 78134 582938
rect 77514 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 78134 582854
rect 77514 547174 78134 582618
rect 77514 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 78134 547174
rect 77514 546854 78134 546938
rect 77514 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 78134 546854
rect 77514 511174 78134 546618
rect 77514 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 78134 511174
rect 77514 510854 78134 510938
rect 77514 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 78134 510854
rect 77514 485308 78134 510618
rect 81234 694894 81854 708122
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 658894 81854 694338
rect 81234 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 81854 658894
rect 81234 658574 81854 658658
rect 81234 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 81854 658574
rect 81234 622894 81854 658338
rect 81234 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 81854 622894
rect 81234 622574 81854 622658
rect 81234 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 81854 622574
rect 81234 586894 81854 622338
rect 81234 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 81854 586894
rect 81234 586574 81854 586658
rect 81234 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 81854 586574
rect 81234 550894 81854 586338
rect 81234 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 81854 550894
rect 81234 550574 81854 550658
rect 81234 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 81854 550574
rect 81234 514894 81854 550338
rect 81234 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 81854 514894
rect 81234 514574 81854 514658
rect 81234 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 81854 514574
rect 81234 485308 81854 514338
rect 84954 698614 85574 710042
rect 102954 711558 103574 711590
rect 102954 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 103574 711558
rect 102954 711238 103574 711322
rect 102954 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 103574 711238
rect 99234 709638 99854 709670
rect 99234 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 99854 709638
rect 99234 709318 99854 709402
rect 99234 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 99854 709318
rect 95514 707718 96134 707750
rect 95514 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 96134 707718
rect 95514 707398 96134 707482
rect 95514 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 96134 707398
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 662614 85574 698058
rect 84954 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 85574 662614
rect 84954 662294 85574 662378
rect 84954 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 85574 662294
rect 84954 626614 85574 662058
rect 84954 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 85574 626614
rect 84954 626294 85574 626378
rect 84954 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 85574 626294
rect 84954 590614 85574 626058
rect 84954 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 85574 590614
rect 84954 590294 85574 590378
rect 84954 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 85574 590294
rect 84954 554614 85574 590058
rect 84954 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 85574 554614
rect 84954 554294 85574 554378
rect 84954 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 85574 554294
rect 84954 518614 85574 554058
rect 84954 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 85574 518614
rect 84954 518294 85574 518378
rect 84954 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 85574 518294
rect 84954 485308 85574 518058
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 669454 92414 705242
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 561454 92414 596898
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 91794 525454 92414 560898
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 88747 503572 88813 503573
rect 88747 503508 88748 503572
rect 88812 503508 88813 503572
rect 88747 503507 88813 503508
rect 88750 498210 88810 503507
rect 88566 498150 88810 498210
rect 88566 491310 88626 498150
rect 88382 491250 88626 491310
rect 88382 483850 88442 491250
rect 89529 490380 89595 490381
rect 89529 490316 89530 490380
rect 89594 490316 89595 490380
rect 89529 490315 89595 490316
rect 91553 490380 91619 490381
rect 91553 490316 91554 490380
rect 91618 490316 91619 490380
rect 91553 490315 91619 490316
rect 89532 489970 89592 490315
rect 91556 489970 91616 490315
rect 89532 489910 89730 489970
rect 89670 484410 89730 489910
rect 91510 489910 91616 489970
rect 89670 484350 91202 484410
rect 91142 483850 91202 484350
rect 88382 483790 88764 483850
rect 88704 483202 88764 483790
rect 91016 483790 91202 483850
rect 91510 483850 91570 489910
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 91794 485308 92414 488898
rect 95514 673174 96134 707162
rect 95514 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 96134 673174
rect 95514 672854 96134 672938
rect 95514 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 96134 672854
rect 95514 637174 96134 672618
rect 95514 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 96134 637174
rect 95514 636854 96134 636938
rect 95514 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 96134 636854
rect 95514 601174 96134 636618
rect 95514 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 96134 601174
rect 95514 600854 96134 600938
rect 95514 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 96134 600854
rect 95514 565174 96134 600618
rect 95514 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 96134 565174
rect 95514 564854 96134 564938
rect 95514 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 96134 564854
rect 95514 529174 96134 564618
rect 95514 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 96134 529174
rect 95514 528854 96134 528938
rect 95514 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 96134 528854
rect 95514 493174 96134 528618
rect 99234 676894 99854 709082
rect 99234 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 99854 676894
rect 99234 676574 99854 676658
rect 99234 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 99854 676574
rect 99234 640894 99854 676338
rect 99234 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 99854 640894
rect 99234 640574 99854 640658
rect 99234 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 99854 640574
rect 99234 604894 99854 640338
rect 99234 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 99854 604894
rect 99234 604574 99854 604658
rect 99234 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 99854 604574
rect 99234 568894 99854 604338
rect 99234 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 99854 568894
rect 99234 568574 99854 568658
rect 99234 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 99854 568574
rect 99234 532894 99854 568338
rect 99234 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 99854 532894
rect 99234 532574 99854 532658
rect 99234 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 99854 532574
rect 96475 503572 96541 503573
rect 96475 503508 96476 503572
rect 96540 503508 96541 503572
rect 96475 503507 96541 503508
rect 98499 503572 98565 503573
rect 98499 503508 98500 503572
rect 98564 503508 98565 503572
rect 98499 503507 98565 503508
rect 95514 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 96134 493174
rect 95514 492854 96134 492938
rect 95514 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 96134 492854
rect 95514 485308 96134 492618
rect 96478 487170 96538 503507
rect 96478 487110 96722 487170
rect 96662 483850 96722 487110
rect 98502 483850 98562 503507
rect 99234 496894 99854 532338
rect 102954 680614 103574 711002
rect 120954 710598 121574 711590
rect 120954 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 121574 710598
rect 120954 710278 121574 710362
rect 120954 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 121574 710278
rect 117234 708678 117854 709670
rect 117234 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 117854 708678
rect 117234 708358 117854 708442
rect 117234 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 117854 708358
rect 113514 706758 114134 707750
rect 113514 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 114134 706758
rect 113514 706438 114134 706522
rect 113514 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 114134 706438
rect 102954 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 103574 680614
rect 102954 680294 103574 680378
rect 102954 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 103574 680294
rect 102954 644614 103574 680058
rect 102954 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 103574 644614
rect 102954 644294 103574 644378
rect 102954 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 103574 644294
rect 102954 608614 103574 644058
rect 102954 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 103574 608614
rect 102954 608294 103574 608378
rect 102954 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 103574 608294
rect 102954 572614 103574 608058
rect 102954 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 103574 572614
rect 102954 572294 103574 572378
rect 102954 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 103574 572294
rect 102954 536614 103574 572058
rect 102954 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 103574 536614
rect 102954 536294 103574 536378
rect 102954 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 103574 536294
rect 101259 503572 101325 503573
rect 101259 503508 101260 503572
rect 101324 503508 101325 503572
rect 101259 503507 101325 503508
rect 99234 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 99854 496894
rect 99234 496574 99854 496658
rect 99234 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 99854 496574
rect 99234 485308 99854 496338
rect 101262 483850 101322 503507
rect 102954 500614 103574 536058
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 103835 503572 103901 503573
rect 103835 503508 103836 503572
rect 103900 503508 103901 503572
rect 103835 503507 103901 503508
rect 106043 503572 106109 503573
rect 106043 503508 106044 503572
rect 106108 503508 106109 503572
rect 106043 503507 106109 503508
rect 102954 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 103574 500614
rect 102954 500294 103574 500378
rect 102954 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 103574 500294
rect 102954 485308 103574 500058
rect 103838 498210 103898 503507
rect 103654 498150 103898 498210
rect 103654 487170 103714 498150
rect 103654 487110 103898 487170
rect 103838 483850 103898 487110
rect 91510 483790 93524 483850
rect 91016 483202 91076 483790
rect 93464 483202 93524 483790
rect 96184 483790 96722 483850
rect 98496 483790 98562 483850
rect 101080 483790 101322 483850
rect 103528 483790 103898 483850
rect 106046 483850 106106 503507
rect 108297 491060 108363 491061
rect 108297 490996 108298 491060
rect 108362 490996 108363 491060
rect 108297 490995 108363 490996
rect 108300 490650 108360 490995
rect 108254 490590 108360 490650
rect 108254 484258 108314 490590
rect 109794 485308 110414 506898
rect 113514 691174 114134 706202
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 655174 114134 690618
rect 113514 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 114134 655174
rect 113514 654854 114134 654938
rect 113514 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 114134 654854
rect 113514 619174 114134 654618
rect 113514 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 114134 619174
rect 113514 618854 114134 618938
rect 113514 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 114134 618854
rect 113514 583174 114134 618618
rect 113514 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 114134 583174
rect 113514 582854 114134 582938
rect 113514 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 114134 582854
rect 113514 547174 114134 582618
rect 113514 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 114134 547174
rect 113514 546854 114134 546938
rect 113514 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 114134 546854
rect 113514 511174 114134 546618
rect 113514 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 114134 511174
rect 113514 510854 114134 510938
rect 113514 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 114134 510854
rect 111977 488340 112043 488341
rect 111977 488276 111978 488340
rect 112042 488276 112043 488340
rect 111977 488275 112043 488276
rect 111980 487930 112040 488275
rect 111980 487870 112178 487930
rect 112118 484410 112178 487870
rect 113514 485308 114134 510618
rect 117234 694894 117854 708122
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 658894 117854 694338
rect 117234 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 117854 658894
rect 117234 658574 117854 658658
rect 117234 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 117854 658574
rect 117234 622894 117854 658338
rect 117234 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 117854 622894
rect 117234 622574 117854 622658
rect 117234 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 117854 622574
rect 117234 586894 117854 622338
rect 117234 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 117854 586894
rect 117234 586574 117854 586658
rect 117234 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 117854 586574
rect 117234 550894 117854 586338
rect 117234 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 117854 550894
rect 117234 550574 117854 550658
rect 117234 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 117854 550574
rect 117234 514894 117854 550338
rect 117234 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 117854 514894
rect 117234 514574 117854 514658
rect 117234 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 117854 514574
rect 116163 503708 116229 503709
rect 116163 503644 116164 503708
rect 116228 503644 116229 503708
rect 116163 503643 116229 503644
rect 116166 485790 116226 503643
rect 116166 485730 116410 485790
rect 112118 484350 113650 484410
rect 108254 484198 108682 484258
rect 106046 483790 106172 483850
rect 96184 483202 96244 483790
rect 98496 483202 98556 483790
rect 101080 483202 101140 483790
rect 103528 483202 103588 483790
rect 106112 483202 106172 483790
rect 108622 483232 108682 484198
rect 113590 483850 113650 484350
rect 116350 483850 116410 485730
rect 117234 485308 117854 514338
rect 120954 698614 121574 710042
rect 138954 711558 139574 711590
rect 138954 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 139574 711558
rect 138954 711238 139574 711322
rect 138954 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 139574 711238
rect 135234 709638 135854 709670
rect 135234 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 135854 709638
rect 135234 709318 135854 709402
rect 135234 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 135854 709318
rect 131514 707718 132134 707750
rect 131514 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 132134 707718
rect 131514 707398 132134 707482
rect 131514 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 132134 707398
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 662614 121574 698058
rect 120954 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 121574 662614
rect 120954 662294 121574 662378
rect 120954 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 121574 662294
rect 120954 626614 121574 662058
rect 120954 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 121574 626614
rect 120954 626294 121574 626378
rect 120954 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 121574 626294
rect 120954 590614 121574 626058
rect 120954 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 121574 590614
rect 120954 590294 121574 590378
rect 120954 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 121574 590294
rect 120954 554614 121574 590058
rect 120954 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 121574 554614
rect 120954 554294 121574 554378
rect 120954 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 121574 554294
rect 120954 518614 121574 554058
rect 120954 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 121574 518614
rect 120954 518294 121574 518378
rect 120954 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 121574 518294
rect 118187 503572 118253 503573
rect 118187 503508 118188 503572
rect 118252 503508 118253 503572
rect 118187 503507 118253 503508
rect 118190 491310 118250 503507
rect 118006 491250 118250 491310
rect 118558 495350 120826 495410
rect 118006 487170 118066 491250
rect 118006 487110 118250 487170
rect 108590 483172 108682 483232
rect 111144 483790 111442 483850
rect 113590 483790 113652 483850
rect 111144 483202 111204 483790
rect 111382 483717 111442 483790
rect 111379 483716 111445 483717
rect 111379 483652 111380 483716
rect 111444 483652 111445 483716
rect 111379 483651 111445 483652
rect 113592 483202 113652 483790
rect 116176 483790 116410 483850
rect 118190 483850 118250 487110
rect 118558 485213 118618 495350
rect 118509 485212 118618 485213
rect 118509 485148 118510 485212
rect 118574 485150 118618 485212
rect 118574 485148 118575 485150
rect 118509 485147 118575 485148
rect 120766 483850 120826 495350
rect 120954 485308 121574 518058
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 127794 669454 128414 705242
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 123523 503572 123589 503573
rect 123523 503508 123524 503572
rect 123588 503508 123589 503572
rect 123523 503507 123589 503508
rect 123891 503572 123957 503573
rect 123891 503508 123892 503572
rect 123956 503508 123957 503572
rect 123891 503507 123957 503508
rect 123526 487170 123586 503507
rect 123526 487110 123770 487170
rect 123710 483850 123770 487110
rect 123894 484410 123954 503507
rect 127794 489454 128414 524898
rect 131514 673174 132134 707162
rect 131514 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 132134 673174
rect 131514 672854 132134 672938
rect 131514 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 132134 672854
rect 131514 637174 132134 672618
rect 131514 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 132134 637174
rect 131514 636854 132134 636938
rect 131514 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 132134 636854
rect 131514 601174 132134 636618
rect 131514 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 132134 601174
rect 131514 600854 132134 600938
rect 131514 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 132134 600854
rect 131514 565174 132134 600618
rect 131514 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 132134 565174
rect 131514 564854 132134 564938
rect 131514 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 132134 564854
rect 131514 529174 132134 564618
rect 131514 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 132134 529174
rect 131514 528854 132134 528938
rect 131514 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 132134 528854
rect 128675 504388 128741 504389
rect 128675 504324 128676 504388
rect 128740 504324 128741 504388
rect 128675 504323 128741 504324
rect 128678 495450 128738 504323
rect 129779 503572 129845 503573
rect 129779 503508 129780 503572
rect 129844 503508 129845 503572
rect 129779 503507 129845 503508
rect 129782 498210 129842 503507
rect 129782 498150 130026 498210
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 127794 485308 128414 488898
rect 128494 495390 128738 495450
rect 123894 484350 126162 484410
rect 118190 483790 118548 483850
rect 120766 483790 120996 483850
rect 116176 483202 116236 483790
rect 118488 483202 118548 483790
rect 120936 483202 120996 483790
rect 123656 483790 123770 483850
rect 126102 483850 126162 484350
rect 128494 483850 128554 495390
rect 129966 483850 130026 498150
rect 131514 493174 132134 528618
rect 135234 676894 135854 709082
rect 135234 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 135854 676894
rect 135234 676574 135854 676658
rect 135234 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 135854 676574
rect 135234 640894 135854 676338
rect 135234 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 135854 640894
rect 135234 640574 135854 640658
rect 135234 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 135854 640574
rect 135234 604894 135854 640338
rect 135234 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 135854 604894
rect 135234 604574 135854 604658
rect 135234 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 135854 604574
rect 135234 568894 135854 604338
rect 135234 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 135854 568894
rect 135234 568574 135854 568658
rect 135234 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 135854 568574
rect 135234 532894 135854 568338
rect 135234 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 135854 532894
rect 135234 532574 135854 532658
rect 135234 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 135854 532574
rect 134931 503708 134997 503709
rect 134931 503644 134932 503708
rect 134996 503644 134997 503708
rect 134931 503643 134997 503644
rect 131514 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 132134 493174
rect 131514 492854 132134 492938
rect 131514 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 132134 492854
rect 131514 485308 132134 492618
rect 133462 491950 133660 492010
rect 133462 483986 133522 491950
rect 133600 491877 133660 491950
rect 133597 491876 133663 491877
rect 133597 491812 133598 491876
rect 133662 491812 133663 491876
rect 133597 491811 133663 491812
rect 134934 491310 134994 503643
rect 134750 491250 134994 491310
rect 135234 496894 135854 532338
rect 135234 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 135854 496894
rect 135234 496574 135854 496658
rect 135234 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 135854 496574
rect 134750 487170 134810 491250
rect 134750 487110 134994 487170
rect 134934 483986 134994 487110
rect 135234 485308 135854 496338
rect 138954 680614 139574 711002
rect 156954 710598 157574 711590
rect 156954 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 157574 710598
rect 156954 710278 157574 710362
rect 156954 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 157574 710278
rect 153234 708678 153854 709670
rect 153234 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 153854 708678
rect 153234 708358 153854 708442
rect 153234 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 153854 708358
rect 149514 706758 150134 707750
rect 149514 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 150134 706758
rect 149514 706438 150134 706522
rect 149514 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 150134 706438
rect 138954 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 139574 680614
rect 138954 680294 139574 680378
rect 138954 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 139574 680294
rect 138954 644614 139574 680058
rect 138954 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 139574 644614
rect 138954 644294 139574 644378
rect 138954 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 139574 644294
rect 138954 608614 139574 644058
rect 138954 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 139574 608614
rect 138954 608294 139574 608378
rect 138954 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 139574 608294
rect 138954 572614 139574 608058
rect 138954 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 139574 572614
rect 138954 572294 139574 572378
rect 138954 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 139574 572294
rect 138954 536614 139574 572058
rect 138954 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 139574 536614
rect 138954 536294 139574 536378
rect 138954 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 139574 536294
rect 138954 500614 139574 536058
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 143211 503572 143277 503573
rect 143211 503508 143212 503572
rect 143276 503508 143277 503572
rect 143211 503507 143277 503508
rect 144867 503572 144933 503573
rect 144867 503508 144868 503572
rect 144932 503508 144933 503572
rect 144867 503507 144933 503508
rect 138954 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 139574 500614
rect 138954 500294 139574 500378
rect 138954 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 139574 500294
rect 138954 485308 139574 500058
rect 143214 492690 143274 503507
rect 144870 502350 144930 503507
rect 143950 502290 144930 502350
rect 143950 492690 144010 502290
rect 141006 492630 143274 492690
rect 143582 492630 144010 492690
rect 141006 491310 141066 492630
rect 143582 492010 143642 492630
rect 139718 491250 141066 491310
rect 141190 491950 143642 492010
rect 133462 483926 133660 483986
rect 134934 483926 135914 483986
rect 133600 483850 133660 483926
rect 126102 483790 126164 483850
rect 128494 483790 128612 483850
rect 129966 483790 131060 483850
rect 123656 483202 123716 483790
rect 126104 483202 126164 483790
rect 128552 483202 128612 483790
rect 131000 483202 131060 483790
rect 133584 483790 133660 483850
rect 135854 483850 135914 483926
rect 139718 483850 139778 491250
rect 141190 483850 141250 491950
rect 145794 485308 146414 506898
rect 149514 691174 150134 706202
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 655174 150134 690618
rect 149514 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 150134 655174
rect 149514 654854 150134 654938
rect 149514 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 150134 654854
rect 149514 619174 150134 654618
rect 149514 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 150134 619174
rect 149514 618854 150134 618938
rect 149514 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 150134 618854
rect 149514 583174 150134 618618
rect 149514 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 150134 583174
rect 149514 582854 150134 582938
rect 149514 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 150134 582854
rect 149514 547174 150134 582618
rect 149514 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 150134 547174
rect 149514 546854 150134 546938
rect 149514 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 150134 546854
rect 149514 511174 150134 546618
rect 149514 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 150134 511174
rect 149514 510854 150134 510938
rect 149514 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 150134 510854
rect 146523 503572 146589 503573
rect 146523 503508 146524 503572
rect 146588 503508 146589 503572
rect 146523 503507 146589 503508
rect 148363 503572 148429 503573
rect 148363 503508 148364 503572
rect 148428 503508 148429 503572
rect 148363 503507 148429 503508
rect 143027 484124 143093 484125
rect 143027 484060 143028 484124
rect 143092 484060 143093 484124
rect 143027 484059 143093 484060
rect 135854 483790 135956 483850
rect 133584 483202 133644 483790
rect 135896 483202 135956 483790
rect 138616 483790 139778 483850
rect 141064 483790 141250 483850
rect 143030 483850 143090 484059
rect 146526 483850 146586 503507
rect 148366 491310 148426 503507
rect 148366 491250 148610 491310
rect 148550 484410 148610 491250
rect 149514 485308 150134 510618
rect 153234 694894 153854 708122
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 658894 153854 694338
rect 153234 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 153854 658894
rect 153234 658574 153854 658658
rect 153234 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 153854 658574
rect 153234 622894 153854 658338
rect 153234 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 153854 622894
rect 153234 622574 153854 622658
rect 153234 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 153854 622574
rect 153234 586894 153854 622338
rect 153234 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 153854 586894
rect 153234 586574 153854 586658
rect 153234 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 153854 586574
rect 153234 550894 153854 586338
rect 153234 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 153854 550894
rect 153234 550574 153854 550658
rect 153234 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 153854 550574
rect 153234 514894 153854 550338
rect 153234 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 153854 514894
rect 153234 514574 153854 514658
rect 153234 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 153854 514574
rect 151123 503708 151189 503709
rect 151123 503644 151124 503708
rect 151188 503644 151189 503708
rect 151123 503643 151189 503644
rect 151126 495450 151186 503643
rect 151080 495410 151186 495450
rect 150942 495390 151186 495410
rect 150942 495350 151140 495390
rect 150942 491310 151002 495350
rect 153009 491740 153075 491741
rect 153009 491676 153010 491740
rect 153074 491676 153075 491740
rect 153009 491675 153075 491676
rect 153012 491330 153072 491675
rect 150758 491250 151002 491310
rect 152966 491270 153072 491330
rect 150758 489290 150818 491250
rect 150758 489230 151002 489290
rect 143030 483790 143572 483850
rect 138616 483202 138676 483790
rect 141064 483202 141124 483790
rect 143512 483202 143572 483790
rect 145960 483790 146586 483850
rect 148366 484350 148610 484410
rect 148366 483850 148426 484350
rect 150942 483850 151002 489230
rect 152966 483850 153026 491270
rect 153234 485308 153854 514338
rect 156954 698614 157574 710042
rect 174954 711558 175574 711590
rect 174954 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 175574 711558
rect 174954 711238 175574 711322
rect 174954 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 175574 711238
rect 171234 709638 171854 709670
rect 171234 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 171854 709638
rect 171234 709318 171854 709402
rect 171234 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 171854 709318
rect 167514 707718 168134 707750
rect 167514 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 168134 707718
rect 167514 707398 168134 707482
rect 167514 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 168134 707398
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 662614 157574 698058
rect 156954 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 157574 662614
rect 156954 662294 157574 662378
rect 156954 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 157574 662294
rect 156954 626614 157574 662058
rect 156954 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 157574 626614
rect 156954 626294 157574 626378
rect 156954 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 157574 626294
rect 156954 590614 157574 626058
rect 156954 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 157574 590614
rect 156954 590294 157574 590378
rect 156954 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 157574 590294
rect 156954 554614 157574 590058
rect 156954 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 157574 554614
rect 156954 554294 157574 554378
rect 156954 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 157574 554294
rect 156954 518614 157574 554058
rect 156954 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 157574 518614
rect 156954 518294 157574 518378
rect 156954 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 157574 518294
rect 155907 503572 155973 503573
rect 155907 503508 155908 503572
rect 155972 503508 155973 503572
rect 155907 503507 155973 503508
rect 155910 483850 155970 503507
rect 156954 485308 157574 518058
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 669454 164414 705242
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 158667 503572 158733 503573
rect 158667 503508 158668 503572
rect 158732 503508 158733 503572
rect 158667 503507 158733 503508
rect 160139 503572 160205 503573
rect 160139 503508 160140 503572
rect 160204 503508 160205 503572
rect 160139 503507 160205 503508
rect 163451 503572 163517 503573
rect 163451 503508 163452 503572
rect 163516 503508 163517 503572
rect 163451 503507 163517 503508
rect 158670 489930 158730 503507
rect 160142 495410 160202 503507
rect 160142 495350 160386 495410
rect 160326 491330 160386 495350
rect 160326 491270 160754 491330
rect 158486 489870 158730 489930
rect 158486 485790 158546 489870
rect 158486 485730 158730 485790
rect 158670 483850 158730 485730
rect 148366 483790 148468 483850
rect 150942 483790 151052 483850
rect 152966 483790 153636 483850
rect 155910 483790 156084 483850
rect 145960 483202 146020 483790
rect 148408 483202 148468 483790
rect 150992 483202 151052 483790
rect 153576 483202 153636 483790
rect 156024 483202 156084 483790
rect 158472 483790 158730 483850
rect 160694 483850 160754 491270
rect 163454 483850 163514 503507
rect 163794 489454 164414 524898
rect 167514 673174 168134 707162
rect 167514 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 168134 673174
rect 167514 672854 168134 672938
rect 167514 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 168134 672854
rect 167514 637174 168134 672618
rect 167514 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 168134 637174
rect 167514 636854 168134 636938
rect 167514 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 168134 636854
rect 167514 601174 168134 636618
rect 167514 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 168134 601174
rect 167514 600854 168134 600938
rect 167514 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 168134 600854
rect 167514 565174 168134 600618
rect 167514 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 168134 565174
rect 167514 564854 168134 564938
rect 167514 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 168134 564854
rect 167514 529174 168134 564618
rect 167514 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 168134 529174
rect 167514 528854 168134 528938
rect 167514 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 168134 528854
rect 165659 503572 165725 503573
rect 165659 503508 165660 503572
rect 165724 503508 165725 503572
rect 165659 503507 165725 503508
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 485308 164414 488898
rect 165662 488550 165722 503507
rect 167514 493174 168134 528618
rect 167514 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 168134 493174
rect 167514 492854 168134 492938
rect 167514 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 168134 492854
rect 165662 488490 166090 488550
rect 166030 487170 166090 488490
rect 166030 487110 166274 487170
rect 166214 483850 166274 487110
rect 167514 485308 168134 492618
rect 171234 676894 171854 709082
rect 171234 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 171854 676894
rect 171234 676574 171854 676658
rect 171234 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 171854 676574
rect 171234 640894 171854 676338
rect 171234 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 171854 640894
rect 171234 640574 171854 640658
rect 171234 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 171854 640574
rect 171234 604894 171854 640338
rect 171234 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 171854 604894
rect 171234 604574 171854 604658
rect 171234 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 171854 604574
rect 171234 568894 171854 604338
rect 171234 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 171854 568894
rect 171234 568574 171854 568658
rect 171234 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 171854 568574
rect 171234 532894 171854 568338
rect 171234 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 171854 532894
rect 171234 532574 171854 532658
rect 171234 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 171854 532574
rect 171234 496894 171854 532338
rect 171234 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 171854 496894
rect 171234 496574 171854 496658
rect 171234 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 171854 496574
rect 171234 485308 171854 496338
rect 174954 680614 175574 711002
rect 192954 710598 193574 711590
rect 192954 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 193574 710598
rect 192954 710278 193574 710362
rect 192954 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 193574 710278
rect 189234 708678 189854 709670
rect 189234 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 189854 708678
rect 189234 708358 189854 708442
rect 189234 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 189854 708358
rect 185514 706758 186134 707750
rect 185514 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 186134 706758
rect 185514 706438 186134 706522
rect 185514 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 186134 706438
rect 174954 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 175574 680614
rect 174954 680294 175574 680378
rect 174954 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 175574 680294
rect 174954 644614 175574 680058
rect 174954 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 175574 644614
rect 174954 644294 175574 644378
rect 174954 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 175574 644294
rect 174954 608614 175574 644058
rect 174954 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 175574 608614
rect 174954 608294 175574 608378
rect 174954 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 175574 608294
rect 174954 572614 175574 608058
rect 174954 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 175574 572614
rect 174954 572294 175574 572378
rect 174954 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 175574 572294
rect 174954 536614 175574 572058
rect 174954 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 175574 536614
rect 174954 536294 175574 536378
rect 174954 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 175574 536294
rect 174954 500614 175574 536058
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 178539 503708 178605 503709
rect 178539 503644 178540 503708
rect 178604 503644 178605 503708
rect 178539 503643 178605 503644
rect 174954 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 175574 500614
rect 174954 500294 175574 500378
rect 174954 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 175574 500294
rect 174954 485308 175574 500058
rect 178542 491310 178602 503643
rect 178358 491250 178602 491310
rect 178358 487170 178418 491250
rect 178358 487110 178602 487170
rect 178542 483850 178602 487110
rect 181794 485308 182414 506898
rect 185514 691174 186134 706202
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 655174 186134 690618
rect 185514 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 186134 655174
rect 185514 654854 186134 654938
rect 185514 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 186134 654854
rect 185514 619174 186134 654618
rect 185514 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 186134 619174
rect 185514 618854 186134 618938
rect 185514 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 186134 618854
rect 185514 583174 186134 618618
rect 185514 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 186134 583174
rect 185514 582854 186134 582938
rect 185514 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 186134 582854
rect 185514 547174 186134 582618
rect 185514 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 186134 547174
rect 185514 546854 186134 546938
rect 185514 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 186134 546854
rect 185514 511174 186134 546618
rect 185514 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 186134 511174
rect 185514 510854 186134 510938
rect 185514 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 186134 510854
rect 185514 485308 186134 510618
rect 189234 694894 189854 708122
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 658894 189854 694338
rect 189234 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 189854 658894
rect 189234 658574 189854 658658
rect 189234 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 189854 658574
rect 189234 622894 189854 658338
rect 189234 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 189854 622894
rect 189234 622574 189854 622658
rect 189234 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 189854 622574
rect 189234 586894 189854 622338
rect 189234 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 189854 586894
rect 189234 586574 189854 586658
rect 189234 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 189854 586574
rect 189234 550894 189854 586338
rect 189234 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 189854 550894
rect 189234 550574 189854 550658
rect 189234 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 189854 550574
rect 189234 514894 189854 550338
rect 189234 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 189854 514894
rect 189234 514574 189854 514658
rect 189234 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 189854 514574
rect 189234 485308 189854 514338
rect 192954 698614 193574 710042
rect 210954 711558 211574 711590
rect 210954 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 211574 711558
rect 210954 711238 211574 711322
rect 210954 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 211574 711238
rect 207234 709638 207854 709670
rect 207234 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 207854 709638
rect 207234 709318 207854 709402
rect 207234 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 207854 709318
rect 203514 707718 204134 707750
rect 203514 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 204134 707718
rect 203514 707398 204134 707482
rect 203514 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 204134 707398
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 662614 193574 698058
rect 192954 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 193574 662614
rect 192954 662294 193574 662378
rect 192954 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 193574 662294
rect 192954 626614 193574 662058
rect 192954 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 193574 626614
rect 192954 626294 193574 626378
rect 192954 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 193574 626294
rect 192954 590614 193574 626058
rect 192954 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 193574 590614
rect 192954 590294 193574 590378
rect 192954 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 193574 590294
rect 192954 554614 193574 590058
rect 192954 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 193574 554614
rect 192954 554294 193574 554378
rect 192954 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 193574 554294
rect 192954 518614 193574 554058
rect 192954 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 193574 518614
rect 192954 518294 193574 518378
rect 192954 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 193574 518294
rect 192954 485308 193574 518058
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 669454 200414 705242
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 525454 200414 560898
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 489454 200414 524898
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 196755 486300 196821 486301
rect 196755 486236 196756 486300
rect 196820 486236 196821 486300
rect 196755 486235 196821 486236
rect 180195 484124 180261 484125
rect 180195 484122 180196 484124
rect 179830 484062 180196 484122
rect 179830 483850 179890 484062
rect 180195 484060 180196 484062
rect 180260 484060 180261 484124
rect 180195 484059 180261 484060
rect 196758 483850 196818 486235
rect 160694 483790 161116 483850
rect 158472 483202 158532 483790
rect 161056 483202 161116 483790
rect 163368 483790 163514 483850
rect 166088 483790 166274 483850
rect 178464 483790 178602 483850
rect 179688 483790 179890 483850
rect 190840 483790 196818 483850
rect 163368 483202 163428 483790
rect 166088 483202 166148 483790
rect 178464 483202 178524 483790
rect 179688 483202 179748 483790
rect 190840 483202 190900 483790
rect 60952 471454 61300 471486
rect 60952 471218 61008 471454
rect 61244 471218 61300 471454
rect 60952 471134 61300 471218
rect 60952 470898 61008 471134
rect 61244 470898 61300 471134
rect 60952 470866 61300 470898
rect 195320 471454 195668 471486
rect 195320 471218 195376 471454
rect 195612 471218 195668 471454
rect 195320 471134 195668 471218
rect 195320 470898 195376 471134
rect 195612 470898 195668 471134
rect 195320 470866 195668 470898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 60272 453454 60620 453486
rect 60272 453218 60328 453454
rect 60564 453218 60620 453454
rect 60272 453134 60620 453218
rect 60272 452898 60328 453134
rect 60564 452898 60620 453134
rect 60272 452866 60620 452898
rect 196000 453454 196348 453486
rect 196000 453218 196056 453454
rect 196292 453218 196348 453454
rect 196000 453134 196348 453218
rect 196000 452898 196056 453134
rect 196292 452898 196348 453134
rect 196000 452866 196348 452898
rect 199794 453454 200414 488898
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 60952 435454 61300 435486
rect 60952 435218 61008 435454
rect 61244 435218 61300 435454
rect 60952 435134 61300 435218
rect 60952 434898 61008 435134
rect 61244 434898 61300 435134
rect 60952 434866 61300 434898
rect 195320 435454 195668 435486
rect 195320 435218 195376 435454
rect 195612 435218 195668 435454
rect 195320 435134 195668 435218
rect 195320 434898 195376 435134
rect 195612 434898 195668 435134
rect 195320 434866 195668 434898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 60272 417454 60620 417486
rect 60272 417218 60328 417454
rect 60564 417218 60620 417454
rect 60272 417134 60620 417218
rect 60272 416898 60328 417134
rect 60564 416898 60620 417134
rect 60272 416866 60620 416898
rect 196000 417454 196348 417486
rect 196000 417218 196056 417454
rect 196292 417218 196348 417454
rect 196000 417134 196348 417218
rect 196000 416898 196056 417134
rect 196292 416898 196348 417134
rect 196000 416866 196348 416898
rect 199794 417454 200414 452898
rect 199794 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 200414 417454
rect 199794 417134 200414 417218
rect 199794 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 200414 417134
rect 76056 399530 76116 400106
rect 76054 399470 76116 399530
rect 77144 399530 77204 400106
rect 78232 399530 78292 400106
rect 79592 399530 79652 400106
rect 77144 399470 77218 399530
rect 78232 399470 78322 399530
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 59514 385174 60134 398000
rect 59514 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 60134 385174
rect 59514 384854 60134 384938
rect 59514 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 60134 384854
rect 59514 349174 60134 384618
rect 59514 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 60134 349174
rect 59514 348854 60134 348938
rect 59514 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 60134 348854
rect 59514 313174 60134 348618
rect 59514 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 60134 313174
rect 59514 312854 60134 312938
rect 59514 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 60134 312854
rect 59514 277174 60134 312618
rect 59514 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 60134 277174
rect 59514 276854 60134 276938
rect 59514 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 60134 276854
rect 59514 241174 60134 276618
rect 59514 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 60134 241174
rect 59514 240854 60134 240938
rect 59514 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 60134 240854
rect 59514 228675 60134 240618
rect 63234 388894 63854 398000
rect 63234 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 63854 388894
rect 63234 388574 63854 388658
rect 63234 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 63854 388574
rect 63234 352894 63854 388338
rect 63234 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 63854 352894
rect 63234 352574 63854 352658
rect 63234 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 63854 352574
rect 63234 316894 63854 352338
rect 63234 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 63854 316894
rect 63234 316574 63854 316658
rect 63234 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 63854 316574
rect 63234 280894 63854 316338
rect 63234 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 63854 280894
rect 63234 280574 63854 280658
rect 63234 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 63854 280574
rect 63234 244894 63854 280338
rect 63234 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 63854 244894
rect 63234 244574 63854 244658
rect 63234 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 63854 244574
rect 63234 228675 63854 244338
rect 66954 392614 67574 398000
rect 66954 392378 66986 392614
rect 67222 392378 67306 392614
rect 67542 392378 67574 392614
rect 66954 392294 67574 392378
rect 66954 392058 66986 392294
rect 67222 392058 67306 392294
rect 67542 392058 67574 392294
rect 66954 356614 67574 392058
rect 66954 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 67574 356614
rect 66954 356294 67574 356378
rect 66954 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 67574 356294
rect 66954 320614 67574 356058
rect 66954 320378 66986 320614
rect 67222 320378 67306 320614
rect 67542 320378 67574 320614
rect 66954 320294 67574 320378
rect 66954 320058 66986 320294
rect 67222 320058 67306 320294
rect 67542 320058 67574 320294
rect 66954 284614 67574 320058
rect 66954 284378 66986 284614
rect 67222 284378 67306 284614
rect 67542 284378 67574 284614
rect 66954 284294 67574 284378
rect 66954 284058 66986 284294
rect 67222 284058 67306 284294
rect 67542 284058 67574 284294
rect 66954 248614 67574 284058
rect 66954 248378 66986 248614
rect 67222 248378 67306 248614
rect 67542 248378 67574 248614
rect 66954 248294 67574 248378
rect 66954 248058 66986 248294
rect 67222 248058 67306 248294
rect 67542 248058 67574 248294
rect 66954 228675 67574 248058
rect 73794 363454 74414 398000
rect 76054 396677 76114 399470
rect 77158 396813 77218 399470
rect 77155 396812 77221 396813
rect 77155 396748 77156 396812
rect 77220 396748 77221 396812
rect 77155 396747 77221 396748
rect 76051 396676 76117 396677
rect 76051 396612 76052 396676
rect 76116 396612 76117 396676
rect 76051 396611 76117 396612
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 327454 74414 362898
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 73794 291454 74414 326898
rect 73794 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 74414 291454
rect 73794 291134 74414 291218
rect 73794 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 74414 291134
rect 73794 255454 74414 290898
rect 73794 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 74414 255454
rect 73794 255134 74414 255218
rect 73794 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 74414 255134
rect 73794 228675 74414 254898
rect 77514 367174 78134 398000
rect 78262 397357 78322 399470
rect 79550 399470 79652 399530
rect 80544 399530 80604 400106
rect 81768 399530 81828 400106
rect 83128 399530 83188 400106
rect 84216 399530 84276 400106
rect 85440 399530 85500 400106
rect 80544 399470 80714 399530
rect 81768 399470 82002 399530
rect 83128 399470 83290 399530
rect 84216 399470 84394 399530
rect 78259 397356 78325 397357
rect 78259 397292 78260 397356
rect 78324 397292 78325 397356
rect 78259 397291 78325 397292
rect 79550 396813 79610 399470
rect 80654 397357 80714 399470
rect 80651 397356 80717 397357
rect 80651 397292 80652 397356
rect 80716 397292 80717 397356
rect 80651 397291 80717 397292
rect 79547 396812 79613 396813
rect 79547 396748 79548 396812
rect 79612 396748 79613 396812
rect 79547 396747 79613 396748
rect 77514 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 78134 367174
rect 77514 366854 78134 366938
rect 77514 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 78134 366854
rect 77514 331174 78134 366618
rect 77514 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 78134 331174
rect 77514 330854 78134 330938
rect 77514 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 78134 330854
rect 77514 295174 78134 330618
rect 77514 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 78134 295174
rect 77514 294854 78134 294938
rect 77514 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 78134 294854
rect 77514 259174 78134 294618
rect 77514 258938 77546 259174
rect 77782 258938 77866 259174
rect 78102 258938 78134 259174
rect 77514 258854 78134 258938
rect 77514 258618 77546 258854
rect 77782 258618 77866 258854
rect 78102 258618 78134 258854
rect 77514 228675 78134 258618
rect 81234 370894 81854 398000
rect 81942 397357 82002 399470
rect 83230 397357 83290 399470
rect 84334 397357 84394 399470
rect 85438 399470 85500 399530
rect 86528 399530 86588 400106
rect 87616 399530 87676 400106
rect 88296 399530 88356 400106
rect 88704 399530 88764 400106
rect 90064 399530 90124 400106
rect 86528 399470 86602 399530
rect 87616 399470 87706 399530
rect 88296 399470 88442 399530
rect 88704 399470 88810 399530
rect 85438 398173 85498 399470
rect 85435 398172 85501 398173
rect 85435 398108 85436 398172
rect 85500 398108 85501 398172
rect 85435 398107 85501 398108
rect 81939 397356 82005 397357
rect 81939 397292 81940 397356
rect 82004 397292 82005 397356
rect 81939 397291 82005 397292
rect 83227 397356 83293 397357
rect 83227 397292 83228 397356
rect 83292 397292 83293 397356
rect 83227 397291 83293 397292
rect 84331 397356 84397 397357
rect 84331 397292 84332 397356
rect 84396 397292 84397 397356
rect 84331 397291 84397 397292
rect 81234 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 81854 370894
rect 81234 370574 81854 370658
rect 81234 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 81854 370574
rect 81234 334894 81854 370338
rect 81234 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 81854 334894
rect 81234 334574 81854 334658
rect 81234 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 81854 334574
rect 81234 298894 81854 334338
rect 81234 298658 81266 298894
rect 81502 298658 81586 298894
rect 81822 298658 81854 298894
rect 81234 298574 81854 298658
rect 81234 298338 81266 298574
rect 81502 298338 81586 298574
rect 81822 298338 81854 298574
rect 81234 262894 81854 298338
rect 81234 262658 81266 262894
rect 81502 262658 81586 262894
rect 81822 262658 81854 262894
rect 81234 262574 81854 262658
rect 81234 262338 81266 262574
rect 81502 262338 81586 262574
rect 81822 262338 81854 262574
rect 81234 228675 81854 262338
rect 84954 374614 85574 398000
rect 86542 396813 86602 399470
rect 87646 397357 87706 399470
rect 87643 397356 87709 397357
rect 87643 397292 87644 397356
rect 87708 397292 87709 397356
rect 87643 397291 87709 397292
rect 88382 396813 88442 399470
rect 88750 397357 88810 399470
rect 90038 399470 90124 399530
rect 90744 399530 90804 400106
rect 91288 399530 91348 400106
rect 92376 399530 92436 400106
rect 93464 399530 93524 400106
rect 90744 399470 90834 399530
rect 91288 399470 91386 399530
rect 92376 399470 92490 399530
rect 90038 397357 90098 399470
rect 88747 397356 88813 397357
rect 88747 397292 88748 397356
rect 88812 397292 88813 397356
rect 88747 397291 88813 397292
rect 90035 397356 90101 397357
rect 90035 397292 90036 397356
rect 90100 397292 90101 397356
rect 90035 397291 90101 397292
rect 90774 396813 90834 399470
rect 91326 397357 91386 399470
rect 92430 398173 92490 399470
rect 93350 399470 93524 399530
rect 93600 399530 93660 400106
rect 94552 399530 94612 400106
rect 93600 399470 93778 399530
rect 92427 398172 92493 398173
rect 92427 398108 92428 398172
rect 92492 398108 92493 398172
rect 92427 398107 92493 398108
rect 91323 397356 91389 397357
rect 91323 397292 91324 397356
rect 91388 397292 91389 397356
rect 91323 397291 91389 397292
rect 86539 396812 86605 396813
rect 86539 396748 86540 396812
rect 86604 396748 86605 396812
rect 86539 396747 86605 396748
rect 88379 396812 88445 396813
rect 88379 396748 88380 396812
rect 88444 396748 88445 396812
rect 88379 396747 88445 396748
rect 90771 396812 90837 396813
rect 90771 396748 90772 396812
rect 90836 396748 90837 396812
rect 90771 396747 90837 396748
rect 84954 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 85574 374614
rect 84954 374294 85574 374378
rect 84954 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 85574 374294
rect 84954 338614 85574 374058
rect 84954 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 85574 338614
rect 84954 338294 85574 338378
rect 84954 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 85574 338294
rect 84954 302614 85574 338058
rect 84954 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 85574 302614
rect 84954 302294 85574 302378
rect 84954 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 85574 302294
rect 84954 266614 85574 302058
rect 84954 266378 84986 266614
rect 85222 266378 85306 266614
rect 85542 266378 85574 266614
rect 84954 266294 85574 266378
rect 84954 266058 84986 266294
rect 85222 266058 85306 266294
rect 85542 266058 85574 266294
rect 84954 230614 85574 266058
rect 84954 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 85574 230614
rect 84954 230294 85574 230378
rect 84954 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 85574 230294
rect 84954 228675 85574 230058
rect 91794 381454 92414 398000
rect 93350 396677 93410 399470
rect 93718 396813 93778 399470
rect 94454 399470 94612 399530
rect 95912 399530 95972 400106
rect 96048 399530 96108 400106
rect 97000 399530 97060 400106
rect 98088 399530 98148 400106
rect 98496 399530 98556 400106
rect 99448 399530 99508 400106
rect 95912 399470 95986 399530
rect 96048 399470 96354 399530
rect 97000 399470 97090 399530
rect 98088 399470 98194 399530
rect 98496 399470 98562 399530
rect 94454 397357 94514 399470
rect 95926 398173 95986 399470
rect 95923 398172 95989 398173
rect 95923 398108 95924 398172
rect 95988 398108 95989 398172
rect 95923 398107 95989 398108
rect 94451 397356 94517 397357
rect 94451 397292 94452 397356
rect 94516 397292 94517 397356
rect 94451 397291 94517 397292
rect 93715 396812 93781 396813
rect 93715 396748 93716 396812
rect 93780 396748 93781 396812
rect 93715 396747 93781 396748
rect 93347 396676 93413 396677
rect 93347 396612 93348 396676
rect 93412 396612 93413 396676
rect 93347 396611 93413 396612
rect 91794 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 92414 381454
rect 91794 381134 92414 381218
rect 91794 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 92414 381134
rect 91794 345454 92414 380898
rect 91794 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 92414 345454
rect 91794 345134 92414 345218
rect 91794 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 92414 345134
rect 91794 309454 92414 344898
rect 91794 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 92414 309454
rect 91794 309134 92414 309218
rect 91794 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 92414 309134
rect 91794 273454 92414 308898
rect 91794 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 92414 273454
rect 91794 273134 92414 273218
rect 91794 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 92414 273134
rect 91794 237454 92414 272898
rect 91794 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 92414 237454
rect 91794 237134 92414 237218
rect 91794 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 92414 237134
rect 91794 228675 92414 236898
rect 95514 385174 96134 398000
rect 96294 396813 96354 399470
rect 97030 397357 97090 399470
rect 97027 397356 97093 397357
rect 97027 397292 97028 397356
rect 97092 397292 97093 397356
rect 97027 397291 97093 397292
rect 96291 396812 96357 396813
rect 96291 396748 96292 396812
rect 96356 396748 96357 396812
rect 96291 396747 96357 396748
rect 98134 396677 98194 399470
rect 98502 396813 98562 399470
rect 99422 399470 99508 399530
rect 100672 399530 100732 400106
rect 101080 399530 101140 400106
rect 100672 399470 100770 399530
rect 99422 398173 99482 399470
rect 99419 398172 99485 398173
rect 99419 398108 99420 398172
rect 99484 398108 99485 398172
rect 99419 398107 99485 398108
rect 98499 396812 98565 396813
rect 98499 396748 98500 396812
rect 98564 396748 98565 396812
rect 98499 396747 98565 396748
rect 98131 396676 98197 396677
rect 98131 396612 98132 396676
rect 98196 396612 98197 396676
rect 98131 396611 98197 396612
rect 95514 384938 95546 385174
rect 95782 384938 95866 385174
rect 96102 384938 96134 385174
rect 95514 384854 96134 384938
rect 95514 384618 95546 384854
rect 95782 384618 95866 384854
rect 96102 384618 96134 384854
rect 95514 349174 96134 384618
rect 95514 348938 95546 349174
rect 95782 348938 95866 349174
rect 96102 348938 96134 349174
rect 95514 348854 96134 348938
rect 95514 348618 95546 348854
rect 95782 348618 95866 348854
rect 96102 348618 96134 348854
rect 95514 313174 96134 348618
rect 95514 312938 95546 313174
rect 95782 312938 95866 313174
rect 96102 312938 96134 313174
rect 95514 312854 96134 312938
rect 95514 312618 95546 312854
rect 95782 312618 95866 312854
rect 96102 312618 96134 312854
rect 95514 277174 96134 312618
rect 95514 276938 95546 277174
rect 95782 276938 95866 277174
rect 96102 276938 96134 277174
rect 95514 276854 96134 276938
rect 95514 276618 95546 276854
rect 95782 276618 95866 276854
rect 96102 276618 96134 276854
rect 95514 241174 96134 276618
rect 95514 240938 95546 241174
rect 95782 240938 95866 241174
rect 96102 240938 96134 241174
rect 95514 240854 96134 240938
rect 95514 240618 95546 240854
rect 95782 240618 95866 240854
rect 96102 240618 96134 240854
rect 95514 228675 96134 240618
rect 99234 388894 99854 398000
rect 100710 397357 100770 399470
rect 101078 399470 101140 399530
rect 101760 399530 101820 400106
rect 102848 399530 102908 400106
rect 101760 399470 101874 399530
rect 100707 397356 100773 397357
rect 100707 397292 100708 397356
rect 100772 397292 100773 397356
rect 100707 397291 100773 397292
rect 101078 396813 101138 399470
rect 101814 397357 101874 399470
rect 102734 399470 102908 399530
rect 103528 399530 103588 400106
rect 103936 399530 103996 400106
rect 105296 399530 105356 400106
rect 105976 399530 106036 400106
rect 106384 399530 106444 400106
rect 107608 399530 107668 400106
rect 108288 399530 108348 400106
rect 103528 399470 103714 399530
rect 103936 399470 104082 399530
rect 105296 399470 105370 399530
rect 105976 399470 106106 399530
rect 106384 399470 106474 399530
rect 101811 397356 101877 397357
rect 101811 397292 101812 397356
rect 101876 397292 101877 397356
rect 101811 397291 101877 397292
rect 102734 396813 102794 399470
rect 101075 396812 101141 396813
rect 101075 396748 101076 396812
rect 101140 396748 101141 396812
rect 101075 396747 101141 396748
rect 102731 396812 102797 396813
rect 102731 396748 102732 396812
rect 102796 396748 102797 396812
rect 102731 396747 102797 396748
rect 99234 388658 99266 388894
rect 99502 388658 99586 388894
rect 99822 388658 99854 388894
rect 99234 388574 99854 388658
rect 99234 388338 99266 388574
rect 99502 388338 99586 388574
rect 99822 388338 99854 388574
rect 99234 352894 99854 388338
rect 99234 352658 99266 352894
rect 99502 352658 99586 352894
rect 99822 352658 99854 352894
rect 99234 352574 99854 352658
rect 99234 352338 99266 352574
rect 99502 352338 99586 352574
rect 99822 352338 99854 352574
rect 99234 316894 99854 352338
rect 99234 316658 99266 316894
rect 99502 316658 99586 316894
rect 99822 316658 99854 316894
rect 99234 316574 99854 316658
rect 99234 316338 99266 316574
rect 99502 316338 99586 316574
rect 99822 316338 99854 316574
rect 99234 280894 99854 316338
rect 99234 280658 99266 280894
rect 99502 280658 99586 280894
rect 99822 280658 99854 280894
rect 99234 280574 99854 280658
rect 99234 280338 99266 280574
rect 99502 280338 99586 280574
rect 99822 280338 99854 280574
rect 99234 244894 99854 280338
rect 99234 244658 99266 244894
rect 99502 244658 99586 244894
rect 99822 244658 99854 244894
rect 99234 244574 99854 244658
rect 99234 244338 99266 244574
rect 99502 244338 99586 244574
rect 99822 244338 99854 244574
rect 99234 228675 99854 244338
rect 102954 392614 103574 398000
rect 103654 396810 103714 399470
rect 104022 397357 104082 399470
rect 104019 397356 104085 397357
rect 104019 397292 104020 397356
rect 104084 397292 104085 397356
rect 104019 397291 104085 397292
rect 105310 396813 105370 399470
rect 106046 396813 106106 399470
rect 106414 397357 106474 399470
rect 107518 399470 107668 399530
rect 108254 399470 108348 399530
rect 108696 399530 108756 400106
rect 109784 399530 109844 400106
rect 108696 399470 108866 399530
rect 106411 397356 106477 397357
rect 106411 397292 106412 397356
rect 106476 397292 106477 397356
rect 106411 397291 106477 397292
rect 107518 396813 107578 399470
rect 103835 396812 103901 396813
rect 103835 396810 103836 396812
rect 103654 396750 103836 396810
rect 103835 396748 103836 396750
rect 103900 396748 103901 396812
rect 103835 396747 103901 396748
rect 105307 396812 105373 396813
rect 105307 396748 105308 396812
rect 105372 396748 105373 396812
rect 105307 396747 105373 396748
rect 106043 396812 106109 396813
rect 106043 396748 106044 396812
rect 106108 396748 106109 396812
rect 106043 396747 106109 396748
rect 107515 396812 107581 396813
rect 107515 396748 107516 396812
rect 107580 396748 107581 396812
rect 107515 396747 107581 396748
rect 108254 396677 108314 399470
rect 108806 396813 108866 399470
rect 109542 399470 109844 399530
rect 111008 399530 111068 400106
rect 111144 399530 111204 400106
rect 112232 399530 112292 400106
rect 113320 399530 113380 400106
rect 111008 399470 111074 399530
rect 111144 399470 111258 399530
rect 109542 397357 109602 399470
rect 109539 397356 109605 397357
rect 109539 397292 109540 397356
rect 109604 397292 109605 397356
rect 109539 397291 109605 397292
rect 108803 396812 108869 396813
rect 108803 396748 108804 396812
rect 108868 396748 108869 396812
rect 108803 396747 108869 396748
rect 108251 396676 108317 396677
rect 108251 396612 108252 396676
rect 108316 396612 108317 396676
rect 108251 396611 108317 396612
rect 102954 392378 102986 392614
rect 103222 392378 103306 392614
rect 103542 392378 103574 392614
rect 102954 392294 103574 392378
rect 102954 392058 102986 392294
rect 103222 392058 103306 392294
rect 103542 392058 103574 392294
rect 102954 356614 103574 392058
rect 102954 356378 102986 356614
rect 103222 356378 103306 356614
rect 103542 356378 103574 356614
rect 102954 356294 103574 356378
rect 102954 356058 102986 356294
rect 103222 356058 103306 356294
rect 103542 356058 103574 356294
rect 102954 320614 103574 356058
rect 102954 320378 102986 320614
rect 103222 320378 103306 320614
rect 103542 320378 103574 320614
rect 102954 320294 103574 320378
rect 102954 320058 102986 320294
rect 103222 320058 103306 320294
rect 103542 320058 103574 320294
rect 102954 284614 103574 320058
rect 102954 284378 102986 284614
rect 103222 284378 103306 284614
rect 103542 284378 103574 284614
rect 102954 284294 103574 284378
rect 102954 284058 102986 284294
rect 103222 284058 103306 284294
rect 103542 284058 103574 284294
rect 102954 248614 103574 284058
rect 102954 248378 102986 248614
rect 103222 248378 103306 248614
rect 103542 248378 103574 248614
rect 102954 248294 103574 248378
rect 102954 248058 102986 248294
rect 103222 248058 103306 248294
rect 103542 248058 103574 248294
rect 102954 228675 103574 248058
rect 109794 363454 110414 398000
rect 111014 396813 111074 399470
rect 111198 397357 111258 399470
rect 112118 399470 112292 399530
rect 113222 399470 113380 399530
rect 112118 397357 112178 399470
rect 113222 397357 113282 399470
rect 113590 398173 113650 400136
rect 114408 399530 114468 400106
rect 114326 399470 114468 399530
rect 113587 398172 113653 398173
rect 113587 398108 113588 398172
rect 113652 398108 113653 398172
rect 113587 398107 113653 398108
rect 111195 397356 111261 397357
rect 111195 397292 111196 397356
rect 111260 397292 111261 397356
rect 111195 397291 111261 397292
rect 112115 397356 112181 397357
rect 112115 397292 112116 397356
rect 112180 397292 112181 397356
rect 112115 397291 112181 397292
rect 113219 397356 113285 397357
rect 113219 397292 113220 397356
rect 113284 397292 113285 397356
rect 113219 397291 113285 397292
rect 111011 396812 111077 396813
rect 111011 396748 111012 396812
rect 111076 396748 111077 396812
rect 111011 396747 111077 396748
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 327454 110414 362898
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 109794 291454 110414 326898
rect 109794 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 110414 291454
rect 109794 291134 110414 291218
rect 109794 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 110414 291134
rect 109794 255454 110414 290898
rect 109794 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 110414 255454
rect 109794 255134 110414 255218
rect 109794 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 110414 255134
rect 109794 228675 110414 254898
rect 113514 367174 114134 398000
rect 114326 397357 114386 399470
rect 115798 397357 115858 400136
rect 115982 400076 116070 400136
rect 114323 397356 114389 397357
rect 114323 397292 114324 397356
rect 114388 397292 114389 397356
rect 114323 397291 114389 397292
rect 115795 397356 115861 397357
rect 115795 397292 115796 397356
rect 115860 397292 115861 397356
rect 115795 397291 115861 397292
rect 115982 396813 116042 400076
rect 116992 399530 117052 400106
rect 118080 399530 118140 400106
rect 118488 399530 118548 400106
rect 119168 399530 119228 400106
rect 120936 399530 120996 400106
rect 116992 399470 117146 399530
rect 118080 399470 118250 399530
rect 118488 399470 118618 399530
rect 117086 397357 117146 399470
rect 117083 397356 117149 397357
rect 117083 397292 117084 397356
rect 117148 397292 117149 397356
rect 117083 397291 117149 397292
rect 115979 396812 116045 396813
rect 115979 396748 115980 396812
rect 116044 396748 116045 396812
rect 115979 396747 116045 396748
rect 113514 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 114134 367174
rect 113514 366854 114134 366938
rect 113514 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 114134 366854
rect 113514 331174 114134 366618
rect 113514 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 114134 331174
rect 113514 330854 114134 330938
rect 113514 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 114134 330854
rect 113514 295174 114134 330618
rect 113514 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 114134 295174
rect 113514 294854 114134 294938
rect 113514 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 114134 294854
rect 113514 259174 114134 294618
rect 113514 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 114134 259174
rect 113514 258854 114134 258938
rect 113514 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 114134 258854
rect 113514 228675 114134 258618
rect 117234 370894 117854 398000
rect 118190 397357 118250 399470
rect 118558 397357 118618 399470
rect 119110 399470 119228 399530
rect 120766 399470 120996 399530
rect 123520 399530 123580 400106
rect 125968 399530 126028 400106
rect 123520 399470 123586 399530
rect 118187 397356 118253 397357
rect 118187 397292 118188 397356
rect 118252 397292 118253 397356
rect 118187 397291 118253 397292
rect 118555 397356 118621 397357
rect 118555 397292 118556 397356
rect 118620 397292 118621 397356
rect 118555 397291 118621 397292
rect 119110 396813 119170 399470
rect 120766 396813 120826 399470
rect 119107 396812 119173 396813
rect 119107 396748 119108 396812
rect 119172 396748 119173 396812
rect 119107 396747 119173 396748
rect 120763 396812 120829 396813
rect 120763 396748 120764 396812
rect 120828 396748 120829 396812
rect 120763 396747 120829 396748
rect 117234 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 117854 370894
rect 117234 370574 117854 370658
rect 117234 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 117854 370574
rect 117234 334894 117854 370338
rect 117234 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 117854 334894
rect 117234 334574 117854 334658
rect 117234 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 117854 334574
rect 117234 298894 117854 334338
rect 117234 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 117854 298894
rect 117234 298574 117854 298658
rect 117234 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 117854 298574
rect 117234 262894 117854 298338
rect 117234 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 117854 262894
rect 117234 262574 117854 262658
rect 117234 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 117854 262574
rect 117234 228675 117854 262338
rect 120954 374614 121574 398000
rect 123526 397357 123586 399470
rect 125918 399470 126028 399530
rect 128280 399530 128340 400106
rect 131000 399530 131060 400106
rect 128280 399470 128554 399530
rect 125918 397357 125978 399470
rect 123523 397356 123589 397357
rect 123523 397292 123524 397356
rect 123588 397292 123589 397356
rect 123523 397291 123589 397292
rect 125915 397356 125981 397357
rect 125915 397292 125916 397356
rect 125980 397292 125981 397356
rect 125915 397291 125981 397292
rect 120954 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 121574 374614
rect 120954 374294 121574 374378
rect 120954 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 121574 374294
rect 120954 338614 121574 374058
rect 120954 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 121574 338614
rect 120954 338294 121574 338378
rect 120954 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 121574 338294
rect 120954 302614 121574 338058
rect 120954 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 121574 302614
rect 120954 302294 121574 302378
rect 120954 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 121574 302294
rect 120954 266614 121574 302058
rect 120954 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 121574 266614
rect 120954 266294 121574 266378
rect 120954 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 121574 266294
rect 120954 230614 121574 266058
rect 120954 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 121574 230614
rect 120954 230294 121574 230378
rect 120954 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 121574 230294
rect 120954 228675 121574 230058
rect 127794 381454 128414 398000
rect 128494 396130 128554 399470
rect 130886 399470 131060 399530
rect 133448 399530 133508 400106
rect 135896 399530 135956 400106
rect 138480 399530 138540 400106
rect 140928 399530 140988 400106
rect 133448 399470 133522 399530
rect 135896 399470 136098 399530
rect 130886 396813 130946 399470
rect 130883 396812 130949 396813
rect 130883 396748 130884 396812
rect 130948 396748 130949 396812
rect 130883 396747 130949 396748
rect 128675 396132 128741 396133
rect 128675 396130 128676 396132
rect 128494 396070 128676 396130
rect 128675 396068 128676 396070
rect 128740 396068 128741 396132
rect 128675 396067 128741 396068
rect 127794 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 128414 381454
rect 127794 381134 128414 381218
rect 127794 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 128414 381134
rect 127794 345454 128414 380898
rect 127794 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 128414 345454
rect 127794 345134 128414 345218
rect 127794 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 128414 345134
rect 127794 309454 128414 344898
rect 127794 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 128414 309454
rect 127794 309134 128414 309218
rect 127794 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 128414 309134
rect 127794 273454 128414 308898
rect 127794 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 128414 273454
rect 127794 273134 128414 273218
rect 127794 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 128414 273134
rect 127794 237454 128414 272898
rect 127794 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 128414 237454
rect 127794 237134 128414 237218
rect 127794 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 128414 237134
rect 127794 228675 128414 236898
rect 131514 385174 132134 398000
rect 133462 396813 133522 399470
rect 133459 396812 133525 396813
rect 133459 396748 133460 396812
rect 133524 396748 133525 396812
rect 133459 396747 133525 396748
rect 131514 384938 131546 385174
rect 131782 384938 131866 385174
rect 132102 384938 132134 385174
rect 131514 384854 132134 384938
rect 131514 384618 131546 384854
rect 131782 384618 131866 384854
rect 132102 384618 132134 384854
rect 131514 349174 132134 384618
rect 131514 348938 131546 349174
rect 131782 348938 131866 349174
rect 132102 348938 132134 349174
rect 131514 348854 132134 348938
rect 131514 348618 131546 348854
rect 131782 348618 131866 348854
rect 132102 348618 132134 348854
rect 131514 313174 132134 348618
rect 131514 312938 131546 313174
rect 131782 312938 131866 313174
rect 132102 312938 132134 313174
rect 131514 312854 132134 312938
rect 131514 312618 131546 312854
rect 131782 312618 131866 312854
rect 132102 312618 132134 312854
rect 131514 277174 132134 312618
rect 131514 276938 131546 277174
rect 131782 276938 131866 277174
rect 132102 276938 132134 277174
rect 131514 276854 132134 276938
rect 131514 276618 131546 276854
rect 131782 276618 131866 276854
rect 132102 276618 132134 276854
rect 131514 241174 132134 276618
rect 131514 240938 131546 241174
rect 131782 240938 131866 241174
rect 132102 240938 132134 241174
rect 131514 240854 132134 240938
rect 131514 240618 131546 240854
rect 131782 240618 131866 240854
rect 132102 240618 132134 240854
rect 131514 228675 132134 240618
rect 135234 388894 135854 398000
rect 136038 397357 136098 399470
rect 138430 399470 138540 399530
rect 140822 399470 140988 399530
rect 143512 399530 143572 400106
rect 145960 399530 146020 400106
rect 148544 399530 148604 400106
rect 150992 399530 151052 400106
rect 143512 399470 143642 399530
rect 145960 399470 146034 399530
rect 148544 399470 148610 399530
rect 138430 397357 138490 399470
rect 136035 397356 136101 397357
rect 136035 397292 136036 397356
rect 136100 397292 136101 397356
rect 136035 397291 136101 397292
rect 138427 397356 138493 397357
rect 138427 397292 138428 397356
rect 138492 397292 138493 397356
rect 138427 397291 138493 397292
rect 135234 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 135854 388894
rect 135234 388574 135854 388658
rect 135234 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 135854 388574
rect 135234 352894 135854 388338
rect 135234 352658 135266 352894
rect 135502 352658 135586 352894
rect 135822 352658 135854 352894
rect 135234 352574 135854 352658
rect 135234 352338 135266 352574
rect 135502 352338 135586 352574
rect 135822 352338 135854 352574
rect 135234 316894 135854 352338
rect 135234 316658 135266 316894
rect 135502 316658 135586 316894
rect 135822 316658 135854 316894
rect 135234 316574 135854 316658
rect 135234 316338 135266 316574
rect 135502 316338 135586 316574
rect 135822 316338 135854 316574
rect 135234 280894 135854 316338
rect 135234 280658 135266 280894
rect 135502 280658 135586 280894
rect 135822 280658 135854 280894
rect 135234 280574 135854 280658
rect 135234 280338 135266 280574
rect 135502 280338 135586 280574
rect 135822 280338 135854 280574
rect 135234 244894 135854 280338
rect 135234 244658 135266 244894
rect 135502 244658 135586 244894
rect 135822 244658 135854 244894
rect 135234 244574 135854 244658
rect 135234 244338 135266 244574
rect 135502 244338 135586 244574
rect 135822 244338 135854 244574
rect 135234 228675 135854 244338
rect 138954 392614 139574 398000
rect 140822 396813 140882 399470
rect 143582 396813 143642 399470
rect 145974 398173 146034 399470
rect 145971 398172 146037 398173
rect 145971 398108 145972 398172
rect 146036 398108 146037 398172
rect 145971 398107 146037 398108
rect 140819 396812 140885 396813
rect 140819 396748 140820 396812
rect 140884 396748 140885 396812
rect 140819 396747 140885 396748
rect 143579 396812 143645 396813
rect 143579 396748 143580 396812
rect 143644 396748 143645 396812
rect 143579 396747 143645 396748
rect 138954 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 139574 392614
rect 138954 392294 139574 392378
rect 138954 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 139574 392294
rect 138954 356614 139574 392058
rect 138954 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 139574 356614
rect 138954 356294 139574 356378
rect 138954 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 139574 356294
rect 138954 320614 139574 356058
rect 138954 320378 138986 320614
rect 139222 320378 139306 320614
rect 139542 320378 139574 320614
rect 138954 320294 139574 320378
rect 138954 320058 138986 320294
rect 139222 320058 139306 320294
rect 139542 320058 139574 320294
rect 138954 284614 139574 320058
rect 138954 284378 138986 284614
rect 139222 284378 139306 284614
rect 139542 284378 139574 284614
rect 138954 284294 139574 284378
rect 138954 284058 138986 284294
rect 139222 284058 139306 284294
rect 139542 284058 139574 284294
rect 138954 248614 139574 284058
rect 138954 248378 138986 248614
rect 139222 248378 139306 248614
rect 139542 248378 139574 248614
rect 138954 248294 139574 248378
rect 138954 248058 138986 248294
rect 139222 248058 139306 248294
rect 139542 248058 139574 248294
rect 138954 228675 139574 248058
rect 145794 363454 146414 398000
rect 148550 396813 148610 399470
rect 150942 399470 151052 399530
rect 153440 399530 153500 400106
rect 155888 399530 155948 400106
rect 158472 399530 158532 400106
rect 160920 399530 160980 400106
rect 153440 399470 154130 399530
rect 155888 399470 155970 399530
rect 158472 399470 158546 399530
rect 148547 396812 148613 396813
rect 148547 396748 148548 396812
rect 148612 396748 148613 396812
rect 148547 396747 148613 396748
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 327454 146414 362898
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 145794 291454 146414 326898
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 255454 146414 290898
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 228675 146414 254898
rect 149514 367174 150134 398000
rect 150942 396813 151002 399470
rect 150939 396812 151005 396813
rect 150939 396748 150940 396812
rect 151004 396748 151005 396812
rect 150939 396747 151005 396748
rect 149514 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 150134 367174
rect 149514 366854 150134 366938
rect 149514 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 150134 366854
rect 149514 331174 150134 366618
rect 149514 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 150134 331174
rect 149514 330854 150134 330938
rect 149514 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 150134 330854
rect 149514 295174 150134 330618
rect 149514 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 150134 295174
rect 149514 294854 150134 294938
rect 149514 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 150134 294854
rect 149514 259174 150134 294618
rect 149514 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 150134 259174
rect 149514 258854 150134 258938
rect 149514 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 150134 258854
rect 149514 228675 150134 258618
rect 153234 370894 153854 398000
rect 154070 396813 154130 399470
rect 155910 397357 155970 399470
rect 155907 397356 155973 397357
rect 155907 397292 155908 397356
rect 155972 397292 155973 397356
rect 155907 397291 155973 397292
rect 154067 396812 154133 396813
rect 154067 396748 154068 396812
rect 154132 396748 154133 396812
rect 154067 396747 154133 396748
rect 153234 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 153854 370894
rect 153234 370574 153854 370658
rect 153234 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 153854 370574
rect 153234 334894 153854 370338
rect 153234 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 153854 334894
rect 153234 334574 153854 334658
rect 153234 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 153854 334574
rect 153234 298894 153854 334338
rect 153234 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 153854 298894
rect 153234 298574 153854 298658
rect 153234 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 153854 298574
rect 153234 262894 153854 298338
rect 153234 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 153854 262894
rect 153234 262574 153854 262658
rect 153234 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 153854 262574
rect 153234 228675 153854 262338
rect 156954 374614 157574 398000
rect 158486 396813 158546 399470
rect 160878 399470 160980 399530
rect 163368 399530 163428 400106
rect 165952 399530 166012 400106
rect 183224 399530 183284 400106
rect 163368 399470 163514 399530
rect 160878 396813 160938 399470
rect 163454 397357 163514 399470
rect 165846 399470 166012 399530
rect 183142 399470 183284 399530
rect 183360 399530 183420 400106
rect 183360 399470 183570 399530
rect 163451 397356 163517 397357
rect 163451 397292 163452 397356
rect 163516 397292 163517 397356
rect 163451 397291 163517 397292
rect 158483 396812 158549 396813
rect 158483 396748 158484 396812
rect 158548 396748 158549 396812
rect 158483 396747 158549 396748
rect 160875 396812 160941 396813
rect 160875 396748 160876 396812
rect 160940 396748 160941 396812
rect 160875 396747 160941 396748
rect 156954 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 157574 374614
rect 156954 374294 157574 374378
rect 156954 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 157574 374294
rect 156954 338614 157574 374058
rect 156954 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 157574 338614
rect 156954 338294 157574 338378
rect 156954 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 157574 338294
rect 156954 302614 157574 338058
rect 156954 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 157574 302614
rect 156954 302294 157574 302378
rect 156954 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 157574 302294
rect 156954 266614 157574 302058
rect 156954 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 157574 266614
rect 156954 266294 157574 266378
rect 156954 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 157574 266294
rect 156954 230614 157574 266058
rect 156954 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 157574 230614
rect 156954 230294 157574 230378
rect 156954 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 157574 230294
rect 156954 228675 157574 230058
rect 163794 381454 164414 398000
rect 165846 396813 165906 399470
rect 165843 396812 165909 396813
rect 165843 396748 165844 396812
rect 165908 396748 165909 396812
rect 165843 396747 165909 396748
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 163794 345454 164414 380898
rect 163794 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 164414 345454
rect 163794 345134 164414 345218
rect 163794 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 164414 345134
rect 163794 309454 164414 344898
rect 163794 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 164414 309454
rect 163794 309134 164414 309218
rect 163794 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 164414 309134
rect 163794 273454 164414 308898
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 163794 237454 164414 272898
rect 163794 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 164414 237454
rect 163794 237134 164414 237218
rect 163794 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 164414 237134
rect 163794 228675 164414 236898
rect 167514 385174 168134 398000
rect 167514 384938 167546 385174
rect 167782 384938 167866 385174
rect 168102 384938 168134 385174
rect 167514 384854 168134 384938
rect 167514 384618 167546 384854
rect 167782 384618 167866 384854
rect 168102 384618 168134 384854
rect 167514 349174 168134 384618
rect 167514 348938 167546 349174
rect 167782 348938 167866 349174
rect 168102 348938 168134 349174
rect 167514 348854 168134 348938
rect 167514 348618 167546 348854
rect 167782 348618 167866 348854
rect 168102 348618 168134 348854
rect 167514 313174 168134 348618
rect 167514 312938 167546 313174
rect 167782 312938 167866 313174
rect 168102 312938 168134 313174
rect 167514 312854 168134 312938
rect 167514 312618 167546 312854
rect 167782 312618 167866 312854
rect 168102 312618 168134 312854
rect 167514 277174 168134 312618
rect 167514 276938 167546 277174
rect 167782 276938 167866 277174
rect 168102 276938 168134 277174
rect 167514 276854 168134 276938
rect 167514 276618 167546 276854
rect 167782 276618 167866 276854
rect 168102 276618 168134 276854
rect 167514 241174 168134 276618
rect 167514 240938 167546 241174
rect 167782 240938 167866 241174
rect 168102 240938 168134 241174
rect 167514 240854 168134 240938
rect 167514 240618 167546 240854
rect 167782 240618 167866 240854
rect 168102 240618 168134 240854
rect 167514 228675 168134 240618
rect 171234 388894 171854 398000
rect 171234 388658 171266 388894
rect 171502 388658 171586 388894
rect 171822 388658 171854 388894
rect 171234 388574 171854 388658
rect 171234 388338 171266 388574
rect 171502 388338 171586 388574
rect 171822 388338 171854 388574
rect 171234 352894 171854 388338
rect 171234 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 171854 352894
rect 171234 352574 171854 352658
rect 171234 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 171854 352574
rect 171234 316894 171854 352338
rect 171234 316658 171266 316894
rect 171502 316658 171586 316894
rect 171822 316658 171854 316894
rect 171234 316574 171854 316658
rect 171234 316338 171266 316574
rect 171502 316338 171586 316574
rect 171822 316338 171854 316574
rect 171234 280894 171854 316338
rect 171234 280658 171266 280894
rect 171502 280658 171586 280894
rect 171822 280658 171854 280894
rect 171234 280574 171854 280658
rect 171234 280338 171266 280574
rect 171502 280338 171586 280574
rect 171822 280338 171854 280574
rect 171234 244894 171854 280338
rect 171234 244658 171266 244894
rect 171502 244658 171586 244894
rect 171822 244658 171854 244894
rect 171234 244574 171854 244658
rect 171234 244338 171266 244574
rect 171502 244338 171586 244574
rect 171822 244338 171854 244574
rect 171234 228675 171854 244338
rect 174954 392614 175574 398000
rect 174954 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 175574 392614
rect 174954 392294 175574 392378
rect 174954 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 175574 392294
rect 174954 356614 175574 392058
rect 174954 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 175574 356614
rect 174954 356294 175574 356378
rect 174954 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 175574 356294
rect 174954 320614 175574 356058
rect 174954 320378 174986 320614
rect 175222 320378 175306 320614
rect 175542 320378 175574 320614
rect 174954 320294 175574 320378
rect 174954 320058 174986 320294
rect 175222 320058 175306 320294
rect 175542 320058 175574 320294
rect 174954 284614 175574 320058
rect 174954 284378 174986 284614
rect 175222 284378 175306 284614
rect 175542 284378 175574 284614
rect 174954 284294 175574 284378
rect 174954 284058 174986 284294
rect 175222 284058 175306 284294
rect 175542 284058 175574 284294
rect 174954 248614 175574 284058
rect 174954 248378 174986 248614
rect 175222 248378 175306 248614
rect 175542 248378 175574 248614
rect 174954 248294 175574 248378
rect 174954 248058 174986 248294
rect 175222 248058 175306 248294
rect 175542 248058 175574 248294
rect 174954 228675 175574 248058
rect 181794 363454 182414 398000
rect 183142 396813 183202 399470
rect 183510 396813 183570 399470
rect 183139 396812 183205 396813
rect 183139 396748 183140 396812
rect 183204 396748 183205 396812
rect 183139 396747 183205 396748
rect 183507 396812 183573 396813
rect 183507 396748 183508 396812
rect 183572 396748 183573 396812
rect 183507 396747 183573 396748
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 255454 182414 290898
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 181794 228675 182414 254898
rect 185514 367174 186134 398000
rect 185514 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 186134 367174
rect 185514 366854 186134 366938
rect 185514 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 186134 366854
rect 185514 331174 186134 366618
rect 185514 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 186134 331174
rect 185514 330854 186134 330938
rect 185514 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 186134 330854
rect 185514 295174 186134 330618
rect 185514 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 186134 295174
rect 185514 294854 186134 294938
rect 185514 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 186134 294854
rect 185514 259174 186134 294618
rect 185514 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 186134 259174
rect 185514 258854 186134 258938
rect 185514 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 186134 258854
rect 185514 228675 186134 258618
rect 189234 370894 189854 398000
rect 189234 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 189854 370894
rect 189234 370574 189854 370658
rect 189234 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 189854 370574
rect 189234 334894 189854 370338
rect 189234 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 189854 334894
rect 189234 334574 189854 334658
rect 189234 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 189854 334574
rect 189234 298894 189854 334338
rect 189234 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 189854 298894
rect 189234 298574 189854 298658
rect 189234 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 189854 298574
rect 189234 262894 189854 298338
rect 189234 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 189854 262894
rect 189234 262574 189854 262658
rect 189234 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 189854 262574
rect 189234 228675 189854 262338
rect 192954 374614 193574 398000
rect 192954 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 193574 374614
rect 192954 374294 193574 374378
rect 192954 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 193574 374294
rect 192954 338614 193574 374058
rect 192954 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 193574 338614
rect 192954 338294 193574 338378
rect 192954 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 193574 338294
rect 192954 302614 193574 338058
rect 192954 302378 192986 302614
rect 193222 302378 193306 302614
rect 193542 302378 193574 302614
rect 192954 302294 193574 302378
rect 192954 302058 192986 302294
rect 193222 302058 193306 302294
rect 193542 302058 193574 302294
rect 192954 266614 193574 302058
rect 192954 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 193574 266614
rect 192954 266294 193574 266378
rect 192954 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 193574 266294
rect 192954 230614 193574 266058
rect 192954 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 193574 230614
rect 192954 230294 193574 230378
rect 192954 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 193574 230294
rect 192954 228675 193574 230058
rect 199794 381454 200414 416898
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 199794 345454 200414 380898
rect 199794 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 200414 345454
rect 199794 345134 200414 345218
rect 199794 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 200414 345134
rect 199794 309454 200414 344898
rect 199794 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 200414 309454
rect 199794 309134 200414 309218
rect 199794 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 200414 309134
rect 199794 273454 200414 308898
rect 199794 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 200414 273454
rect 199794 273134 200414 273218
rect 199794 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 200414 273134
rect 199794 237454 200414 272898
rect 199794 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 200414 237454
rect 199794 237134 200414 237218
rect 199794 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 200414 237134
rect 199794 228675 200414 236898
rect 203514 673174 204134 707162
rect 203514 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 204134 673174
rect 203514 672854 204134 672938
rect 203514 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 204134 672854
rect 203514 637174 204134 672618
rect 203514 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 204134 637174
rect 203514 636854 204134 636938
rect 203514 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 204134 636854
rect 203514 601174 204134 636618
rect 203514 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 204134 601174
rect 203514 600854 204134 600938
rect 203514 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 204134 600854
rect 203514 565174 204134 600618
rect 203514 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 204134 565174
rect 203514 564854 204134 564938
rect 203514 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 204134 564854
rect 203514 529174 204134 564618
rect 203514 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 204134 529174
rect 203514 528854 204134 528938
rect 203514 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 204134 528854
rect 203514 493174 204134 528618
rect 203514 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 204134 493174
rect 203514 492854 204134 492938
rect 203514 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 204134 492854
rect 203514 457174 204134 492618
rect 203514 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 204134 457174
rect 203514 456854 204134 456938
rect 203514 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 204134 456854
rect 203514 421174 204134 456618
rect 203514 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 204134 421174
rect 203514 420854 204134 420938
rect 203514 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 204134 420854
rect 203514 385174 204134 420618
rect 203514 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 204134 385174
rect 203514 384854 204134 384938
rect 203514 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 204134 384854
rect 203514 349174 204134 384618
rect 203514 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 204134 349174
rect 203514 348854 204134 348938
rect 203514 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 204134 348854
rect 203514 313174 204134 348618
rect 203514 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 204134 313174
rect 203514 312854 204134 312938
rect 203514 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 204134 312854
rect 203514 277174 204134 312618
rect 203514 276938 203546 277174
rect 203782 276938 203866 277174
rect 204102 276938 204134 277174
rect 203514 276854 204134 276938
rect 203514 276618 203546 276854
rect 203782 276618 203866 276854
rect 204102 276618 204134 276854
rect 203514 241174 204134 276618
rect 203514 240938 203546 241174
rect 203782 240938 203866 241174
rect 204102 240938 204134 241174
rect 203514 240854 204134 240938
rect 203514 240618 203546 240854
rect 203782 240618 203866 240854
rect 204102 240618 204134 240854
rect 203514 228675 204134 240618
rect 207234 676894 207854 709082
rect 207234 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 207854 676894
rect 207234 676574 207854 676658
rect 207234 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 207854 676574
rect 207234 640894 207854 676338
rect 207234 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 207854 640894
rect 207234 640574 207854 640658
rect 207234 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 207854 640574
rect 207234 604894 207854 640338
rect 207234 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 207854 604894
rect 207234 604574 207854 604658
rect 207234 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 207854 604574
rect 207234 568894 207854 604338
rect 207234 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 207854 568894
rect 207234 568574 207854 568658
rect 207234 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 207854 568574
rect 207234 532894 207854 568338
rect 207234 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 207854 532894
rect 207234 532574 207854 532658
rect 207234 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 207854 532574
rect 207234 496894 207854 532338
rect 207234 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 207854 496894
rect 207234 496574 207854 496658
rect 207234 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 207854 496574
rect 207234 460894 207854 496338
rect 207234 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 207854 460894
rect 207234 460574 207854 460658
rect 207234 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 207854 460574
rect 207234 424894 207854 460338
rect 207234 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 207854 424894
rect 207234 424574 207854 424658
rect 207234 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 207854 424574
rect 207234 388894 207854 424338
rect 207234 388658 207266 388894
rect 207502 388658 207586 388894
rect 207822 388658 207854 388894
rect 207234 388574 207854 388658
rect 207234 388338 207266 388574
rect 207502 388338 207586 388574
rect 207822 388338 207854 388574
rect 207234 352894 207854 388338
rect 207234 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 207854 352894
rect 207234 352574 207854 352658
rect 207234 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 207854 352574
rect 207234 316894 207854 352338
rect 207234 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 207854 316894
rect 207234 316574 207854 316658
rect 207234 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 207854 316574
rect 207234 280894 207854 316338
rect 207234 280658 207266 280894
rect 207502 280658 207586 280894
rect 207822 280658 207854 280894
rect 207234 280574 207854 280658
rect 207234 280338 207266 280574
rect 207502 280338 207586 280574
rect 207822 280338 207854 280574
rect 207234 244894 207854 280338
rect 207234 244658 207266 244894
rect 207502 244658 207586 244894
rect 207822 244658 207854 244894
rect 207234 244574 207854 244658
rect 207234 244338 207266 244574
rect 207502 244338 207586 244574
rect 207822 244338 207854 244574
rect 207234 228675 207854 244338
rect 210954 680614 211574 711002
rect 228954 710598 229574 711590
rect 228954 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 229574 710598
rect 228954 710278 229574 710362
rect 228954 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 229574 710278
rect 225234 708678 225854 709670
rect 225234 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 225854 708678
rect 225234 708358 225854 708442
rect 225234 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 225854 708358
rect 221514 706758 222134 707750
rect 221514 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 222134 706758
rect 221514 706438 222134 706522
rect 221514 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 222134 706438
rect 210954 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 211574 680614
rect 210954 680294 211574 680378
rect 210954 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 211574 680294
rect 210954 644614 211574 680058
rect 210954 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 211574 644614
rect 210954 644294 211574 644378
rect 210954 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 211574 644294
rect 210954 608614 211574 644058
rect 210954 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 211574 608614
rect 210954 608294 211574 608378
rect 210954 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 211574 608294
rect 210954 572614 211574 608058
rect 210954 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 211574 572614
rect 210954 572294 211574 572378
rect 210954 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 211574 572294
rect 210954 536614 211574 572058
rect 210954 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 211574 536614
rect 210954 536294 211574 536378
rect 210954 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 211574 536294
rect 210954 500614 211574 536058
rect 210954 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 211574 500614
rect 210954 500294 211574 500378
rect 210954 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 211574 500294
rect 210954 464614 211574 500058
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 507454 218414 542898
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217794 485308 218414 506898
rect 221514 691174 222134 706202
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 655174 222134 690618
rect 221514 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 222134 655174
rect 221514 654854 222134 654938
rect 221514 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 222134 654854
rect 221514 619174 222134 654618
rect 221514 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 222134 619174
rect 221514 618854 222134 618938
rect 221514 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 222134 618854
rect 221514 583174 222134 618618
rect 221514 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 222134 583174
rect 221514 582854 222134 582938
rect 221514 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 222134 582854
rect 221514 547174 222134 582618
rect 221514 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 222134 547174
rect 221514 546854 222134 546938
rect 221514 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 222134 546854
rect 221514 511174 222134 546618
rect 221514 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 222134 511174
rect 221514 510854 222134 510938
rect 221514 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 222134 510854
rect 218651 505204 218717 505205
rect 218651 505140 218652 505204
rect 218716 505140 218717 505204
rect 218651 505139 218717 505140
rect 210954 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 211574 464614
rect 210954 464294 211574 464378
rect 210954 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 211574 464294
rect 210954 428614 211574 464058
rect 210954 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 211574 428614
rect 210954 428294 211574 428378
rect 210954 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 211574 428294
rect 210954 392614 211574 428058
rect 210954 392378 210986 392614
rect 211222 392378 211306 392614
rect 211542 392378 211574 392614
rect 210954 392294 211574 392378
rect 210954 392058 210986 392294
rect 211222 392058 211306 392294
rect 211542 392058 211574 392294
rect 210954 356614 211574 392058
rect 210954 356378 210986 356614
rect 211222 356378 211306 356614
rect 211542 356378 211574 356614
rect 210954 356294 211574 356378
rect 210954 356058 210986 356294
rect 211222 356058 211306 356294
rect 211542 356058 211574 356294
rect 210954 320614 211574 356058
rect 210954 320378 210986 320614
rect 211222 320378 211306 320614
rect 211542 320378 211574 320614
rect 210954 320294 211574 320378
rect 210954 320058 210986 320294
rect 211222 320058 211306 320294
rect 211542 320058 211574 320294
rect 210954 284614 211574 320058
rect 210954 284378 210986 284614
rect 211222 284378 211306 284614
rect 211542 284378 211574 284614
rect 210954 284294 211574 284378
rect 210954 284058 210986 284294
rect 211222 284058 211306 284294
rect 211542 284058 211574 284294
rect 210954 248614 211574 284058
rect 210954 248378 210986 248614
rect 211222 248378 211306 248614
rect 211542 248378 211574 248614
rect 210954 248294 211574 248378
rect 210954 248058 210986 248294
rect 211222 248058 211306 248294
rect 211542 248058 211574 248294
rect 210954 228675 211574 248058
rect 217794 363454 218414 398000
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 327454 218414 362898
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 217794 291454 218414 326898
rect 217794 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 218414 291454
rect 217794 291134 218414 291218
rect 217794 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 218414 291134
rect 217794 255454 218414 290898
rect 217794 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 218414 255454
rect 217794 255134 218414 255218
rect 217794 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 218414 255134
rect 217794 228675 218414 254898
rect 218654 230349 218714 505139
rect 219755 486028 219821 486029
rect 219755 485964 219756 486028
rect 219820 485964 219821 486028
rect 219755 485963 219821 485964
rect 219758 480997 219818 485963
rect 221514 485308 222134 510618
rect 225234 694894 225854 708122
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 658894 225854 694338
rect 225234 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 225854 658894
rect 225234 658574 225854 658658
rect 225234 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 225854 658574
rect 225234 622894 225854 658338
rect 225234 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 225854 622894
rect 225234 622574 225854 622658
rect 225234 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 225854 622574
rect 225234 586894 225854 622338
rect 225234 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 225854 586894
rect 225234 586574 225854 586658
rect 225234 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 225854 586574
rect 225234 550894 225854 586338
rect 225234 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 225854 550894
rect 225234 550574 225854 550658
rect 225234 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 225854 550574
rect 225234 514894 225854 550338
rect 225234 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 225854 514894
rect 225234 514574 225854 514658
rect 225234 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 225854 514574
rect 225234 485308 225854 514338
rect 228954 698614 229574 710042
rect 246954 711558 247574 711590
rect 246954 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 247574 711558
rect 246954 711238 247574 711322
rect 246954 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 247574 711238
rect 243234 709638 243854 709670
rect 243234 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 243854 709638
rect 243234 709318 243854 709402
rect 243234 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 243854 709318
rect 239514 707718 240134 707750
rect 239514 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 240134 707718
rect 239514 707398 240134 707482
rect 239514 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 240134 707398
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 662614 229574 698058
rect 228954 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 229574 662614
rect 228954 662294 229574 662378
rect 228954 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 229574 662294
rect 228954 626614 229574 662058
rect 228954 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 229574 626614
rect 228954 626294 229574 626378
rect 228954 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 229574 626294
rect 228954 590614 229574 626058
rect 228954 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 229574 590614
rect 228954 590294 229574 590378
rect 228954 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 229574 590294
rect 228954 554614 229574 590058
rect 228954 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 229574 554614
rect 228954 554294 229574 554378
rect 228954 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 229574 554294
rect 228954 518614 229574 554058
rect 228954 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 229574 518614
rect 228954 518294 229574 518378
rect 228954 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 229574 518294
rect 228954 485308 229574 518058
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 235794 669454 236414 705242
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561454 236414 596898
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 525454 236414 560898
rect 235794 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 236414 525454
rect 235794 525134 236414 525218
rect 235794 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 236414 525134
rect 235794 489454 236414 524898
rect 235794 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 236414 489454
rect 235794 489134 236414 489218
rect 235794 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 236414 489134
rect 235794 485308 236414 488898
rect 239514 673174 240134 707162
rect 239514 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 240134 673174
rect 239514 672854 240134 672938
rect 239514 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 240134 672854
rect 239514 637174 240134 672618
rect 239514 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 240134 637174
rect 239514 636854 240134 636938
rect 239514 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 240134 636854
rect 239514 601174 240134 636618
rect 239514 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 240134 601174
rect 239514 600854 240134 600938
rect 239514 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 240134 600854
rect 239514 565174 240134 600618
rect 239514 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 240134 565174
rect 239514 564854 240134 564938
rect 239514 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 240134 564854
rect 239514 529174 240134 564618
rect 239514 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 240134 529174
rect 239514 528854 240134 528938
rect 239514 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 240134 528854
rect 239514 493174 240134 528618
rect 239514 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 240134 493174
rect 239514 492854 240134 492938
rect 239514 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 240134 492854
rect 239514 485308 240134 492618
rect 243234 676894 243854 709082
rect 243234 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 243854 676894
rect 243234 676574 243854 676658
rect 243234 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 243854 676574
rect 243234 640894 243854 676338
rect 243234 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 243854 640894
rect 243234 640574 243854 640658
rect 243234 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 243854 640574
rect 243234 604894 243854 640338
rect 243234 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 243854 604894
rect 243234 604574 243854 604658
rect 243234 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 243854 604574
rect 243234 568894 243854 604338
rect 243234 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 243854 568894
rect 243234 568574 243854 568658
rect 243234 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 243854 568574
rect 243234 532894 243854 568338
rect 243234 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 243854 532894
rect 243234 532574 243854 532658
rect 243234 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 243854 532574
rect 243234 496894 243854 532338
rect 243234 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 243854 496894
rect 243234 496574 243854 496658
rect 243234 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 243854 496574
rect 243234 485308 243854 496338
rect 246954 680614 247574 711002
rect 264954 710598 265574 711590
rect 264954 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 265574 710598
rect 264954 710278 265574 710362
rect 264954 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 265574 710278
rect 261234 708678 261854 709670
rect 261234 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 261854 708678
rect 261234 708358 261854 708442
rect 261234 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 261854 708358
rect 257514 706758 258134 707750
rect 257514 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 258134 706758
rect 257514 706438 258134 706522
rect 257514 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 258134 706438
rect 246954 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 247574 680614
rect 246954 680294 247574 680378
rect 246954 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 247574 680294
rect 246954 644614 247574 680058
rect 246954 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 247574 644614
rect 246954 644294 247574 644378
rect 246954 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 247574 644294
rect 246954 608614 247574 644058
rect 246954 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 247574 608614
rect 246954 608294 247574 608378
rect 246954 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 247574 608294
rect 246954 572614 247574 608058
rect 246954 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 247574 572614
rect 246954 572294 247574 572378
rect 246954 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 247574 572294
rect 246954 536614 247574 572058
rect 246954 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 247574 536614
rect 246954 536294 247574 536378
rect 246954 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 247574 536294
rect 246954 500614 247574 536058
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 507454 254414 542898
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 248459 504252 248525 504253
rect 248459 504188 248460 504252
rect 248524 504188 248525 504252
rect 248459 504187 248525 504188
rect 246954 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 247574 500614
rect 246954 500294 247574 500378
rect 246954 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 247574 500294
rect 246954 485308 247574 500058
rect 248462 487170 248522 504187
rect 251035 503572 251101 503573
rect 251035 503508 251036 503572
rect 251100 503508 251101 503572
rect 251035 503507 251101 503508
rect 248462 487110 248706 487170
rect 248646 483850 248706 487110
rect 251038 483850 251098 503507
rect 253289 487660 253355 487661
rect 253289 487596 253290 487660
rect 253354 487596 253355 487660
rect 253289 487595 253355 487596
rect 253292 487250 253352 487595
rect 248646 483790 248764 483850
rect 248704 483202 248764 483790
rect 251016 483790 251098 483850
rect 253246 487190 253352 487250
rect 253246 483850 253306 487190
rect 253794 485308 254414 506898
rect 257514 691174 258134 706202
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 655174 258134 690618
rect 257514 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 258134 655174
rect 257514 654854 258134 654938
rect 257514 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 258134 654854
rect 257514 619174 258134 654618
rect 257514 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 258134 619174
rect 257514 618854 258134 618938
rect 257514 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 258134 618854
rect 257514 583174 258134 618618
rect 257514 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 258134 583174
rect 257514 582854 258134 582938
rect 257514 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 258134 582854
rect 257514 547174 258134 582618
rect 257514 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 258134 547174
rect 257514 546854 258134 546938
rect 257514 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 258134 546854
rect 257514 511174 258134 546618
rect 257514 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 258134 511174
rect 257514 510854 258134 510938
rect 257514 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 258134 510854
rect 256187 503844 256253 503845
rect 256187 503780 256188 503844
rect 256252 503780 256253 503844
rect 256187 503779 256253 503780
rect 256190 483850 256250 503779
rect 257514 485308 258134 510618
rect 261234 694894 261854 708122
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 658894 261854 694338
rect 261234 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 261854 658894
rect 261234 658574 261854 658658
rect 261234 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 261854 658574
rect 261234 622894 261854 658338
rect 261234 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 261854 622894
rect 261234 622574 261854 622658
rect 261234 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 261854 622574
rect 261234 586894 261854 622338
rect 261234 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 261854 586894
rect 261234 586574 261854 586658
rect 261234 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 261854 586574
rect 261234 550894 261854 586338
rect 261234 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 261854 550894
rect 261234 550574 261854 550658
rect 261234 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 261854 550574
rect 261234 514894 261854 550338
rect 261234 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 261854 514894
rect 261234 514574 261854 514658
rect 261234 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 261854 514574
rect 258395 503980 258461 503981
rect 258395 503916 258396 503980
rect 258460 503916 258461 503980
rect 258395 503915 258461 503916
rect 258398 495450 258458 503915
rect 260971 503572 261037 503573
rect 260971 503508 260972 503572
rect 261036 503508 261037 503572
rect 260971 503507 261037 503508
rect 258214 495390 258458 495450
rect 258214 494070 258274 495390
rect 258214 494010 258458 494070
rect 258398 487170 258458 494010
rect 260974 487170 261034 503507
rect 258398 487110 258642 487170
rect 260974 487110 261140 487170
rect 258582 483850 258642 487110
rect 261080 486570 261140 487110
rect 260974 486510 261140 486570
rect 260974 485210 261034 486510
rect 261234 485308 261854 514338
rect 264954 698614 265574 710042
rect 282954 711558 283574 711590
rect 282954 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 283574 711558
rect 282954 711238 283574 711322
rect 282954 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 283574 711238
rect 279234 709638 279854 709670
rect 279234 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 279854 709638
rect 279234 709318 279854 709402
rect 279234 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 279854 709318
rect 275514 707718 276134 707750
rect 275514 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 276134 707718
rect 275514 707398 276134 707482
rect 275514 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 276134 707398
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 662614 265574 698058
rect 264954 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 265574 662614
rect 264954 662294 265574 662378
rect 264954 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 265574 662294
rect 264954 626614 265574 662058
rect 264954 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 265574 626614
rect 264954 626294 265574 626378
rect 264954 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 265574 626294
rect 264954 590614 265574 626058
rect 264954 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 265574 590614
rect 264954 590294 265574 590378
rect 264954 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 265574 590294
rect 264954 554614 265574 590058
rect 264954 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 265574 554614
rect 264954 554294 265574 554378
rect 264954 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 265574 554294
rect 264954 518614 265574 554058
rect 264954 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 265574 518614
rect 264954 518294 265574 518378
rect 264954 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 265574 518294
rect 263685 487660 263751 487661
rect 263685 487596 263686 487660
rect 263750 487596 263751 487660
rect 263685 487595 263751 487596
rect 263688 487250 263748 487595
rect 263550 487190 263748 487250
rect 260974 485150 261218 485210
rect 261158 483850 261218 485150
rect 263550 483850 263610 487190
rect 264954 485308 265574 518058
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 271794 669454 272414 705242
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 525454 272414 560898
rect 271794 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 272414 525454
rect 271794 525134 272414 525218
rect 271794 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 272414 525134
rect 266123 503572 266189 503573
rect 266123 503508 266124 503572
rect 266188 503508 266189 503572
rect 266123 503507 266189 503508
rect 267779 503572 267845 503573
rect 267779 503508 267780 503572
rect 267844 503508 267845 503572
rect 267779 503507 267845 503508
rect 270539 503572 270605 503573
rect 270539 503508 270540 503572
rect 270604 503508 270605 503572
rect 270539 503507 270605 503508
rect 266126 483850 266186 503507
rect 253246 483790 253524 483850
rect 251016 483202 251076 483790
rect 253464 483202 253524 483790
rect 256184 483790 256250 483850
rect 258496 483790 258642 483850
rect 261080 483790 261218 483850
rect 263528 483790 263610 483850
rect 266112 483790 266186 483850
rect 267782 483850 267842 503507
rect 270542 483850 270602 503507
rect 271794 489454 272414 524898
rect 275514 673174 276134 707162
rect 275514 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 276134 673174
rect 275514 672854 276134 672938
rect 275514 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 276134 672854
rect 275514 637174 276134 672618
rect 275514 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 276134 637174
rect 275514 636854 276134 636938
rect 275514 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 276134 636854
rect 275514 601174 276134 636618
rect 275514 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 276134 601174
rect 275514 600854 276134 600938
rect 275514 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 276134 600854
rect 275514 565174 276134 600618
rect 275514 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 276134 565174
rect 275514 564854 276134 564938
rect 275514 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 276134 564854
rect 275514 529174 276134 564618
rect 275514 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 276134 529174
rect 275514 528854 276134 528938
rect 275514 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 276134 528854
rect 273299 503572 273365 503573
rect 273299 503508 273300 503572
rect 273364 503508 273365 503572
rect 273299 503507 273365 503508
rect 271794 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 272414 489454
rect 271794 489134 272414 489218
rect 271794 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 272414 489134
rect 271794 485308 272414 488898
rect 273302 483850 273362 503507
rect 275514 493174 276134 528618
rect 279234 676894 279854 709082
rect 279234 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 279854 676894
rect 279234 676574 279854 676658
rect 279234 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 279854 676574
rect 279234 640894 279854 676338
rect 279234 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 279854 640894
rect 279234 640574 279854 640658
rect 279234 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 279854 640574
rect 279234 604894 279854 640338
rect 279234 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 279854 604894
rect 279234 604574 279854 604658
rect 279234 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 279854 604574
rect 279234 568894 279854 604338
rect 279234 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 279854 568894
rect 279234 568574 279854 568658
rect 279234 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 279854 568574
rect 279234 532894 279854 568338
rect 279234 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 279854 532894
rect 279234 532574 279854 532658
rect 279234 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 279854 532574
rect 278451 503708 278517 503709
rect 278451 503644 278452 503708
rect 278516 503644 278517 503708
rect 278451 503643 278517 503644
rect 276243 503572 276309 503573
rect 276243 503508 276244 503572
rect 276308 503508 276309 503572
rect 276243 503507 276309 503508
rect 275514 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 276134 493174
rect 275514 492854 276134 492938
rect 275514 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 276134 492854
rect 275514 485308 276134 492618
rect 276246 483850 276306 503507
rect 267782 483790 268620 483850
rect 270542 483790 271204 483850
rect 273302 483790 273652 483850
rect 256184 483202 256244 483790
rect 258496 483202 258556 483790
rect 261080 483202 261140 483790
rect 263528 483202 263588 483790
rect 266112 483202 266172 483790
rect 268560 483202 268620 483790
rect 271144 483202 271204 483790
rect 273592 483202 273652 483790
rect 276176 483790 276306 483850
rect 278454 483850 278514 503643
rect 279234 496894 279854 532338
rect 282954 680614 283574 711002
rect 300954 710598 301574 711590
rect 300954 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 301574 710598
rect 300954 710278 301574 710362
rect 300954 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 301574 710278
rect 297234 708678 297854 709670
rect 297234 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 297854 708678
rect 297234 708358 297854 708442
rect 297234 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 297854 708358
rect 293514 706758 294134 707750
rect 293514 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 294134 706758
rect 293514 706438 294134 706522
rect 293514 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 294134 706438
rect 282954 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 283574 680614
rect 282954 680294 283574 680378
rect 282954 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 283574 680294
rect 282954 644614 283574 680058
rect 282954 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 283574 644614
rect 282954 644294 283574 644378
rect 282954 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 283574 644294
rect 282954 608614 283574 644058
rect 282954 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 283574 608614
rect 282954 608294 283574 608378
rect 282954 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 283574 608294
rect 282954 572614 283574 608058
rect 282954 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 283574 572614
rect 282954 572294 283574 572378
rect 282954 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 283574 572294
rect 282954 536614 283574 572058
rect 282954 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 283574 536614
rect 282954 536294 283574 536378
rect 282954 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 283574 536294
rect 280107 503572 280173 503573
rect 280107 503508 280108 503572
rect 280172 503508 280173 503572
rect 280107 503507 280173 503508
rect 279234 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 279854 496894
rect 279234 496574 279854 496658
rect 279234 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 279854 496574
rect 279234 485308 279854 496338
rect 280110 488550 280170 503507
rect 282954 500614 283574 536058
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 288571 503708 288637 503709
rect 288571 503644 288572 503708
rect 288636 503644 288637 503708
rect 288571 503643 288637 503644
rect 285627 503572 285693 503573
rect 285627 503508 285628 503572
rect 285692 503508 285693 503572
rect 285627 503507 285693 503508
rect 282954 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 283574 500614
rect 282954 500294 283574 500378
rect 282954 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 283574 500294
rect 280110 488490 280906 488550
rect 280846 483850 280906 488490
rect 282954 485308 283574 500058
rect 285630 487930 285690 503507
rect 285630 487870 286058 487930
rect 284385 487660 284451 487661
rect 284385 487596 284386 487660
rect 284450 487596 284451 487660
rect 284385 487595 284451 487596
rect 284388 487250 284448 487595
rect 283790 487190 284448 487250
rect 283790 483850 283850 487190
rect 278454 483790 278548 483850
rect 280846 483790 280996 483850
rect 276176 483202 276236 483790
rect 278488 483202 278548 483790
rect 280936 483202 280996 483790
rect 283656 483790 283850 483850
rect 285998 483850 286058 487870
rect 288574 483850 288634 503643
rect 289794 485308 290414 506898
rect 293514 691174 294134 706202
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 655174 294134 690618
rect 293514 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 294134 655174
rect 293514 654854 294134 654938
rect 293514 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 294134 654854
rect 293514 619174 294134 654618
rect 293514 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 294134 619174
rect 293514 618854 294134 618938
rect 293514 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 294134 618854
rect 293514 583174 294134 618618
rect 293514 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 294134 583174
rect 293514 582854 294134 582938
rect 293514 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 294134 582854
rect 293514 547174 294134 582618
rect 293514 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 294134 547174
rect 293514 546854 294134 546938
rect 293514 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 294134 546854
rect 293514 511174 294134 546618
rect 293514 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 294134 511174
rect 293514 510854 294134 510938
rect 293514 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 294134 510854
rect 290963 503572 291029 503573
rect 290963 503508 290964 503572
rect 291028 503508 291029 503572
rect 290963 503507 291029 503508
rect 292619 503572 292685 503573
rect 292619 503508 292620 503572
rect 292684 503508 292685 503572
rect 292619 503507 292685 503508
rect 285998 483790 286164 483850
rect 283656 483202 283716 483790
rect 286104 483202 286164 483790
rect 288552 483790 288634 483850
rect 290966 483850 291026 503507
rect 292622 494050 292682 503507
rect 292622 493990 292866 494050
rect 292806 485890 292866 493990
rect 292806 485830 293418 485890
rect 293358 483850 293418 485830
rect 293514 485308 294134 510618
rect 297234 694894 297854 708122
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 658894 297854 694338
rect 297234 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 297854 658894
rect 297234 658574 297854 658658
rect 297234 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 297854 658574
rect 297234 622894 297854 658338
rect 297234 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 297854 622894
rect 297234 622574 297854 622658
rect 297234 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 297854 622574
rect 297234 586894 297854 622338
rect 297234 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 297854 586894
rect 297234 586574 297854 586658
rect 297234 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 297854 586574
rect 297234 550894 297854 586338
rect 297234 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 297854 550894
rect 297234 550574 297854 550658
rect 297234 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 297854 550574
rect 297234 514894 297854 550338
rect 297234 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 297854 514894
rect 297234 514574 297854 514658
rect 297234 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 297854 514574
rect 295379 503572 295445 503573
rect 295379 503508 295380 503572
rect 295444 503508 295445 503572
rect 295379 503507 295445 503508
rect 295382 483850 295442 503507
rect 297234 485308 297854 514338
rect 300954 698614 301574 710042
rect 318954 711558 319574 711590
rect 318954 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 319574 711558
rect 318954 711238 319574 711322
rect 318954 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 319574 711238
rect 315234 709638 315854 709670
rect 315234 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 315854 709638
rect 315234 709318 315854 709402
rect 315234 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 315854 709318
rect 311514 707718 312134 707750
rect 311514 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 312134 707718
rect 311514 707398 312134 707482
rect 311514 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 312134 707398
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 662614 301574 698058
rect 300954 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 301574 662614
rect 300954 662294 301574 662378
rect 300954 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 301574 662294
rect 300954 626614 301574 662058
rect 300954 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 301574 626614
rect 300954 626294 301574 626378
rect 300954 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 301574 626294
rect 300954 590614 301574 626058
rect 300954 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 301574 590614
rect 300954 590294 301574 590378
rect 300954 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 301574 590294
rect 300954 554614 301574 590058
rect 300954 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 301574 554614
rect 300954 554294 301574 554378
rect 300954 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 301574 554294
rect 300954 518614 301574 554058
rect 300954 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 301574 518614
rect 300954 518294 301574 518378
rect 300954 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 301574 518294
rect 300954 492693 301574 518058
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 669454 308414 705242
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 298139 492692 298205 492693
rect 298139 492628 298140 492692
rect 298204 492628 298205 492692
rect 300899 492692 301574 492693
rect 300899 492690 300900 492692
rect 298139 492627 298205 492628
rect 300718 492630 300900 492690
rect 298142 483850 298202 492627
rect 300718 485210 300778 492630
rect 300899 492628 300900 492630
rect 300964 492628 301574 492692
rect 300899 492627 301574 492628
rect 302187 492692 302253 492693
rect 302187 492628 302188 492692
rect 302252 492628 302253 492692
rect 302187 492627 302253 492628
rect 304947 492692 305013 492693
rect 304947 492628 304948 492692
rect 305012 492628 305013 492692
rect 307707 492692 307773 492693
rect 307707 492690 307708 492692
rect 304947 492627 305013 492628
rect 307526 492630 307708 492690
rect 300954 485308 301574 492627
rect 300718 485150 300962 485210
rect 300902 483850 300962 485150
rect 302190 483850 302250 492627
rect 304950 483850 305010 492627
rect 307526 485210 307586 492630
rect 307707 492628 307708 492630
rect 307772 492628 307773 492692
rect 307707 492627 307773 492628
rect 307794 489454 308414 524898
rect 311514 673174 312134 707162
rect 311514 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 312134 673174
rect 311514 672854 312134 672938
rect 311514 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 312134 672854
rect 311514 637174 312134 672618
rect 311514 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 312134 637174
rect 311514 636854 312134 636938
rect 311514 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 312134 636854
rect 311514 601174 312134 636618
rect 311514 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 312134 601174
rect 311514 600854 312134 600938
rect 311514 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 312134 600854
rect 311514 565174 312134 600618
rect 311514 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 312134 565174
rect 311514 564854 312134 564938
rect 311514 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 312134 564854
rect 311514 529174 312134 564618
rect 311514 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 312134 529174
rect 311514 528854 312134 528938
rect 311514 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 312134 528854
rect 311514 493174 312134 528618
rect 311514 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 312134 493174
rect 311514 492854 312134 492938
rect 310467 492692 310533 492693
rect 310467 492628 310468 492692
rect 310532 492628 310533 492692
rect 310467 492627 310533 492628
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 307794 485308 308414 488898
rect 307526 485150 308322 485210
rect 308262 483850 308322 485150
rect 310470 483850 310530 492627
rect 311514 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 312134 492854
rect 315234 676894 315854 709082
rect 315234 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 315854 676894
rect 315234 676574 315854 676658
rect 315234 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 315854 676574
rect 315234 640894 315854 676338
rect 315234 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 315854 640894
rect 315234 640574 315854 640658
rect 315234 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 315854 640574
rect 315234 604894 315854 640338
rect 315234 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 315854 604894
rect 315234 604574 315854 604658
rect 315234 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 315854 604574
rect 315234 568894 315854 604338
rect 315234 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 315854 568894
rect 315234 568574 315854 568658
rect 315234 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 315854 568574
rect 315234 532894 315854 568338
rect 315234 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 315854 532894
rect 315234 532574 315854 532658
rect 315234 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 315854 532574
rect 315234 496894 315854 532338
rect 315234 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 315854 496894
rect 315234 496574 315854 496658
rect 315234 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 315854 496574
rect 313227 492692 313293 492693
rect 313227 492628 313228 492692
rect 313292 492628 313293 492692
rect 313227 492627 313293 492628
rect 311514 485308 312134 492618
rect 313230 483850 313290 492627
rect 315234 485308 315854 496338
rect 318954 680614 319574 711002
rect 336954 710598 337574 711590
rect 336954 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 337574 710598
rect 336954 710278 337574 710362
rect 336954 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 337574 710278
rect 333234 708678 333854 709670
rect 333234 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 333854 708678
rect 333234 708358 333854 708442
rect 333234 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 333854 708358
rect 329514 706758 330134 707750
rect 329514 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 330134 706758
rect 329514 706438 330134 706522
rect 329514 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 330134 706438
rect 318954 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 319574 680614
rect 318954 680294 319574 680378
rect 318954 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 319574 680294
rect 318954 644614 319574 680058
rect 318954 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 319574 644614
rect 318954 644294 319574 644378
rect 318954 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 319574 644294
rect 318954 608614 319574 644058
rect 318954 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 319574 608614
rect 318954 608294 319574 608378
rect 318954 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 319574 608294
rect 318954 572614 319574 608058
rect 318954 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 319574 572614
rect 318954 572294 319574 572378
rect 318954 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 319574 572294
rect 318954 536614 319574 572058
rect 318954 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 319574 536614
rect 318954 536294 319574 536378
rect 318954 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 319574 536294
rect 318954 500614 319574 536058
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 323347 503572 323413 503573
rect 323347 503508 323348 503572
rect 323412 503508 323413 503572
rect 323347 503507 323413 503508
rect 318954 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 319574 500614
rect 318954 500294 319574 500378
rect 318954 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 319574 500294
rect 316021 492692 316087 492693
rect 316021 492690 316022 492692
rect 315990 492628 316022 492690
rect 316086 492628 316087 492692
rect 315990 492627 316087 492628
rect 317459 492692 317525 492693
rect 317459 492628 317460 492692
rect 317524 492628 317525 492692
rect 317459 492627 317525 492628
rect 315990 489930 316050 492627
rect 315990 489870 316234 489930
rect 316174 483850 316234 489870
rect 317462 488550 317522 492627
rect 317462 488490 318442 488550
rect 290966 483790 291060 483850
rect 293358 483790 293644 483850
rect 295382 483790 295956 483850
rect 298142 483790 298676 483850
rect 300902 483790 301124 483850
rect 302190 483790 303572 483850
rect 304950 483790 306020 483850
rect 308262 483790 308468 483850
rect 310470 483790 311052 483850
rect 313230 483790 313636 483850
rect 288552 483202 288612 483790
rect 291000 483202 291060 483790
rect 293584 483202 293644 483790
rect 295896 483202 295956 483790
rect 298616 483202 298676 483790
rect 301064 483202 301124 483790
rect 303512 483202 303572 483790
rect 305960 483202 306020 483790
rect 308408 483202 308468 483790
rect 310992 483202 311052 483790
rect 313576 483202 313636 483790
rect 316024 483790 316234 483850
rect 318382 483850 318442 488490
rect 318954 485308 319574 500058
rect 320219 492692 320285 492693
rect 320219 492628 320220 492692
rect 320284 492628 320285 492692
rect 320219 492627 320285 492628
rect 320222 488550 320282 492627
rect 323350 488550 323410 503507
rect 320038 488490 320282 488550
rect 323166 488490 323410 488550
rect 320038 485890 320098 488490
rect 320038 485830 320190 485890
rect 320130 485790 320190 485830
rect 320130 485730 320834 485790
rect 320774 483850 320834 485730
rect 323166 484410 323226 488490
rect 325794 485308 326414 506898
rect 329514 691174 330134 706202
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 655174 330134 690618
rect 329514 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 330134 655174
rect 329514 654854 330134 654938
rect 329514 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 330134 654854
rect 329514 619174 330134 654618
rect 329514 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 330134 619174
rect 329514 618854 330134 618938
rect 329514 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 330134 618854
rect 329514 583174 330134 618618
rect 329514 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 330134 583174
rect 329514 582854 330134 582938
rect 329514 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 330134 582854
rect 329514 547174 330134 582618
rect 329514 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 330134 547174
rect 329514 546854 330134 546938
rect 329514 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 330134 546854
rect 329514 511174 330134 546618
rect 329514 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 330134 511174
rect 329514 510854 330134 510938
rect 329514 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 330134 510854
rect 326613 488340 326679 488341
rect 326613 488276 326614 488340
rect 326678 488276 326679 488340
rect 326613 488275 326679 488276
rect 326616 487930 326676 488275
rect 326616 487870 326722 487930
rect 323166 484350 323410 484410
rect 318382 483790 318532 483850
rect 320774 483790 321116 483850
rect 316024 483202 316084 483790
rect 318472 483202 318532 483790
rect 321056 483202 321116 483790
rect 323350 483714 323410 484350
rect 326662 483850 326722 487870
rect 329514 485308 330134 510618
rect 333234 694894 333854 708122
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 658894 333854 694338
rect 333234 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 333854 658894
rect 333234 658574 333854 658658
rect 333234 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 333854 658574
rect 333234 622894 333854 658338
rect 333234 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 333854 622894
rect 333234 622574 333854 622658
rect 333234 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 333854 622574
rect 333234 586894 333854 622338
rect 333234 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 333854 586894
rect 333234 586574 333854 586658
rect 333234 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 333854 586574
rect 333234 550894 333854 586338
rect 333234 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 333854 550894
rect 333234 550574 333854 550658
rect 333234 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 333854 550574
rect 333234 514894 333854 550338
rect 333234 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 333854 514894
rect 333234 514574 333854 514658
rect 333234 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 333854 514574
rect 333234 485308 333854 514338
rect 336954 698614 337574 710042
rect 354954 711558 355574 711590
rect 354954 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 355574 711558
rect 354954 711238 355574 711322
rect 354954 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 355574 711238
rect 351234 709638 351854 709670
rect 351234 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 351854 709638
rect 351234 709318 351854 709402
rect 351234 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 351854 709318
rect 347514 707718 348134 707750
rect 347514 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 348134 707718
rect 347514 707398 348134 707482
rect 347514 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 348134 707398
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 662614 337574 698058
rect 336954 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 337574 662614
rect 336954 662294 337574 662378
rect 336954 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 337574 662294
rect 336954 626614 337574 662058
rect 336954 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 337574 626614
rect 336954 626294 337574 626378
rect 336954 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 337574 626294
rect 336954 590614 337574 626058
rect 336954 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 337574 590614
rect 336954 590294 337574 590378
rect 336954 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 337574 590294
rect 336954 554614 337574 590058
rect 336954 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 337574 554614
rect 336954 554294 337574 554378
rect 336954 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 337574 554294
rect 336954 518614 337574 554058
rect 336954 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 337574 518614
rect 336954 518294 337574 518378
rect 336954 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 337574 518294
rect 336954 485308 337574 518058
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 343794 669454 344414 705242
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 525454 344414 560898
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 339355 492692 339421 492693
rect 339355 492628 339356 492692
rect 339420 492628 339421 492692
rect 339355 492627 339421 492628
rect 339539 492692 339605 492693
rect 339539 492628 339540 492692
rect 339604 492628 339605 492692
rect 339539 492627 339605 492628
rect 339358 483850 339418 492627
rect 326088 483790 326722 483850
rect 338464 483790 339418 483850
rect 339542 483850 339602 492627
rect 343794 489454 344414 524898
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 343794 485308 344414 488898
rect 347514 673174 348134 707162
rect 347514 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 348134 673174
rect 347514 672854 348134 672938
rect 347514 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 348134 672854
rect 347514 637174 348134 672618
rect 347514 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 348134 637174
rect 347514 636854 348134 636938
rect 347514 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 348134 636854
rect 347514 601174 348134 636618
rect 347514 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 348134 601174
rect 347514 600854 348134 600938
rect 347514 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 348134 600854
rect 347514 565174 348134 600618
rect 347514 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 348134 565174
rect 347514 564854 348134 564938
rect 347514 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 348134 564854
rect 347514 529174 348134 564618
rect 347514 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 348134 529174
rect 347514 528854 348134 528938
rect 347514 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 348134 528854
rect 347514 493174 348134 528618
rect 347514 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 348134 493174
rect 347514 492854 348134 492938
rect 347514 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 348134 492854
rect 347514 485308 348134 492618
rect 351234 676894 351854 709082
rect 351234 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 351854 676894
rect 351234 676574 351854 676658
rect 351234 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 351854 676574
rect 351234 640894 351854 676338
rect 351234 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 351854 640894
rect 351234 640574 351854 640658
rect 351234 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 351854 640574
rect 351234 604894 351854 640338
rect 351234 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 351854 604894
rect 351234 604574 351854 604658
rect 351234 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 351854 604574
rect 351234 568894 351854 604338
rect 351234 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 351854 568894
rect 351234 568574 351854 568658
rect 351234 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 351854 568574
rect 351234 532894 351854 568338
rect 351234 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 351854 532894
rect 351234 532574 351854 532658
rect 351234 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 351854 532574
rect 351234 496894 351854 532338
rect 351234 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 351854 496894
rect 351234 496574 351854 496658
rect 351234 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 351854 496574
rect 351234 485308 351854 496338
rect 354954 680614 355574 711002
rect 372954 710598 373574 711590
rect 372954 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 373574 710598
rect 372954 710278 373574 710362
rect 372954 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 373574 710278
rect 369234 708678 369854 709670
rect 369234 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 369854 708678
rect 369234 708358 369854 708442
rect 369234 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 369854 708358
rect 365514 706758 366134 707750
rect 365514 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 366134 706758
rect 365514 706438 366134 706522
rect 365514 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 366134 706438
rect 354954 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 355574 680614
rect 354954 680294 355574 680378
rect 354954 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 355574 680294
rect 354954 644614 355574 680058
rect 354954 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 355574 644614
rect 354954 644294 355574 644378
rect 354954 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 355574 644294
rect 354954 608614 355574 644058
rect 354954 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 355574 608614
rect 354954 608294 355574 608378
rect 354954 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 355574 608294
rect 354954 572614 355574 608058
rect 354954 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 355574 572614
rect 354954 572294 355574 572378
rect 354954 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 355574 572294
rect 354954 536614 355574 572058
rect 354954 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 355574 536614
rect 354954 536294 355574 536378
rect 354954 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 355574 536294
rect 354954 500614 355574 536058
rect 354954 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 355574 500614
rect 354954 500294 355574 500378
rect 354954 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 355574 500294
rect 354954 485308 355574 500058
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 356835 485484 356901 485485
rect 356835 485420 356836 485484
rect 356900 485420 356901 485484
rect 356835 485419 356901 485420
rect 356838 485210 356898 485419
rect 350950 485150 356898 485210
rect 350950 483850 351010 485150
rect 339542 483790 339748 483850
rect 323350 483654 323428 483714
rect 323368 483202 323428 483654
rect 326088 483202 326148 483790
rect 338464 483202 338524 483790
rect 339688 483202 339748 483790
rect 350840 483790 351010 483850
rect 350840 483202 350900 483790
rect 219755 480996 219821 480997
rect 219755 480932 219756 480996
rect 219820 480932 219821 480996
rect 219755 480931 219821 480932
rect 220952 471454 221300 471486
rect 220952 471218 221008 471454
rect 221244 471218 221300 471454
rect 220952 471134 221300 471218
rect 220952 470898 221008 471134
rect 221244 470898 221300 471134
rect 220952 470866 221300 470898
rect 355320 471454 355668 471486
rect 355320 471218 355376 471454
rect 355612 471218 355668 471454
rect 355320 471134 355668 471218
rect 355320 470898 355376 471134
rect 355612 470898 355668 471134
rect 355320 470866 355668 470898
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 220272 453454 220620 453486
rect 220272 453218 220328 453454
rect 220564 453218 220620 453454
rect 220272 453134 220620 453218
rect 220272 452898 220328 453134
rect 220564 452898 220620 453134
rect 220272 452866 220620 452898
rect 356000 453454 356348 453486
rect 356000 453218 356056 453454
rect 356292 453218 356348 453454
rect 356000 453134 356348 453218
rect 356000 452898 356056 453134
rect 356292 452898 356348 453134
rect 356000 452866 356348 452898
rect 220952 435454 221300 435486
rect 220952 435218 221008 435454
rect 221244 435218 221300 435454
rect 220952 435134 221300 435218
rect 220952 434898 221008 435134
rect 221244 434898 221300 435134
rect 220952 434866 221300 434898
rect 355320 435454 355668 435486
rect 355320 435218 355376 435454
rect 355612 435218 355668 435454
rect 355320 435134 355668 435218
rect 355320 434898 355376 435134
rect 355612 434898 355668 435134
rect 355320 434866 355668 434898
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 220272 417454 220620 417486
rect 220272 417218 220328 417454
rect 220564 417218 220620 417454
rect 220272 417134 220620 417218
rect 220272 416898 220328 417134
rect 220564 416898 220620 417134
rect 220272 416866 220620 416898
rect 356000 417454 356348 417486
rect 356000 417218 356056 417454
rect 356292 417218 356348 417454
rect 356000 417134 356348 417218
rect 356000 416898 356056 417134
rect 356292 416898 356348 417134
rect 356000 416866 356348 416898
rect 236056 399530 236116 400106
rect 237144 399530 237204 400106
rect 238232 399530 238292 400106
rect 239592 399530 239652 400106
rect 235950 399470 236116 399530
rect 237054 399470 237204 399530
rect 238158 399470 238292 399530
rect 239262 399470 239652 399530
rect 240544 399530 240604 400106
rect 241768 399530 241828 400106
rect 243128 399530 243188 400106
rect 240544 399470 240610 399530
rect 235950 398173 236010 399470
rect 235947 398172 236013 398173
rect 235947 398108 235948 398172
rect 236012 398108 236013 398172
rect 235947 398107 236013 398108
rect 226379 398036 226445 398037
rect 221514 367174 222134 398000
rect 221514 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 222134 367174
rect 221514 366854 222134 366938
rect 221514 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 222134 366854
rect 221514 331174 222134 366618
rect 221514 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 222134 331174
rect 221514 330854 222134 330938
rect 221514 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 222134 330854
rect 221514 295174 222134 330618
rect 221514 294938 221546 295174
rect 221782 294938 221866 295174
rect 222102 294938 222134 295174
rect 221514 294854 222134 294938
rect 221514 294618 221546 294854
rect 221782 294618 221866 294854
rect 222102 294618 222134 294854
rect 221514 259174 222134 294618
rect 221514 258938 221546 259174
rect 221782 258938 221866 259174
rect 222102 258938 222134 259174
rect 221514 258854 222134 258938
rect 221514 258618 221546 258854
rect 221782 258618 221866 258854
rect 222102 258618 222134 258854
rect 218651 230348 218717 230349
rect 218651 230284 218652 230348
rect 218716 230284 218717 230348
rect 218651 230283 218717 230284
rect 221514 228675 222134 258618
rect 225234 370894 225854 398000
rect 226379 397972 226380 398036
rect 226444 397972 226445 398036
rect 226379 397971 226445 397972
rect 225234 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 225854 370894
rect 225234 370574 225854 370658
rect 225234 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 225854 370574
rect 225234 334894 225854 370338
rect 225234 334658 225266 334894
rect 225502 334658 225586 334894
rect 225822 334658 225854 334894
rect 225234 334574 225854 334658
rect 225234 334338 225266 334574
rect 225502 334338 225586 334574
rect 225822 334338 225854 334574
rect 225234 298894 225854 334338
rect 225234 298658 225266 298894
rect 225502 298658 225586 298894
rect 225822 298658 225854 298894
rect 225234 298574 225854 298658
rect 225234 298338 225266 298574
rect 225502 298338 225586 298574
rect 225822 298338 225854 298574
rect 225234 262894 225854 298338
rect 225234 262658 225266 262894
rect 225502 262658 225586 262894
rect 225822 262658 225854 262894
rect 225234 262574 225854 262658
rect 225234 262338 225266 262574
rect 225502 262338 225586 262574
rect 225822 262338 225854 262574
rect 224907 233068 224973 233069
rect 224907 233004 224908 233068
rect 224972 233004 224973 233068
rect 224907 233003 224973 233004
rect 224910 230890 224970 233003
rect 224726 230830 224970 230890
rect 224726 229530 224786 230830
rect 224907 230348 224973 230349
rect 224907 230284 224908 230348
rect 224972 230284 224973 230348
rect 224907 230283 224973 230284
rect 224910 230210 224970 230283
rect 224910 230150 225154 230210
rect 224726 229470 224970 229530
rect 64208 219454 64528 219486
rect 64208 219218 64250 219454
rect 64486 219218 64528 219454
rect 64208 219134 64528 219218
rect 64208 218898 64250 219134
rect 64486 218898 64528 219134
rect 64208 218866 64528 218898
rect 94928 219454 95248 219486
rect 94928 219218 94970 219454
rect 95206 219218 95248 219454
rect 94928 219134 95248 219218
rect 94928 218898 94970 219134
rect 95206 218898 95248 219134
rect 94928 218866 95248 218898
rect 125648 219454 125968 219486
rect 125648 219218 125690 219454
rect 125926 219218 125968 219454
rect 125648 219134 125968 219218
rect 125648 218898 125690 219134
rect 125926 218898 125968 219134
rect 125648 218866 125968 218898
rect 156368 219454 156688 219486
rect 156368 219218 156410 219454
rect 156646 219218 156688 219454
rect 156368 219134 156688 219218
rect 156368 218898 156410 219134
rect 156646 218898 156688 219134
rect 156368 218866 156688 218898
rect 187088 219454 187408 219486
rect 187088 219218 187130 219454
rect 187366 219218 187408 219454
rect 187088 219134 187408 219218
rect 187088 218898 187130 219134
rect 187366 218898 187408 219134
rect 187088 218866 187408 218898
rect 217808 219454 218128 219486
rect 217808 219218 217850 219454
rect 218086 219218 218128 219454
rect 217808 219134 218128 219218
rect 217808 218898 217850 219134
rect 218086 218898 218128 219134
rect 217808 218866 218128 218898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 79568 201454 79888 201486
rect 79568 201218 79610 201454
rect 79846 201218 79888 201454
rect 79568 201134 79888 201218
rect 79568 200898 79610 201134
rect 79846 200898 79888 201134
rect 79568 200866 79888 200898
rect 110288 201454 110608 201486
rect 110288 201218 110330 201454
rect 110566 201218 110608 201454
rect 110288 201134 110608 201218
rect 110288 200898 110330 201134
rect 110566 200898 110608 201134
rect 110288 200866 110608 200898
rect 141008 201454 141328 201486
rect 141008 201218 141050 201454
rect 141286 201218 141328 201454
rect 141008 201134 141328 201218
rect 141008 200898 141050 201134
rect 141286 200898 141328 201134
rect 141008 200866 141328 200898
rect 171728 201454 172048 201486
rect 171728 201218 171770 201454
rect 172006 201218 172048 201454
rect 171728 201134 172048 201218
rect 171728 200898 171770 201134
rect 172006 200898 172048 201134
rect 171728 200866 172048 200898
rect 202448 201454 202768 201486
rect 202448 201218 202490 201454
rect 202726 201218 202768 201454
rect 202448 201134 202768 201218
rect 202448 200898 202490 201134
rect 202726 200898 202768 201134
rect 202448 200866 202768 200898
rect 64208 183454 64528 183486
rect 64208 183218 64250 183454
rect 64486 183218 64528 183454
rect 64208 183134 64528 183218
rect 64208 182898 64250 183134
rect 64486 182898 64528 183134
rect 64208 182866 64528 182898
rect 94928 183454 95248 183486
rect 94928 183218 94970 183454
rect 95206 183218 95248 183454
rect 94928 183134 95248 183218
rect 94928 182898 94970 183134
rect 95206 182898 95248 183134
rect 94928 182866 95248 182898
rect 125648 183454 125968 183486
rect 125648 183218 125690 183454
rect 125926 183218 125968 183454
rect 125648 183134 125968 183218
rect 125648 182898 125690 183134
rect 125926 182898 125968 183134
rect 125648 182866 125968 182898
rect 156368 183454 156688 183486
rect 156368 183218 156410 183454
rect 156646 183218 156688 183454
rect 156368 183134 156688 183218
rect 156368 182898 156410 183134
rect 156646 182898 156688 183134
rect 156368 182866 156688 182898
rect 187088 183454 187408 183486
rect 187088 183218 187130 183454
rect 187366 183218 187408 183454
rect 187088 183134 187408 183218
rect 187088 182898 187130 183134
rect 187366 182898 187408 183134
rect 187088 182866 187408 182898
rect 217808 183454 218128 183486
rect 217808 183218 217850 183454
rect 218086 183218 218128 183454
rect 217808 183134 218128 183218
rect 217808 182898 217850 183134
rect 218086 182898 218128 183134
rect 217808 182866 218128 182898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 79568 165454 79888 165486
rect 79568 165218 79610 165454
rect 79846 165218 79888 165454
rect 79568 165134 79888 165218
rect 79568 164898 79610 165134
rect 79846 164898 79888 165134
rect 79568 164866 79888 164898
rect 110288 165454 110608 165486
rect 110288 165218 110330 165454
rect 110566 165218 110608 165454
rect 110288 165134 110608 165218
rect 110288 164898 110330 165134
rect 110566 164898 110608 165134
rect 110288 164866 110608 164898
rect 141008 165454 141328 165486
rect 141008 165218 141050 165454
rect 141286 165218 141328 165454
rect 141008 165134 141328 165218
rect 141008 164898 141050 165134
rect 141286 164898 141328 165134
rect 141008 164866 141328 164898
rect 171728 165454 172048 165486
rect 171728 165218 171770 165454
rect 172006 165218 172048 165454
rect 171728 165134 172048 165218
rect 171728 164898 171770 165134
rect 172006 164898 172048 165134
rect 171728 164866 172048 164898
rect 202448 165454 202768 165486
rect 202448 165218 202490 165454
rect 202726 165218 202768 165454
rect 202448 165134 202768 165218
rect 202448 164898 202490 165134
rect 202726 164898 202768 165134
rect 202448 164866 202768 164898
rect 64208 147454 64528 147486
rect 64208 147218 64250 147454
rect 64486 147218 64528 147454
rect 64208 147134 64528 147218
rect 64208 146898 64250 147134
rect 64486 146898 64528 147134
rect 64208 146866 64528 146898
rect 94928 147454 95248 147486
rect 94928 147218 94970 147454
rect 95206 147218 95248 147454
rect 94928 147134 95248 147218
rect 94928 146898 94970 147134
rect 95206 146898 95248 147134
rect 94928 146866 95248 146898
rect 125648 147454 125968 147486
rect 125648 147218 125690 147454
rect 125926 147218 125968 147454
rect 125648 147134 125968 147218
rect 125648 146898 125690 147134
rect 125926 146898 125968 147134
rect 125648 146866 125968 146898
rect 156368 147454 156688 147486
rect 156368 147218 156410 147454
rect 156646 147218 156688 147454
rect 156368 147134 156688 147218
rect 156368 146898 156410 147134
rect 156646 146898 156688 147134
rect 156368 146866 156688 146898
rect 187088 147454 187408 147486
rect 187088 147218 187130 147454
rect 187366 147218 187408 147454
rect 187088 147134 187408 147218
rect 187088 146898 187130 147134
rect 187366 146898 187408 147134
rect 187088 146866 187408 146898
rect 217808 147454 218128 147486
rect 217808 147218 217850 147454
rect 218086 147218 218128 147454
rect 217808 147134 218128 147218
rect 217808 146898 217850 147134
rect 218086 146898 218128 147134
rect 217808 146866 218128 146898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 79568 129454 79888 129486
rect 79568 129218 79610 129454
rect 79846 129218 79888 129454
rect 79568 129134 79888 129218
rect 79568 128898 79610 129134
rect 79846 128898 79888 129134
rect 79568 128866 79888 128898
rect 110288 129454 110608 129486
rect 110288 129218 110330 129454
rect 110566 129218 110608 129454
rect 110288 129134 110608 129218
rect 110288 128898 110330 129134
rect 110566 128898 110608 129134
rect 110288 128866 110608 128898
rect 141008 129454 141328 129486
rect 141008 129218 141050 129454
rect 141286 129218 141328 129454
rect 141008 129134 141328 129218
rect 141008 128898 141050 129134
rect 141286 128898 141328 129134
rect 141008 128866 141328 128898
rect 171728 129454 172048 129486
rect 171728 129218 171770 129454
rect 172006 129218 172048 129454
rect 171728 129134 172048 129218
rect 171728 128898 171770 129134
rect 172006 128898 172048 129134
rect 171728 128866 172048 128898
rect 202448 129454 202768 129486
rect 202448 129218 202490 129454
rect 202726 129218 202768 129454
rect 202448 129134 202768 129218
rect 202448 128898 202490 129134
rect 202726 128898 202768 129134
rect 202448 128866 202768 128898
rect 64208 111454 64528 111486
rect 64208 111218 64250 111454
rect 64486 111218 64528 111454
rect 64208 111134 64528 111218
rect 64208 110898 64250 111134
rect 64486 110898 64528 111134
rect 64208 110866 64528 110898
rect 94928 111454 95248 111486
rect 94928 111218 94970 111454
rect 95206 111218 95248 111454
rect 94928 111134 95248 111218
rect 94928 110898 94970 111134
rect 95206 110898 95248 111134
rect 94928 110866 95248 110898
rect 125648 111454 125968 111486
rect 125648 111218 125690 111454
rect 125926 111218 125968 111454
rect 125648 111134 125968 111218
rect 125648 110898 125690 111134
rect 125926 110898 125968 111134
rect 125648 110866 125968 110898
rect 156368 111454 156688 111486
rect 156368 111218 156410 111454
rect 156646 111218 156688 111454
rect 156368 111134 156688 111218
rect 156368 110898 156410 111134
rect 156646 110898 156688 111134
rect 156368 110866 156688 110898
rect 187088 111454 187408 111486
rect 187088 111218 187130 111454
rect 187366 111218 187408 111454
rect 187088 111134 187408 111218
rect 187088 110898 187130 111134
rect 187366 110898 187408 111134
rect 187088 110866 187408 110898
rect 217808 111454 218128 111486
rect 217808 111218 217850 111454
rect 218086 111218 218128 111454
rect 217808 111134 218128 111218
rect 217808 110898 217850 111134
rect 218086 110898 218128 111134
rect 217808 110866 218128 110898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 79568 93454 79888 93486
rect 79568 93218 79610 93454
rect 79846 93218 79888 93454
rect 79568 93134 79888 93218
rect 79568 92898 79610 93134
rect 79846 92898 79888 93134
rect 79568 92866 79888 92898
rect 110288 93454 110608 93486
rect 110288 93218 110330 93454
rect 110566 93218 110608 93454
rect 110288 93134 110608 93218
rect 110288 92898 110330 93134
rect 110566 92898 110608 93134
rect 110288 92866 110608 92898
rect 141008 93454 141328 93486
rect 141008 93218 141050 93454
rect 141286 93218 141328 93454
rect 141008 93134 141328 93218
rect 141008 92898 141050 93134
rect 141286 92898 141328 93134
rect 141008 92866 141328 92898
rect 171728 93454 172048 93486
rect 171728 93218 171770 93454
rect 172006 93218 172048 93454
rect 171728 93134 172048 93218
rect 171728 92898 171770 93134
rect 172006 92898 172048 93134
rect 171728 92866 172048 92898
rect 202448 93454 202768 93486
rect 202448 93218 202490 93454
rect 202726 93218 202768 93454
rect 202448 93134 202768 93218
rect 202448 92898 202490 93134
rect 202726 92898 202768 93134
rect 202448 92866 202768 92898
rect 64208 75454 64528 75486
rect 64208 75218 64250 75454
rect 64486 75218 64528 75454
rect 64208 75134 64528 75218
rect 64208 74898 64250 75134
rect 64486 74898 64528 75134
rect 64208 74866 64528 74898
rect 94928 75454 95248 75486
rect 94928 75218 94970 75454
rect 95206 75218 95248 75454
rect 94928 75134 95248 75218
rect 94928 74898 94970 75134
rect 95206 74898 95248 75134
rect 94928 74866 95248 74898
rect 125648 75454 125968 75486
rect 125648 75218 125690 75454
rect 125926 75218 125968 75454
rect 125648 75134 125968 75218
rect 125648 74898 125690 75134
rect 125926 74898 125968 75134
rect 125648 74866 125968 74898
rect 156368 75454 156688 75486
rect 156368 75218 156410 75454
rect 156646 75218 156688 75454
rect 156368 75134 156688 75218
rect 156368 74898 156410 75134
rect 156646 74898 156688 75134
rect 156368 74866 156688 74898
rect 187088 75454 187408 75486
rect 187088 75218 187130 75454
rect 187366 75218 187408 75454
rect 187088 75134 187408 75218
rect 187088 74898 187130 75134
rect 187366 74898 187408 75134
rect 187088 74866 187408 74898
rect 217808 75454 218128 75486
rect 217808 75218 217850 75454
rect 218086 75218 218128 75454
rect 217808 75134 218128 75218
rect 217808 74898 217850 75134
rect 218086 74898 218128 75134
rect 217808 74866 218128 74898
rect 60595 63612 60661 63613
rect 60595 63548 60596 63612
rect 60660 63548 60661 63612
rect 60595 63547 60661 63548
rect 60598 60349 60658 63547
rect 60595 60348 60661 60349
rect 60595 60284 60596 60348
rect 60660 60284 60661 60348
rect 60595 60283 60661 60284
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -1306 56414 20898
rect 55794 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 56414 -1306
rect 55794 -1626 56414 -1542
rect 55794 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 56414 -1626
rect 55794 -1894 56414 -1862
rect 59514 25174 60134 58000
rect 59514 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 60134 25174
rect 59514 24854 60134 24938
rect 59514 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 60134 24854
rect 59514 -3226 60134 24618
rect 59514 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 60134 -3226
rect 59514 -3546 60134 -3462
rect 59514 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 60134 -3546
rect 59514 -3814 60134 -3782
rect 63234 28894 63854 58000
rect 63234 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 63854 28894
rect 63234 28574 63854 28658
rect 63234 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 63854 28574
rect 63234 -5146 63854 28338
rect 63234 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 63854 -5146
rect 63234 -5466 63854 -5382
rect 63234 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 63854 -5466
rect 63234 -5734 63854 -5702
rect 66954 32614 67574 58000
rect 66954 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 67574 32614
rect 66954 32294 67574 32378
rect 66954 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 67574 32294
rect 48954 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 49574 -6106
rect 48954 -6426 49574 -6342
rect 48954 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 49574 -6426
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 32058
rect 73794 39454 74414 58000
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 77514 43174 78134 58000
rect 77514 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 78134 43174
rect 77514 42854 78134 42938
rect 77514 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 78134 42854
rect 77514 7174 78134 42618
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -2266 78134 6618
rect 77514 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 78134 -2266
rect 77514 -2586 78134 -2502
rect 77514 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 78134 -2586
rect 77514 -3814 78134 -2822
rect 81234 46894 81854 58000
rect 81234 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 81854 46894
rect 81234 46574 81854 46658
rect 81234 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 81854 46574
rect 81234 10894 81854 46338
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -4186 81854 10338
rect 81234 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 81854 -4186
rect 81234 -4506 81854 -4422
rect 81234 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 81854 -4506
rect 81234 -5734 81854 -4742
rect 84954 50614 85574 58000
rect 84954 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 85574 50614
rect 84954 50294 85574 50378
rect 84954 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 85574 50294
rect 84954 14614 85574 50058
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 66954 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 67574 -7066
rect 66954 -7386 67574 -7302
rect 66954 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 67574 -7386
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 14058
rect 91794 57454 92414 58000
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -1306 92414 20898
rect 91794 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 92414 -1306
rect 91794 -1626 92414 -1542
rect 91794 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 92414 -1626
rect 91794 -1894 92414 -1862
rect 95514 25174 96134 58000
rect 95514 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 96134 25174
rect 95514 24854 96134 24938
rect 95514 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 96134 24854
rect 95514 -3226 96134 24618
rect 95514 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 96134 -3226
rect 95514 -3546 96134 -3462
rect 95514 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 96134 -3546
rect 95514 -3814 96134 -3782
rect 99234 28894 99854 58000
rect 99234 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 99854 28894
rect 99234 28574 99854 28658
rect 99234 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 99854 28574
rect 99234 -5146 99854 28338
rect 99234 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 99854 -5146
rect 99234 -5466 99854 -5382
rect 99234 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 99854 -5466
rect 99234 -5734 99854 -5702
rect 102954 32614 103574 58000
rect 102954 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 103574 32614
rect 102954 32294 103574 32378
rect 102954 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 103574 32294
rect 84954 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 85574 -6106
rect 84954 -6426 85574 -6342
rect 84954 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 85574 -6426
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 32058
rect 109794 39454 110414 58000
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 113514 43174 114134 58000
rect 113514 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 114134 43174
rect 113514 42854 114134 42938
rect 113514 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 114134 42854
rect 113514 7174 114134 42618
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -2266 114134 6618
rect 113514 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 114134 -2266
rect 113514 -2586 114134 -2502
rect 113514 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 114134 -2586
rect 113514 -3814 114134 -2822
rect 117234 46894 117854 58000
rect 117234 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 117854 46894
rect 117234 46574 117854 46658
rect 117234 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 117854 46574
rect 117234 10894 117854 46338
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -4186 117854 10338
rect 117234 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 117854 -4186
rect 117234 -4506 117854 -4422
rect 117234 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 117854 -4506
rect 117234 -5734 117854 -4742
rect 120954 50614 121574 58000
rect 120954 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 121574 50614
rect 120954 50294 121574 50378
rect 120954 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 121574 50294
rect 120954 14614 121574 50058
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 102954 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 103574 -7066
rect 102954 -7386 103574 -7302
rect 102954 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 103574 -7386
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 14058
rect 127794 57454 128414 58000
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -1306 128414 20898
rect 127794 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 128414 -1306
rect 127794 -1626 128414 -1542
rect 127794 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 128414 -1626
rect 127794 -1894 128414 -1862
rect 131514 25174 132134 58000
rect 131514 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 132134 25174
rect 131514 24854 132134 24938
rect 131514 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 132134 24854
rect 131514 -3226 132134 24618
rect 131514 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 132134 -3226
rect 131514 -3546 132134 -3462
rect 131514 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 132134 -3546
rect 131514 -3814 132134 -3782
rect 135234 28894 135854 58000
rect 135234 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 135854 28894
rect 135234 28574 135854 28658
rect 135234 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 135854 28574
rect 135234 -5146 135854 28338
rect 135234 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 135854 -5146
rect 135234 -5466 135854 -5382
rect 135234 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 135854 -5466
rect 135234 -5734 135854 -5702
rect 138954 32614 139574 58000
rect 138954 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 139574 32614
rect 138954 32294 139574 32378
rect 138954 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 139574 32294
rect 120954 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 121574 -6106
rect 120954 -6426 121574 -6342
rect 120954 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 121574 -6426
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 32058
rect 145794 39454 146414 58000
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 149514 43174 150134 58000
rect 149514 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 150134 43174
rect 149514 42854 150134 42938
rect 149514 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 150134 42854
rect 149514 7174 150134 42618
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -2266 150134 6618
rect 149514 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 150134 -2266
rect 149514 -2586 150134 -2502
rect 149514 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 150134 -2586
rect 149514 -3814 150134 -2822
rect 153234 46894 153854 58000
rect 153234 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 153854 46894
rect 153234 46574 153854 46658
rect 153234 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 153854 46574
rect 153234 10894 153854 46338
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -4186 153854 10338
rect 153234 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 153854 -4186
rect 153234 -4506 153854 -4422
rect 153234 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 153854 -4506
rect 153234 -5734 153854 -4742
rect 156954 50614 157574 58000
rect 156954 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 157574 50614
rect 156954 50294 157574 50378
rect 156954 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 157574 50294
rect 156954 14614 157574 50058
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 138954 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 139574 -7066
rect 138954 -7386 139574 -7302
rect 138954 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 139574 -7386
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 14058
rect 163794 57454 164414 58000
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -1306 164414 20898
rect 163794 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 164414 -1306
rect 163794 -1626 164414 -1542
rect 163794 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 164414 -1626
rect 163794 -1894 164414 -1862
rect 167514 25174 168134 58000
rect 167514 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 168134 25174
rect 167514 24854 168134 24938
rect 167514 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 168134 24854
rect 167514 -3226 168134 24618
rect 167514 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 168134 -3226
rect 167514 -3546 168134 -3462
rect 167514 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 168134 -3546
rect 167514 -3814 168134 -3782
rect 171234 28894 171854 58000
rect 171234 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 171854 28894
rect 171234 28574 171854 28658
rect 171234 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 171854 28574
rect 171234 -5146 171854 28338
rect 171234 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 171854 -5146
rect 171234 -5466 171854 -5382
rect 171234 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 171854 -5466
rect 171234 -5734 171854 -5702
rect 174954 32614 175574 58000
rect 174954 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 175574 32614
rect 174954 32294 175574 32378
rect 174954 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 175574 32294
rect 156954 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 157574 -6106
rect 156954 -6426 157574 -6342
rect 156954 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 157574 -6426
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 32058
rect 181794 39454 182414 58000
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 185514 43174 186134 58000
rect 185514 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 186134 43174
rect 185514 42854 186134 42938
rect 185514 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 186134 42854
rect 185514 7174 186134 42618
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -2266 186134 6618
rect 185514 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 186134 -2266
rect 185514 -2586 186134 -2502
rect 185514 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 186134 -2586
rect 185514 -3814 186134 -2822
rect 189234 46894 189854 58000
rect 189234 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 189854 46894
rect 189234 46574 189854 46658
rect 189234 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 189854 46574
rect 189234 10894 189854 46338
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -4186 189854 10338
rect 189234 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 189854 -4186
rect 189234 -4506 189854 -4422
rect 189234 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 189854 -4506
rect 189234 -5734 189854 -4742
rect 192954 50614 193574 58000
rect 192954 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 193574 50614
rect 192954 50294 193574 50378
rect 192954 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 193574 50294
rect 192954 14614 193574 50058
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 174954 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 175574 -7066
rect 174954 -7386 175574 -7302
rect 174954 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 175574 -7386
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 14058
rect 199794 57454 200414 58000
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -1306 200414 20898
rect 199794 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 200414 -1306
rect 199794 -1626 200414 -1542
rect 199794 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 200414 -1626
rect 199794 -1894 200414 -1862
rect 203514 25174 204134 58000
rect 203514 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 204134 25174
rect 203514 24854 204134 24938
rect 203514 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 204134 24854
rect 203514 -3226 204134 24618
rect 203514 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 204134 -3226
rect 203514 -3546 204134 -3462
rect 203514 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 204134 -3546
rect 203514 -3814 204134 -3782
rect 207234 28894 207854 58000
rect 207234 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 207854 28894
rect 207234 28574 207854 28658
rect 207234 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 207854 28574
rect 207234 -5146 207854 28338
rect 207234 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 207854 -5146
rect 207234 -5466 207854 -5382
rect 207234 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 207854 -5466
rect 207234 -5734 207854 -5702
rect 210954 32614 211574 58000
rect 210954 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 211574 32614
rect 210954 32294 211574 32378
rect 210954 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 211574 32294
rect 192954 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 193574 -6106
rect 192954 -6426 193574 -6342
rect 192954 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 193574 -6426
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 32058
rect 217794 39454 218414 58000
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 221514 43174 222134 58000
rect 224910 57493 224970 229470
rect 224907 57492 224973 57493
rect 224907 57428 224908 57492
rect 224972 57428 224973 57492
rect 224907 57427 224973 57428
rect 224907 56948 224973 56949
rect 224907 56884 224908 56948
rect 224972 56884 224973 56948
rect 224907 56883 224973 56884
rect 224910 56810 224970 56883
rect 225094 56810 225154 230150
rect 225234 228675 225854 262338
rect 226011 227492 226077 227493
rect 226011 227428 226012 227492
rect 226076 227428 226077 227492
rect 226011 227427 226077 227428
rect 224910 56750 225154 56810
rect 221514 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 222134 43174
rect 221514 42854 222134 42938
rect 221514 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 222134 42854
rect 221514 7174 222134 42618
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -2266 222134 6618
rect 221514 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 222134 -2266
rect 221514 -2586 222134 -2502
rect 221514 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 222134 -2586
rect 221514 -3814 222134 -2822
rect 225234 46894 225854 58000
rect 226014 57357 226074 227427
rect 226382 85373 226442 397971
rect 228954 374614 229574 398000
rect 228954 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 229574 374614
rect 228954 374294 229574 374378
rect 228954 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 229574 374294
rect 228954 338614 229574 374058
rect 228954 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 229574 338614
rect 228954 338294 229574 338378
rect 228954 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 229574 338294
rect 228954 302614 229574 338058
rect 228954 302378 228986 302614
rect 229222 302378 229306 302614
rect 229542 302378 229574 302614
rect 228954 302294 229574 302378
rect 228954 302058 228986 302294
rect 229222 302058 229306 302294
rect 229542 302058 229574 302294
rect 228954 266614 229574 302058
rect 228954 266378 228986 266614
rect 229222 266378 229306 266614
rect 229542 266378 229574 266614
rect 228954 266294 229574 266378
rect 228954 266058 228986 266294
rect 229222 266058 229306 266294
rect 229542 266058 229574 266294
rect 226747 242180 226813 242181
rect 226747 242116 226748 242180
rect 226812 242116 226813 242180
rect 226747 242115 226813 242116
rect 226563 227900 226629 227901
rect 226563 227836 226564 227900
rect 226628 227836 226629 227900
rect 226563 227835 226629 227836
rect 226379 85372 226445 85373
rect 226379 85308 226380 85372
rect 226444 85308 226445 85372
rect 226379 85307 226445 85308
rect 226566 69325 226626 227835
rect 226750 115021 226810 242115
rect 228403 236060 228469 236061
rect 228403 235996 228404 236060
rect 228468 235996 228469 236060
rect 228403 235995 228469 235996
rect 228219 233340 228285 233341
rect 228219 233276 228220 233340
rect 228284 233276 228285 233340
rect 228219 233275 228285 233276
rect 226931 232524 226997 232525
rect 226931 232460 226932 232524
rect 226996 232460 226997 232524
rect 226931 232459 226997 232460
rect 226747 115020 226813 115021
rect 226747 114956 226748 115020
rect 226812 114956 226813 115020
rect 226747 114955 226813 114956
rect 226934 106997 226994 232459
rect 227299 220964 227365 220965
rect 227299 220900 227300 220964
rect 227364 220900 227365 220964
rect 227299 220899 227365 220900
rect 227302 219605 227362 220899
rect 227299 219604 227365 219605
rect 227299 219540 227300 219604
rect 227364 219540 227365 219604
rect 227299 219539 227365 219540
rect 228222 111893 228282 233275
rect 228406 218109 228466 235995
rect 228954 230614 229574 266058
rect 228954 230378 228986 230614
rect 229222 230378 229306 230614
rect 229542 230378 229574 230614
rect 228954 230294 229574 230378
rect 228954 230058 228986 230294
rect 229222 230058 229306 230294
rect 229542 230058 229574 230294
rect 228403 218108 228469 218109
rect 228403 218044 228404 218108
rect 228468 218044 228469 218108
rect 228403 218043 228469 218044
rect 228954 194614 229574 230058
rect 228954 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 229574 194614
rect 228954 194294 229574 194378
rect 228954 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 229574 194294
rect 228954 158614 229574 194058
rect 228954 158378 228986 158614
rect 229222 158378 229306 158614
rect 229542 158378 229574 158614
rect 228954 158294 229574 158378
rect 228954 158058 228986 158294
rect 229222 158058 229306 158294
rect 229542 158058 229574 158294
rect 228954 122614 229574 158058
rect 228954 122378 228986 122614
rect 229222 122378 229306 122614
rect 229542 122378 229574 122614
rect 228954 122294 229574 122378
rect 228954 122058 228986 122294
rect 229222 122058 229306 122294
rect 229542 122058 229574 122294
rect 228219 111892 228285 111893
rect 228219 111828 228220 111892
rect 228284 111828 228285 111892
rect 228219 111827 228285 111828
rect 226931 106996 226997 106997
rect 226931 106932 226932 106996
rect 226996 106932 226997 106996
rect 226931 106931 226997 106932
rect 228954 86614 229574 122058
rect 228954 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 229574 86614
rect 228954 86294 229574 86378
rect 228954 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 229574 86294
rect 226563 69324 226629 69325
rect 226563 69260 226564 69324
rect 226628 69260 226629 69324
rect 226563 69259 226629 69260
rect 226011 57356 226077 57357
rect 226011 57292 226012 57356
rect 226076 57292 226077 57356
rect 226011 57291 226077 57292
rect 225234 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 225854 46894
rect 225234 46574 225854 46658
rect 225234 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 225854 46574
rect 225234 10894 225854 46338
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -4186 225854 10338
rect 225234 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 225854 -4186
rect 225234 -4506 225854 -4422
rect 225234 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 225854 -4506
rect 225234 -5734 225854 -4742
rect 228954 50614 229574 86058
rect 228954 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 229574 50614
rect 228954 50294 229574 50378
rect 228954 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 229574 50294
rect 228954 14614 229574 50058
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 210954 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 211574 -7066
rect 210954 -7386 211574 -7302
rect 210954 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 211574 -7386
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 14058
rect 235794 381454 236414 398000
rect 237054 397357 237114 399470
rect 238158 397357 238218 399470
rect 239262 397357 239322 399470
rect 237051 397356 237117 397357
rect 237051 397292 237052 397356
rect 237116 397292 237117 397356
rect 237051 397291 237117 397292
rect 238155 397356 238221 397357
rect 238155 397292 238156 397356
rect 238220 397292 238221 397356
rect 238155 397291 238221 397292
rect 239259 397356 239325 397357
rect 239259 397292 239260 397356
rect 239324 397292 239325 397356
rect 239259 397291 239325 397292
rect 235794 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 236414 381454
rect 235794 381134 236414 381218
rect 235794 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 236414 381134
rect 235794 345454 236414 380898
rect 235794 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 236414 345454
rect 235794 345134 236414 345218
rect 235794 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 236414 345134
rect 235794 309454 236414 344898
rect 235794 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 236414 309454
rect 235794 309134 236414 309218
rect 235794 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 236414 309134
rect 235794 273454 236414 308898
rect 235794 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 236414 273454
rect 235794 273134 236414 273218
rect 235794 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 236414 273134
rect 235794 237454 236414 272898
rect 235794 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 236414 237454
rect 235794 237134 236414 237218
rect 235794 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 236414 237134
rect 235794 201454 236414 236898
rect 235794 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 236414 201454
rect 235794 201134 236414 201218
rect 235794 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 236414 201134
rect 235794 165454 236414 200898
rect 235794 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 236414 165454
rect 235794 165134 236414 165218
rect 235794 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 236414 165134
rect 235794 129454 236414 164898
rect 235794 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 236414 129454
rect 235794 129134 236414 129218
rect 235794 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 236414 129134
rect 235794 93454 236414 128898
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -1306 236414 20898
rect 235794 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 236414 -1306
rect 235794 -1626 236414 -1542
rect 235794 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 236414 -1626
rect 235794 -1894 236414 -1862
rect 239514 385174 240134 398000
rect 240550 397357 240610 399470
rect 241654 399470 241828 399530
rect 242942 399470 243188 399530
rect 244216 399530 244276 400106
rect 245440 399530 245500 400106
rect 246528 399530 246588 400106
rect 244216 399470 244290 399530
rect 241654 397357 241714 399470
rect 240547 397356 240613 397357
rect 240547 397292 240548 397356
rect 240612 397292 240613 397356
rect 240547 397291 240613 397292
rect 241651 397356 241717 397357
rect 241651 397292 241652 397356
rect 241716 397292 241717 397356
rect 241651 397291 241717 397292
rect 242942 396813 243002 399470
rect 242939 396812 243005 396813
rect 242939 396748 242940 396812
rect 243004 396748 243005 396812
rect 242939 396747 243005 396748
rect 239514 384938 239546 385174
rect 239782 384938 239866 385174
rect 240102 384938 240134 385174
rect 239514 384854 240134 384938
rect 239514 384618 239546 384854
rect 239782 384618 239866 384854
rect 240102 384618 240134 384854
rect 239514 349174 240134 384618
rect 239514 348938 239546 349174
rect 239782 348938 239866 349174
rect 240102 348938 240134 349174
rect 239514 348854 240134 348938
rect 239514 348618 239546 348854
rect 239782 348618 239866 348854
rect 240102 348618 240134 348854
rect 239514 313174 240134 348618
rect 239514 312938 239546 313174
rect 239782 312938 239866 313174
rect 240102 312938 240134 313174
rect 239514 312854 240134 312938
rect 239514 312618 239546 312854
rect 239782 312618 239866 312854
rect 240102 312618 240134 312854
rect 239514 277174 240134 312618
rect 239514 276938 239546 277174
rect 239782 276938 239866 277174
rect 240102 276938 240134 277174
rect 239514 276854 240134 276938
rect 239514 276618 239546 276854
rect 239782 276618 239866 276854
rect 240102 276618 240134 276854
rect 239514 241174 240134 276618
rect 239514 240938 239546 241174
rect 239782 240938 239866 241174
rect 240102 240938 240134 241174
rect 239514 240854 240134 240938
rect 239514 240618 239546 240854
rect 239782 240618 239866 240854
rect 240102 240618 240134 240854
rect 239514 205174 240134 240618
rect 239514 204938 239546 205174
rect 239782 204938 239866 205174
rect 240102 204938 240134 205174
rect 239514 204854 240134 204938
rect 239514 204618 239546 204854
rect 239782 204618 239866 204854
rect 240102 204618 240134 204854
rect 239514 169174 240134 204618
rect 239514 168938 239546 169174
rect 239782 168938 239866 169174
rect 240102 168938 240134 169174
rect 239514 168854 240134 168938
rect 239514 168618 239546 168854
rect 239782 168618 239866 168854
rect 240102 168618 240134 168854
rect 239514 133174 240134 168618
rect 239514 132938 239546 133174
rect 239782 132938 239866 133174
rect 240102 132938 240134 133174
rect 239514 132854 240134 132938
rect 239514 132618 239546 132854
rect 239782 132618 239866 132854
rect 240102 132618 240134 132854
rect 239514 97174 240134 132618
rect 239514 96938 239546 97174
rect 239782 96938 239866 97174
rect 240102 96938 240134 97174
rect 239514 96854 240134 96938
rect 239514 96618 239546 96854
rect 239782 96618 239866 96854
rect 240102 96618 240134 96854
rect 239514 61174 240134 96618
rect 239514 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 240134 61174
rect 239514 60854 240134 60938
rect 239514 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 240134 60854
rect 239514 25174 240134 60618
rect 239514 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 240134 25174
rect 239514 24854 240134 24938
rect 239514 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 240134 24854
rect 239514 -3226 240134 24618
rect 239514 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 240134 -3226
rect 239514 -3546 240134 -3462
rect 239514 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 240134 -3546
rect 239514 -3814 240134 -3782
rect 243234 388894 243854 398000
rect 244230 396813 244290 399470
rect 245334 399470 245500 399530
rect 246438 399470 246588 399530
rect 247616 399530 247676 400106
rect 248296 399530 248356 400106
rect 248704 399530 248764 400106
rect 247616 399470 247786 399530
rect 244227 396812 244293 396813
rect 244227 396748 244228 396812
rect 244292 396748 244293 396812
rect 244227 396747 244293 396748
rect 245334 396677 245394 399470
rect 246438 396813 246498 399470
rect 246435 396812 246501 396813
rect 246435 396748 246436 396812
rect 246500 396748 246501 396812
rect 246435 396747 246501 396748
rect 245331 396676 245397 396677
rect 245331 396612 245332 396676
rect 245396 396612 245397 396676
rect 245331 396611 245397 396612
rect 243234 388658 243266 388894
rect 243502 388658 243586 388894
rect 243822 388658 243854 388894
rect 243234 388574 243854 388658
rect 243234 388338 243266 388574
rect 243502 388338 243586 388574
rect 243822 388338 243854 388574
rect 243234 352894 243854 388338
rect 243234 352658 243266 352894
rect 243502 352658 243586 352894
rect 243822 352658 243854 352894
rect 243234 352574 243854 352658
rect 243234 352338 243266 352574
rect 243502 352338 243586 352574
rect 243822 352338 243854 352574
rect 243234 316894 243854 352338
rect 243234 316658 243266 316894
rect 243502 316658 243586 316894
rect 243822 316658 243854 316894
rect 243234 316574 243854 316658
rect 243234 316338 243266 316574
rect 243502 316338 243586 316574
rect 243822 316338 243854 316574
rect 243234 280894 243854 316338
rect 243234 280658 243266 280894
rect 243502 280658 243586 280894
rect 243822 280658 243854 280894
rect 243234 280574 243854 280658
rect 243234 280338 243266 280574
rect 243502 280338 243586 280574
rect 243822 280338 243854 280574
rect 243234 244894 243854 280338
rect 243234 244658 243266 244894
rect 243502 244658 243586 244894
rect 243822 244658 243854 244894
rect 243234 244574 243854 244658
rect 243234 244338 243266 244574
rect 243502 244338 243586 244574
rect 243822 244338 243854 244574
rect 243234 208894 243854 244338
rect 243234 208658 243266 208894
rect 243502 208658 243586 208894
rect 243822 208658 243854 208894
rect 243234 208574 243854 208658
rect 243234 208338 243266 208574
rect 243502 208338 243586 208574
rect 243822 208338 243854 208574
rect 243234 172894 243854 208338
rect 243234 172658 243266 172894
rect 243502 172658 243586 172894
rect 243822 172658 243854 172894
rect 243234 172574 243854 172658
rect 243234 172338 243266 172574
rect 243502 172338 243586 172574
rect 243822 172338 243854 172574
rect 243234 136894 243854 172338
rect 243234 136658 243266 136894
rect 243502 136658 243586 136894
rect 243822 136658 243854 136894
rect 243234 136574 243854 136658
rect 243234 136338 243266 136574
rect 243502 136338 243586 136574
rect 243822 136338 243854 136574
rect 243234 100894 243854 136338
rect 243234 100658 243266 100894
rect 243502 100658 243586 100894
rect 243822 100658 243854 100894
rect 243234 100574 243854 100658
rect 243234 100338 243266 100574
rect 243502 100338 243586 100574
rect 243822 100338 243854 100574
rect 243234 64894 243854 100338
rect 243234 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 243854 64894
rect 243234 64574 243854 64658
rect 243234 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 243854 64574
rect 243234 28894 243854 64338
rect 243234 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 243854 28894
rect 243234 28574 243854 28658
rect 243234 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 243854 28574
rect 243234 -5146 243854 28338
rect 243234 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 243854 -5146
rect 243234 -5466 243854 -5382
rect 243234 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 243854 -5466
rect 243234 -5734 243854 -5702
rect 246954 392614 247574 398000
rect 247726 397357 247786 399470
rect 248278 399470 248356 399530
rect 248646 399470 248764 399530
rect 250064 399530 250124 400106
rect 250744 399530 250804 400106
rect 251288 399530 251348 400106
rect 252376 399530 252436 400106
rect 253464 399530 253524 400106
rect 250064 399470 250178 399530
rect 247723 397356 247789 397357
rect 247723 397292 247724 397356
rect 247788 397292 247789 397356
rect 247723 397291 247789 397292
rect 248278 396813 248338 399470
rect 248646 396813 248706 399470
rect 250118 396813 250178 399470
rect 250670 399470 250804 399530
rect 251222 399470 251348 399530
rect 252326 399470 252436 399530
rect 253430 399470 253524 399530
rect 253600 399530 253660 400106
rect 254552 399530 254612 400106
rect 255912 399530 255972 400106
rect 253600 399470 253674 399530
rect 250670 397357 250730 399470
rect 250667 397356 250733 397357
rect 250667 397292 250668 397356
rect 250732 397292 250733 397356
rect 250667 397291 250733 397292
rect 251222 397221 251282 399470
rect 252326 397357 252386 399470
rect 253430 397357 253490 399470
rect 252323 397356 252389 397357
rect 252323 397292 252324 397356
rect 252388 397292 252389 397356
rect 252323 397291 252389 397292
rect 253427 397356 253493 397357
rect 253427 397292 253428 397356
rect 253492 397292 253493 397356
rect 253427 397291 253493 397292
rect 251219 397220 251285 397221
rect 251219 397156 251220 397220
rect 251284 397156 251285 397220
rect 251219 397155 251285 397156
rect 253614 396813 253674 399470
rect 254534 399470 254612 399530
rect 255822 399470 255972 399530
rect 256048 399530 256108 400106
rect 257000 399530 257060 400106
rect 256048 399470 256250 399530
rect 248275 396812 248341 396813
rect 248275 396748 248276 396812
rect 248340 396748 248341 396812
rect 248275 396747 248341 396748
rect 248643 396812 248709 396813
rect 248643 396748 248644 396812
rect 248708 396748 248709 396812
rect 248643 396747 248709 396748
rect 250115 396812 250181 396813
rect 250115 396748 250116 396812
rect 250180 396748 250181 396812
rect 250115 396747 250181 396748
rect 253611 396812 253677 396813
rect 253611 396748 253612 396812
rect 253676 396748 253677 396812
rect 253611 396747 253677 396748
rect 246954 392378 246986 392614
rect 247222 392378 247306 392614
rect 247542 392378 247574 392614
rect 246954 392294 247574 392378
rect 246954 392058 246986 392294
rect 247222 392058 247306 392294
rect 247542 392058 247574 392294
rect 246954 356614 247574 392058
rect 246954 356378 246986 356614
rect 247222 356378 247306 356614
rect 247542 356378 247574 356614
rect 246954 356294 247574 356378
rect 246954 356058 246986 356294
rect 247222 356058 247306 356294
rect 247542 356058 247574 356294
rect 246954 320614 247574 356058
rect 246954 320378 246986 320614
rect 247222 320378 247306 320614
rect 247542 320378 247574 320614
rect 246954 320294 247574 320378
rect 246954 320058 246986 320294
rect 247222 320058 247306 320294
rect 247542 320058 247574 320294
rect 246954 284614 247574 320058
rect 246954 284378 246986 284614
rect 247222 284378 247306 284614
rect 247542 284378 247574 284614
rect 246954 284294 247574 284378
rect 246954 284058 246986 284294
rect 247222 284058 247306 284294
rect 247542 284058 247574 284294
rect 246954 248614 247574 284058
rect 246954 248378 246986 248614
rect 247222 248378 247306 248614
rect 247542 248378 247574 248614
rect 246954 248294 247574 248378
rect 246954 248058 246986 248294
rect 247222 248058 247306 248294
rect 247542 248058 247574 248294
rect 246954 212614 247574 248058
rect 246954 212378 246986 212614
rect 247222 212378 247306 212614
rect 247542 212378 247574 212614
rect 246954 212294 247574 212378
rect 246954 212058 246986 212294
rect 247222 212058 247306 212294
rect 247542 212058 247574 212294
rect 246954 176614 247574 212058
rect 246954 176378 246986 176614
rect 247222 176378 247306 176614
rect 247542 176378 247574 176614
rect 246954 176294 247574 176378
rect 246954 176058 246986 176294
rect 247222 176058 247306 176294
rect 247542 176058 247574 176294
rect 246954 140614 247574 176058
rect 246954 140378 246986 140614
rect 247222 140378 247306 140614
rect 247542 140378 247574 140614
rect 246954 140294 247574 140378
rect 246954 140058 246986 140294
rect 247222 140058 247306 140294
rect 247542 140058 247574 140294
rect 246954 104614 247574 140058
rect 246954 104378 246986 104614
rect 247222 104378 247306 104614
rect 247542 104378 247574 104614
rect 246954 104294 247574 104378
rect 246954 104058 246986 104294
rect 247222 104058 247306 104294
rect 247542 104058 247574 104294
rect 246954 68614 247574 104058
rect 246954 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 247574 68614
rect 246954 68294 247574 68378
rect 246954 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 247574 68294
rect 246954 32614 247574 68058
rect 246954 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 247574 32614
rect 246954 32294 247574 32378
rect 246954 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 247574 32294
rect 228954 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 229574 -6106
rect 228954 -6426 229574 -6342
rect 228954 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 229574 -6426
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 32058
rect 253794 363454 254414 398000
rect 254534 396813 254594 399470
rect 255822 396813 255882 399470
rect 254531 396812 254597 396813
rect 254531 396748 254532 396812
rect 254596 396748 254597 396812
rect 254531 396747 254597 396748
rect 255819 396812 255885 396813
rect 255819 396748 255820 396812
rect 255884 396748 255885 396812
rect 255819 396747 255885 396748
rect 256190 396677 256250 399470
rect 256926 399470 257060 399530
rect 258088 399530 258148 400106
rect 258496 399530 258556 400106
rect 258088 399470 258274 399530
rect 256926 396813 256986 399470
rect 256923 396812 256989 396813
rect 256923 396748 256924 396812
rect 256988 396748 256989 396812
rect 256923 396747 256989 396748
rect 256187 396676 256253 396677
rect 256187 396612 256188 396676
rect 256252 396612 256253 396676
rect 256187 396611 256253 396612
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 253794 327454 254414 362898
rect 253794 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 254414 327454
rect 253794 327134 254414 327218
rect 253794 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 254414 327134
rect 253794 291454 254414 326898
rect 253794 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 254414 291454
rect 253794 291134 254414 291218
rect 253794 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 254414 291134
rect 253794 255454 254414 290898
rect 253794 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 254414 255454
rect 253794 255134 254414 255218
rect 253794 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 254414 255134
rect 253794 219454 254414 254898
rect 253794 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 254414 219454
rect 253794 219134 254414 219218
rect 253794 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 254414 219134
rect 253794 183454 254414 218898
rect 253794 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 254414 183454
rect 253794 183134 254414 183218
rect 253794 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 254414 183134
rect 253794 147454 254414 182898
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 253794 111454 254414 146898
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 257514 367174 258134 398000
rect 258214 396810 258274 399470
rect 258398 399470 258556 399530
rect 259448 399530 259508 400106
rect 260672 399530 260732 400106
rect 261080 399530 261140 400106
rect 259448 399470 259562 399530
rect 258398 396949 258458 399470
rect 258395 396948 258461 396949
rect 258395 396884 258396 396948
rect 258460 396884 258461 396948
rect 258395 396883 258461 396884
rect 259502 396813 259562 399470
rect 260606 399470 260732 399530
rect 260974 399470 261140 399530
rect 261760 399530 261820 400106
rect 262848 399530 262908 400106
rect 261760 399470 262138 399530
rect 260606 397357 260666 399470
rect 260603 397356 260669 397357
rect 260603 397292 260604 397356
rect 260668 397292 260669 397356
rect 260603 397291 260669 397292
rect 260974 396813 261034 399470
rect 258395 396812 258461 396813
rect 258395 396810 258396 396812
rect 258214 396750 258396 396810
rect 258395 396748 258396 396750
rect 258460 396748 258461 396812
rect 258395 396747 258461 396748
rect 259499 396812 259565 396813
rect 259499 396748 259500 396812
rect 259564 396748 259565 396812
rect 259499 396747 259565 396748
rect 260971 396812 261037 396813
rect 260971 396748 260972 396812
rect 261036 396748 261037 396812
rect 260971 396747 261037 396748
rect 257514 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 258134 367174
rect 257514 366854 258134 366938
rect 257514 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 258134 366854
rect 257514 331174 258134 366618
rect 257514 330938 257546 331174
rect 257782 330938 257866 331174
rect 258102 330938 258134 331174
rect 257514 330854 258134 330938
rect 257514 330618 257546 330854
rect 257782 330618 257866 330854
rect 258102 330618 258134 330854
rect 257514 295174 258134 330618
rect 257514 294938 257546 295174
rect 257782 294938 257866 295174
rect 258102 294938 258134 295174
rect 257514 294854 258134 294938
rect 257514 294618 257546 294854
rect 257782 294618 257866 294854
rect 258102 294618 258134 294854
rect 257514 259174 258134 294618
rect 257514 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 258134 259174
rect 257514 258854 258134 258938
rect 257514 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 258134 258854
rect 257514 223174 258134 258618
rect 257514 222938 257546 223174
rect 257782 222938 257866 223174
rect 258102 222938 258134 223174
rect 257514 222854 258134 222938
rect 257514 222618 257546 222854
rect 257782 222618 257866 222854
rect 258102 222618 258134 222854
rect 257514 187174 258134 222618
rect 257514 186938 257546 187174
rect 257782 186938 257866 187174
rect 258102 186938 258134 187174
rect 257514 186854 258134 186938
rect 257514 186618 257546 186854
rect 257782 186618 257866 186854
rect 258102 186618 258134 186854
rect 257514 151174 258134 186618
rect 257514 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 258134 151174
rect 257514 150854 258134 150938
rect 257514 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 258134 150854
rect 257514 115174 258134 150618
rect 257514 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 258134 115174
rect 257514 114854 258134 114938
rect 257514 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 258134 114854
rect 257514 79174 258134 114618
rect 257514 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 258134 79174
rect 257514 78854 258134 78938
rect 257514 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 258134 78854
rect 257514 43174 258134 78618
rect 257514 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 258134 43174
rect 257514 42854 258134 42938
rect 257514 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 258134 42854
rect 257514 7174 258134 42618
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -2266 258134 6618
rect 257514 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 258134 -2266
rect 257514 -2586 258134 -2502
rect 257514 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 258134 -2586
rect 257514 -3814 258134 -2822
rect 261234 370894 261854 398000
rect 262078 397357 262138 399470
rect 262814 399470 262908 399530
rect 263528 399530 263588 400106
rect 263936 399530 263996 400106
rect 265296 399530 265356 400106
rect 265976 399530 266036 400106
rect 266384 399530 266444 400106
rect 267608 399530 267668 400106
rect 263528 399470 263610 399530
rect 262075 397356 262141 397357
rect 262075 397292 262076 397356
rect 262140 397292 262141 397356
rect 262075 397291 262141 397292
rect 262814 396813 262874 399470
rect 263550 396813 263610 399470
rect 263918 399470 263996 399530
rect 265206 399470 265356 399530
rect 265942 399470 266036 399530
rect 266310 399470 266444 399530
rect 267598 399470 267668 399530
rect 268288 399530 268348 400106
rect 268696 399530 268756 400106
rect 269784 399530 269844 400106
rect 271008 399530 271068 400106
rect 268288 399470 268394 399530
rect 268696 399470 268762 399530
rect 269784 399470 269866 399530
rect 262811 396812 262877 396813
rect 262811 396748 262812 396812
rect 262876 396748 262877 396812
rect 262811 396747 262877 396748
rect 263547 396812 263613 396813
rect 263547 396748 263548 396812
rect 263612 396748 263613 396812
rect 263547 396747 263613 396748
rect 263918 396677 263978 399470
rect 265206 398173 265266 399470
rect 265203 398172 265269 398173
rect 265203 398108 265204 398172
rect 265268 398108 265269 398172
rect 265203 398107 265269 398108
rect 263915 396676 263981 396677
rect 263915 396612 263916 396676
rect 263980 396612 263981 396676
rect 263915 396611 263981 396612
rect 261234 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 261854 370894
rect 261234 370574 261854 370658
rect 261234 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 261854 370574
rect 261234 334894 261854 370338
rect 261234 334658 261266 334894
rect 261502 334658 261586 334894
rect 261822 334658 261854 334894
rect 261234 334574 261854 334658
rect 261234 334338 261266 334574
rect 261502 334338 261586 334574
rect 261822 334338 261854 334574
rect 261234 298894 261854 334338
rect 261234 298658 261266 298894
rect 261502 298658 261586 298894
rect 261822 298658 261854 298894
rect 261234 298574 261854 298658
rect 261234 298338 261266 298574
rect 261502 298338 261586 298574
rect 261822 298338 261854 298574
rect 261234 262894 261854 298338
rect 261234 262658 261266 262894
rect 261502 262658 261586 262894
rect 261822 262658 261854 262894
rect 261234 262574 261854 262658
rect 261234 262338 261266 262574
rect 261502 262338 261586 262574
rect 261822 262338 261854 262574
rect 261234 226894 261854 262338
rect 261234 226658 261266 226894
rect 261502 226658 261586 226894
rect 261822 226658 261854 226894
rect 261234 226574 261854 226658
rect 261234 226338 261266 226574
rect 261502 226338 261586 226574
rect 261822 226338 261854 226574
rect 261234 190894 261854 226338
rect 261234 190658 261266 190894
rect 261502 190658 261586 190894
rect 261822 190658 261854 190894
rect 261234 190574 261854 190658
rect 261234 190338 261266 190574
rect 261502 190338 261586 190574
rect 261822 190338 261854 190574
rect 261234 154894 261854 190338
rect 261234 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 261854 154894
rect 261234 154574 261854 154658
rect 261234 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 261854 154574
rect 261234 118894 261854 154338
rect 261234 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 261854 118894
rect 261234 118574 261854 118658
rect 261234 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 261854 118574
rect 261234 82894 261854 118338
rect 261234 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 261854 82894
rect 261234 82574 261854 82658
rect 261234 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 261854 82574
rect 261234 46894 261854 82338
rect 261234 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 261854 46894
rect 261234 46574 261854 46658
rect 261234 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 261854 46574
rect 261234 10894 261854 46338
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -4186 261854 10338
rect 261234 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 261854 -4186
rect 261234 -4506 261854 -4422
rect 261234 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 261854 -4506
rect 261234 -5734 261854 -4742
rect 264954 374614 265574 398000
rect 265942 397357 266002 399470
rect 265939 397356 266005 397357
rect 265939 397292 265940 397356
rect 266004 397292 266005 397356
rect 265939 397291 266005 397292
rect 266310 396813 266370 399470
rect 266307 396812 266373 396813
rect 266307 396748 266308 396812
rect 266372 396748 266373 396812
rect 266307 396747 266373 396748
rect 267598 396677 267658 399470
rect 268334 397357 268394 399470
rect 268331 397356 268397 397357
rect 268331 397292 268332 397356
rect 268396 397292 268397 397356
rect 268331 397291 268397 397292
rect 268702 396813 268762 399470
rect 269806 396813 269866 399470
rect 270910 399470 271068 399530
rect 271144 399530 271204 400106
rect 272232 399530 272292 400106
rect 273320 399530 273380 400106
rect 273592 399530 273652 400106
rect 274408 399530 274468 400106
rect 275768 399530 275828 400106
rect 271144 399470 271338 399530
rect 272232 399470 272626 399530
rect 270910 397357 270970 399470
rect 270907 397356 270973 397357
rect 270907 397292 270908 397356
rect 270972 397292 270973 397356
rect 270907 397291 270973 397292
rect 271278 396813 271338 399470
rect 268699 396812 268765 396813
rect 268699 396748 268700 396812
rect 268764 396748 268765 396812
rect 268699 396747 268765 396748
rect 269803 396812 269869 396813
rect 269803 396748 269804 396812
rect 269868 396748 269869 396812
rect 269803 396747 269869 396748
rect 271275 396812 271341 396813
rect 271275 396748 271276 396812
rect 271340 396748 271341 396812
rect 271275 396747 271341 396748
rect 267595 396676 267661 396677
rect 267595 396612 267596 396676
rect 267660 396612 267661 396676
rect 267595 396611 267661 396612
rect 264954 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 265574 374614
rect 264954 374294 265574 374378
rect 264954 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 265574 374294
rect 264954 338614 265574 374058
rect 264954 338378 264986 338614
rect 265222 338378 265306 338614
rect 265542 338378 265574 338614
rect 264954 338294 265574 338378
rect 264954 338058 264986 338294
rect 265222 338058 265306 338294
rect 265542 338058 265574 338294
rect 264954 302614 265574 338058
rect 264954 302378 264986 302614
rect 265222 302378 265306 302614
rect 265542 302378 265574 302614
rect 264954 302294 265574 302378
rect 264954 302058 264986 302294
rect 265222 302058 265306 302294
rect 265542 302058 265574 302294
rect 264954 266614 265574 302058
rect 264954 266378 264986 266614
rect 265222 266378 265306 266614
rect 265542 266378 265574 266614
rect 264954 266294 265574 266378
rect 264954 266058 264986 266294
rect 265222 266058 265306 266294
rect 265542 266058 265574 266294
rect 264954 230614 265574 266058
rect 264954 230378 264986 230614
rect 265222 230378 265306 230614
rect 265542 230378 265574 230614
rect 264954 230294 265574 230378
rect 264954 230058 264986 230294
rect 265222 230058 265306 230294
rect 265542 230058 265574 230294
rect 264954 194614 265574 230058
rect 264954 194378 264986 194614
rect 265222 194378 265306 194614
rect 265542 194378 265574 194614
rect 264954 194294 265574 194378
rect 264954 194058 264986 194294
rect 265222 194058 265306 194294
rect 265542 194058 265574 194294
rect 264954 158614 265574 194058
rect 264954 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 265574 158614
rect 264954 158294 265574 158378
rect 264954 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 265574 158294
rect 264954 122614 265574 158058
rect 264954 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 265574 122614
rect 264954 122294 265574 122378
rect 264954 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 265574 122294
rect 264954 86614 265574 122058
rect 264954 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 265574 86614
rect 264954 86294 265574 86378
rect 264954 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 265574 86294
rect 264954 50614 265574 86058
rect 264954 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 265574 50614
rect 264954 50294 265574 50378
rect 264954 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 265574 50294
rect 264954 14614 265574 50058
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 246954 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 247574 -7066
rect 246954 -7386 247574 -7302
rect 246954 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 247574 -7386
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 14058
rect 271794 381454 272414 398000
rect 272566 397357 272626 399470
rect 273302 399470 273380 399530
rect 273486 399470 273652 399530
rect 274406 399470 274468 399530
rect 275326 399470 275828 399530
rect 276040 399530 276100 400106
rect 276992 399530 277052 400106
rect 276040 399470 276306 399530
rect 272563 397356 272629 397357
rect 272563 397292 272564 397356
rect 272628 397292 272629 397356
rect 272563 397291 272629 397292
rect 273302 396813 273362 399470
rect 273486 397221 273546 399470
rect 274406 397357 274466 399470
rect 274403 397356 274469 397357
rect 274403 397292 274404 397356
rect 274468 397292 274469 397356
rect 274403 397291 274469 397292
rect 273483 397220 273549 397221
rect 273483 397156 273484 397220
rect 273548 397156 273549 397220
rect 273483 397155 273549 397156
rect 275326 396813 275386 399470
rect 273299 396812 273365 396813
rect 273299 396748 273300 396812
rect 273364 396748 273365 396812
rect 273299 396747 273365 396748
rect 275323 396812 275389 396813
rect 275323 396748 275324 396812
rect 275388 396748 275389 396812
rect 275323 396747 275389 396748
rect 271794 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 272414 381454
rect 271794 381134 272414 381218
rect 271794 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 272414 381134
rect 271794 345454 272414 380898
rect 271794 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 272414 345454
rect 271794 345134 272414 345218
rect 271794 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 272414 345134
rect 271794 309454 272414 344898
rect 271794 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 272414 309454
rect 271794 309134 272414 309218
rect 271794 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 272414 309134
rect 271794 273454 272414 308898
rect 271794 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 272414 273454
rect 271794 273134 272414 273218
rect 271794 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 272414 273134
rect 271794 237454 272414 272898
rect 271794 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 272414 237454
rect 271794 237134 272414 237218
rect 271794 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 272414 237134
rect 271794 201454 272414 236898
rect 271794 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 272414 201454
rect 271794 201134 272414 201218
rect 271794 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 272414 201134
rect 271794 165454 272414 200898
rect 271794 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 272414 165454
rect 271794 165134 272414 165218
rect 271794 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 272414 165134
rect 271794 129454 272414 164898
rect 271794 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 272414 129454
rect 271794 129134 272414 129218
rect 271794 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 272414 129134
rect 271794 93454 272414 128898
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -1306 272414 20898
rect 271794 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 272414 -1306
rect 271794 -1626 272414 -1542
rect 271794 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 272414 -1626
rect 271794 -1894 272414 -1862
rect 275514 385174 276134 398000
rect 276246 397357 276306 399470
rect 276982 399470 277052 399530
rect 278080 399530 278140 400106
rect 278488 399530 278548 400106
rect 279168 399530 279228 400106
rect 280936 399530 280996 400106
rect 278080 399470 278146 399530
rect 276982 397357 277042 399470
rect 278086 397357 278146 399470
rect 278454 399470 278548 399530
rect 279006 399470 279228 399530
rect 280846 399470 280996 399530
rect 283520 399530 283580 400106
rect 285968 399530 286028 400106
rect 288280 399530 288340 400106
rect 291000 399530 291060 400106
rect 293448 399530 293508 400106
rect 283520 399470 283850 399530
rect 285968 399470 286058 399530
rect 276243 397356 276309 397357
rect 276243 397292 276244 397356
rect 276308 397292 276309 397356
rect 276243 397291 276309 397292
rect 276979 397356 277045 397357
rect 276979 397292 276980 397356
rect 277044 397292 277045 397356
rect 276979 397291 277045 397292
rect 278083 397356 278149 397357
rect 278083 397292 278084 397356
rect 278148 397292 278149 397356
rect 278083 397291 278149 397292
rect 278454 396813 278514 399470
rect 279006 397357 279066 399470
rect 279003 397356 279069 397357
rect 279003 397292 279004 397356
rect 279068 397292 279069 397356
rect 279003 397291 279069 397292
rect 278451 396812 278517 396813
rect 278451 396748 278452 396812
rect 278516 396748 278517 396812
rect 278451 396747 278517 396748
rect 275514 384938 275546 385174
rect 275782 384938 275866 385174
rect 276102 384938 276134 385174
rect 275514 384854 276134 384938
rect 275514 384618 275546 384854
rect 275782 384618 275866 384854
rect 276102 384618 276134 384854
rect 275514 349174 276134 384618
rect 275514 348938 275546 349174
rect 275782 348938 275866 349174
rect 276102 348938 276134 349174
rect 275514 348854 276134 348938
rect 275514 348618 275546 348854
rect 275782 348618 275866 348854
rect 276102 348618 276134 348854
rect 275514 313174 276134 348618
rect 275514 312938 275546 313174
rect 275782 312938 275866 313174
rect 276102 312938 276134 313174
rect 275514 312854 276134 312938
rect 275514 312618 275546 312854
rect 275782 312618 275866 312854
rect 276102 312618 276134 312854
rect 275514 277174 276134 312618
rect 275514 276938 275546 277174
rect 275782 276938 275866 277174
rect 276102 276938 276134 277174
rect 275514 276854 276134 276938
rect 275514 276618 275546 276854
rect 275782 276618 275866 276854
rect 276102 276618 276134 276854
rect 275514 241174 276134 276618
rect 275514 240938 275546 241174
rect 275782 240938 275866 241174
rect 276102 240938 276134 241174
rect 275514 240854 276134 240938
rect 275514 240618 275546 240854
rect 275782 240618 275866 240854
rect 276102 240618 276134 240854
rect 275514 205174 276134 240618
rect 275514 204938 275546 205174
rect 275782 204938 275866 205174
rect 276102 204938 276134 205174
rect 275514 204854 276134 204938
rect 275514 204618 275546 204854
rect 275782 204618 275866 204854
rect 276102 204618 276134 204854
rect 275514 169174 276134 204618
rect 275514 168938 275546 169174
rect 275782 168938 275866 169174
rect 276102 168938 276134 169174
rect 275514 168854 276134 168938
rect 275514 168618 275546 168854
rect 275782 168618 275866 168854
rect 276102 168618 276134 168854
rect 275514 133174 276134 168618
rect 275514 132938 275546 133174
rect 275782 132938 275866 133174
rect 276102 132938 276134 133174
rect 275514 132854 276134 132938
rect 275514 132618 275546 132854
rect 275782 132618 275866 132854
rect 276102 132618 276134 132854
rect 275514 97174 276134 132618
rect 275514 96938 275546 97174
rect 275782 96938 275866 97174
rect 276102 96938 276134 97174
rect 275514 96854 276134 96938
rect 275514 96618 275546 96854
rect 275782 96618 275866 96854
rect 276102 96618 276134 96854
rect 275514 61174 276134 96618
rect 275514 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 276134 61174
rect 275514 60854 276134 60938
rect 275514 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 276134 60854
rect 275514 25174 276134 60618
rect 275514 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 276134 25174
rect 275514 24854 276134 24938
rect 275514 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 276134 24854
rect 275514 -3226 276134 24618
rect 275514 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 276134 -3226
rect 275514 -3546 276134 -3462
rect 275514 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 276134 -3546
rect 275514 -3814 276134 -3782
rect 279234 388894 279854 398000
rect 280846 396813 280906 399470
rect 280843 396812 280909 396813
rect 280843 396748 280844 396812
rect 280908 396748 280909 396812
rect 280843 396747 280909 396748
rect 279234 388658 279266 388894
rect 279502 388658 279586 388894
rect 279822 388658 279854 388894
rect 279234 388574 279854 388658
rect 279234 388338 279266 388574
rect 279502 388338 279586 388574
rect 279822 388338 279854 388574
rect 279234 352894 279854 388338
rect 279234 352658 279266 352894
rect 279502 352658 279586 352894
rect 279822 352658 279854 352894
rect 279234 352574 279854 352658
rect 279234 352338 279266 352574
rect 279502 352338 279586 352574
rect 279822 352338 279854 352574
rect 279234 316894 279854 352338
rect 279234 316658 279266 316894
rect 279502 316658 279586 316894
rect 279822 316658 279854 316894
rect 279234 316574 279854 316658
rect 279234 316338 279266 316574
rect 279502 316338 279586 316574
rect 279822 316338 279854 316574
rect 279234 280894 279854 316338
rect 279234 280658 279266 280894
rect 279502 280658 279586 280894
rect 279822 280658 279854 280894
rect 279234 280574 279854 280658
rect 279234 280338 279266 280574
rect 279502 280338 279586 280574
rect 279822 280338 279854 280574
rect 279234 244894 279854 280338
rect 279234 244658 279266 244894
rect 279502 244658 279586 244894
rect 279822 244658 279854 244894
rect 279234 244574 279854 244658
rect 279234 244338 279266 244574
rect 279502 244338 279586 244574
rect 279822 244338 279854 244574
rect 279234 208894 279854 244338
rect 279234 208658 279266 208894
rect 279502 208658 279586 208894
rect 279822 208658 279854 208894
rect 279234 208574 279854 208658
rect 279234 208338 279266 208574
rect 279502 208338 279586 208574
rect 279822 208338 279854 208574
rect 279234 172894 279854 208338
rect 279234 172658 279266 172894
rect 279502 172658 279586 172894
rect 279822 172658 279854 172894
rect 279234 172574 279854 172658
rect 279234 172338 279266 172574
rect 279502 172338 279586 172574
rect 279822 172338 279854 172574
rect 279234 136894 279854 172338
rect 279234 136658 279266 136894
rect 279502 136658 279586 136894
rect 279822 136658 279854 136894
rect 279234 136574 279854 136658
rect 279234 136338 279266 136574
rect 279502 136338 279586 136574
rect 279822 136338 279854 136574
rect 279234 100894 279854 136338
rect 279234 100658 279266 100894
rect 279502 100658 279586 100894
rect 279822 100658 279854 100894
rect 279234 100574 279854 100658
rect 279234 100338 279266 100574
rect 279502 100338 279586 100574
rect 279822 100338 279854 100574
rect 279234 64894 279854 100338
rect 279234 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 279854 64894
rect 279234 64574 279854 64658
rect 279234 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 279854 64574
rect 279234 28894 279854 64338
rect 279234 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 279854 28894
rect 279234 28574 279854 28658
rect 279234 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 279854 28574
rect 279234 -5146 279854 28338
rect 279234 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 279854 -5146
rect 279234 -5466 279854 -5382
rect 279234 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 279854 -5466
rect 279234 -5734 279854 -5702
rect 282954 392614 283574 398000
rect 283790 397357 283850 399470
rect 283787 397356 283853 397357
rect 283787 397292 283788 397356
rect 283852 397292 283853 397356
rect 283787 397291 283853 397292
rect 285998 396813 286058 399470
rect 288206 399470 288340 399530
rect 290966 399470 291060 399530
rect 293358 399470 293508 399530
rect 295896 399530 295956 400106
rect 298480 399530 298540 400106
rect 300928 399530 300988 400106
rect 303512 399530 303572 400106
rect 305960 399530 306020 400106
rect 295896 399470 295994 399530
rect 298480 399470 298570 399530
rect 288206 396813 288266 399470
rect 285995 396812 286061 396813
rect 285995 396748 285996 396812
rect 286060 396748 286061 396812
rect 285995 396747 286061 396748
rect 288203 396812 288269 396813
rect 288203 396748 288204 396812
rect 288268 396748 288269 396812
rect 288203 396747 288269 396748
rect 282954 392378 282986 392614
rect 283222 392378 283306 392614
rect 283542 392378 283574 392614
rect 282954 392294 283574 392378
rect 282954 392058 282986 392294
rect 283222 392058 283306 392294
rect 283542 392058 283574 392294
rect 282954 356614 283574 392058
rect 282954 356378 282986 356614
rect 283222 356378 283306 356614
rect 283542 356378 283574 356614
rect 282954 356294 283574 356378
rect 282954 356058 282986 356294
rect 283222 356058 283306 356294
rect 283542 356058 283574 356294
rect 282954 320614 283574 356058
rect 282954 320378 282986 320614
rect 283222 320378 283306 320614
rect 283542 320378 283574 320614
rect 282954 320294 283574 320378
rect 282954 320058 282986 320294
rect 283222 320058 283306 320294
rect 283542 320058 283574 320294
rect 282954 284614 283574 320058
rect 282954 284378 282986 284614
rect 283222 284378 283306 284614
rect 283542 284378 283574 284614
rect 282954 284294 283574 284378
rect 282954 284058 282986 284294
rect 283222 284058 283306 284294
rect 283542 284058 283574 284294
rect 282954 248614 283574 284058
rect 282954 248378 282986 248614
rect 283222 248378 283306 248614
rect 283542 248378 283574 248614
rect 282954 248294 283574 248378
rect 282954 248058 282986 248294
rect 283222 248058 283306 248294
rect 283542 248058 283574 248294
rect 282954 212614 283574 248058
rect 282954 212378 282986 212614
rect 283222 212378 283306 212614
rect 283542 212378 283574 212614
rect 282954 212294 283574 212378
rect 282954 212058 282986 212294
rect 283222 212058 283306 212294
rect 283542 212058 283574 212294
rect 282954 176614 283574 212058
rect 282954 176378 282986 176614
rect 283222 176378 283306 176614
rect 283542 176378 283574 176614
rect 282954 176294 283574 176378
rect 282954 176058 282986 176294
rect 283222 176058 283306 176294
rect 283542 176058 283574 176294
rect 282954 140614 283574 176058
rect 282954 140378 282986 140614
rect 283222 140378 283306 140614
rect 283542 140378 283574 140614
rect 282954 140294 283574 140378
rect 282954 140058 282986 140294
rect 283222 140058 283306 140294
rect 283542 140058 283574 140294
rect 282954 104614 283574 140058
rect 282954 104378 282986 104614
rect 283222 104378 283306 104614
rect 283542 104378 283574 104614
rect 282954 104294 283574 104378
rect 282954 104058 282986 104294
rect 283222 104058 283306 104294
rect 283542 104058 283574 104294
rect 282954 68614 283574 104058
rect 282954 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 283574 68614
rect 282954 68294 283574 68378
rect 282954 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 283574 68294
rect 282954 32614 283574 68058
rect 282954 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 283574 32614
rect 282954 32294 283574 32378
rect 282954 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 283574 32294
rect 264954 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 265574 -6106
rect 264954 -6426 265574 -6342
rect 264954 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 265574 -6426
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 32058
rect 289794 363454 290414 398000
rect 290966 397357 291026 399470
rect 290963 397356 291029 397357
rect 290963 397292 290964 397356
rect 291028 397292 291029 397356
rect 290963 397291 291029 397292
rect 293358 396813 293418 399470
rect 293355 396812 293421 396813
rect 293355 396748 293356 396812
rect 293420 396748 293421 396812
rect 293355 396747 293421 396748
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 289794 327454 290414 362898
rect 289794 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 290414 327454
rect 289794 327134 290414 327218
rect 289794 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 290414 327134
rect 289794 291454 290414 326898
rect 289794 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 290414 291454
rect 289794 291134 290414 291218
rect 289794 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 290414 291134
rect 289794 255454 290414 290898
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 289794 219454 290414 254898
rect 289794 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 290414 219454
rect 289794 219134 290414 219218
rect 289794 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 290414 219134
rect 289794 183454 290414 218898
rect 289794 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 290414 183454
rect 289794 183134 290414 183218
rect 289794 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 290414 183134
rect 289794 147454 290414 182898
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 111454 290414 146898
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 289794 75454 290414 110898
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 293514 367174 294134 398000
rect 295934 396813 295994 399470
rect 295931 396812 295997 396813
rect 295931 396748 295932 396812
rect 295996 396748 295997 396812
rect 295931 396747 295997 396748
rect 293514 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 294134 367174
rect 293514 366854 294134 366938
rect 293514 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 294134 366854
rect 293514 331174 294134 366618
rect 293514 330938 293546 331174
rect 293782 330938 293866 331174
rect 294102 330938 294134 331174
rect 293514 330854 294134 330938
rect 293514 330618 293546 330854
rect 293782 330618 293866 330854
rect 294102 330618 294134 330854
rect 293514 295174 294134 330618
rect 293514 294938 293546 295174
rect 293782 294938 293866 295174
rect 294102 294938 294134 295174
rect 293514 294854 294134 294938
rect 293514 294618 293546 294854
rect 293782 294618 293866 294854
rect 294102 294618 294134 294854
rect 293514 259174 294134 294618
rect 293514 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 294134 259174
rect 293514 258854 294134 258938
rect 293514 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 294134 258854
rect 293514 223174 294134 258618
rect 293514 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 294134 223174
rect 293514 222854 294134 222938
rect 293514 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 294134 222854
rect 293514 187174 294134 222618
rect 293514 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 294134 187174
rect 293514 186854 294134 186938
rect 293514 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 294134 186854
rect 293514 151174 294134 186618
rect 293514 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 294134 151174
rect 293514 150854 294134 150938
rect 293514 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 294134 150854
rect 293514 115174 294134 150618
rect 293514 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 294134 115174
rect 293514 114854 294134 114938
rect 293514 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 294134 114854
rect 293514 79174 294134 114618
rect 293514 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 294134 79174
rect 293514 78854 294134 78938
rect 293514 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 294134 78854
rect 293514 43174 294134 78618
rect 293514 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 294134 43174
rect 293514 42854 294134 42938
rect 293514 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 294134 42854
rect 293514 7174 294134 42618
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -2266 294134 6618
rect 293514 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 294134 -2266
rect 293514 -2586 294134 -2502
rect 293514 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 294134 -2586
rect 293514 -3814 294134 -2822
rect 297234 370894 297854 398000
rect 298510 397357 298570 399470
rect 300902 399470 300988 399530
rect 303478 399470 303572 399530
rect 305870 399470 306020 399530
rect 308544 399530 308604 400106
rect 310992 399530 311052 400106
rect 313440 399530 313500 400106
rect 315888 399530 315948 400106
rect 318472 399530 318532 400106
rect 308544 399470 308690 399530
rect 310992 399470 311082 399530
rect 300902 398173 300962 399470
rect 300899 398172 300965 398173
rect 300899 398108 300900 398172
rect 300964 398108 300965 398172
rect 300899 398107 300965 398108
rect 298507 397356 298573 397357
rect 298507 397292 298508 397356
rect 298572 397292 298573 397356
rect 298507 397291 298573 397292
rect 297234 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 297854 370894
rect 297234 370574 297854 370658
rect 297234 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 297854 370574
rect 297234 334894 297854 370338
rect 297234 334658 297266 334894
rect 297502 334658 297586 334894
rect 297822 334658 297854 334894
rect 297234 334574 297854 334658
rect 297234 334338 297266 334574
rect 297502 334338 297586 334574
rect 297822 334338 297854 334574
rect 297234 298894 297854 334338
rect 297234 298658 297266 298894
rect 297502 298658 297586 298894
rect 297822 298658 297854 298894
rect 297234 298574 297854 298658
rect 297234 298338 297266 298574
rect 297502 298338 297586 298574
rect 297822 298338 297854 298574
rect 297234 262894 297854 298338
rect 297234 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 297854 262894
rect 297234 262574 297854 262658
rect 297234 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 297854 262574
rect 297234 226894 297854 262338
rect 297234 226658 297266 226894
rect 297502 226658 297586 226894
rect 297822 226658 297854 226894
rect 297234 226574 297854 226658
rect 297234 226338 297266 226574
rect 297502 226338 297586 226574
rect 297822 226338 297854 226574
rect 297234 190894 297854 226338
rect 297234 190658 297266 190894
rect 297502 190658 297586 190894
rect 297822 190658 297854 190894
rect 297234 190574 297854 190658
rect 297234 190338 297266 190574
rect 297502 190338 297586 190574
rect 297822 190338 297854 190574
rect 297234 154894 297854 190338
rect 297234 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 297854 154894
rect 297234 154574 297854 154658
rect 297234 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 297854 154574
rect 297234 118894 297854 154338
rect 297234 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 297854 118894
rect 297234 118574 297854 118658
rect 297234 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 297854 118574
rect 297234 82894 297854 118338
rect 297234 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 297854 82894
rect 297234 82574 297854 82658
rect 297234 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 297854 82574
rect 297234 46894 297854 82338
rect 297234 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 297854 46894
rect 297234 46574 297854 46658
rect 297234 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 297854 46574
rect 297234 10894 297854 46338
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -4186 297854 10338
rect 297234 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 297854 -4186
rect 297234 -4506 297854 -4422
rect 297234 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 297854 -4506
rect 297234 -5734 297854 -4742
rect 300954 374614 301574 398000
rect 303478 396813 303538 399470
rect 305870 396813 305930 399470
rect 303475 396812 303541 396813
rect 303475 396748 303476 396812
rect 303540 396748 303541 396812
rect 303475 396747 303541 396748
rect 305867 396812 305933 396813
rect 305867 396748 305868 396812
rect 305932 396748 305933 396812
rect 305867 396747 305933 396748
rect 300954 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 301574 374614
rect 300954 374294 301574 374378
rect 300954 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 301574 374294
rect 300954 338614 301574 374058
rect 300954 338378 300986 338614
rect 301222 338378 301306 338614
rect 301542 338378 301574 338614
rect 300954 338294 301574 338378
rect 300954 338058 300986 338294
rect 301222 338058 301306 338294
rect 301542 338058 301574 338294
rect 300954 302614 301574 338058
rect 300954 302378 300986 302614
rect 301222 302378 301306 302614
rect 301542 302378 301574 302614
rect 300954 302294 301574 302378
rect 300954 302058 300986 302294
rect 301222 302058 301306 302294
rect 301542 302058 301574 302294
rect 300954 266614 301574 302058
rect 300954 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 301574 266614
rect 300954 266294 301574 266378
rect 300954 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 301574 266294
rect 300954 230614 301574 266058
rect 300954 230378 300986 230614
rect 301222 230378 301306 230614
rect 301542 230378 301574 230614
rect 300954 230294 301574 230378
rect 300954 230058 300986 230294
rect 301222 230058 301306 230294
rect 301542 230058 301574 230294
rect 300954 194614 301574 230058
rect 300954 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 301574 194614
rect 300954 194294 301574 194378
rect 300954 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 301574 194294
rect 300954 158614 301574 194058
rect 300954 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 301574 158614
rect 300954 158294 301574 158378
rect 300954 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 301574 158294
rect 300954 122614 301574 158058
rect 300954 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 301574 122614
rect 300954 122294 301574 122378
rect 300954 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 301574 122294
rect 300954 86614 301574 122058
rect 300954 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 301574 86614
rect 300954 86294 301574 86378
rect 300954 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 301574 86294
rect 300954 50614 301574 86058
rect 300954 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 301574 50614
rect 300954 50294 301574 50378
rect 300954 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 301574 50294
rect 300954 14614 301574 50058
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 282954 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 283574 -7066
rect 282954 -7386 283574 -7302
rect 282954 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 283574 -7386
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 14058
rect 307794 381454 308414 398000
rect 308630 396813 308690 399470
rect 311022 396813 311082 399470
rect 313414 399470 313500 399530
rect 315806 399470 315948 399530
rect 318382 399470 318532 399530
rect 320920 399530 320980 400106
rect 323368 399530 323428 400106
rect 325952 399530 326012 400106
rect 343224 399530 343284 400106
rect 320920 399470 321018 399530
rect 308627 396812 308693 396813
rect 308627 396748 308628 396812
rect 308692 396748 308693 396812
rect 308627 396747 308693 396748
rect 311019 396812 311085 396813
rect 311019 396748 311020 396812
rect 311084 396748 311085 396812
rect 311019 396747 311085 396748
rect 307794 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 308414 381454
rect 307794 381134 308414 381218
rect 307794 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 308414 381134
rect 307794 345454 308414 380898
rect 307794 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 308414 345454
rect 307794 345134 308414 345218
rect 307794 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 308414 345134
rect 307794 309454 308414 344898
rect 307794 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 308414 309454
rect 307794 309134 308414 309218
rect 307794 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 308414 309134
rect 307794 273454 308414 308898
rect 307794 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 308414 273454
rect 307794 273134 308414 273218
rect 307794 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 308414 273134
rect 307794 237454 308414 272898
rect 307794 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 308414 237454
rect 307794 237134 308414 237218
rect 307794 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 308414 237134
rect 307794 201454 308414 236898
rect 307794 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 308414 201454
rect 307794 201134 308414 201218
rect 307794 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 308414 201134
rect 307794 165454 308414 200898
rect 307794 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 308414 165454
rect 307794 165134 308414 165218
rect 307794 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 308414 165134
rect 307794 129454 308414 164898
rect 307794 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 308414 129454
rect 307794 129134 308414 129218
rect 307794 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 308414 129134
rect 307794 93454 308414 128898
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -1306 308414 20898
rect 307794 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 308414 -1306
rect 307794 -1626 308414 -1542
rect 307794 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 308414 -1626
rect 307794 -1894 308414 -1862
rect 311514 385174 312134 398000
rect 313414 396813 313474 399470
rect 315806 398173 315866 399470
rect 315803 398172 315869 398173
rect 315803 398108 315804 398172
rect 315868 398108 315869 398172
rect 315803 398107 315869 398108
rect 313411 396812 313477 396813
rect 313411 396748 313412 396812
rect 313476 396748 313477 396812
rect 313411 396747 313477 396748
rect 311514 384938 311546 385174
rect 311782 384938 311866 385174
rect 312102 384938 312134 385174
rect 311514 384854 312134 384938
rect 311514 384618 311546 384854
rect 311782 384618 311866 384854
rect 312102 384618 312134 384854
rect 311514 349174 312134 384618
rect 311514 348938 311546 349174
rect 311782 348938 311866 349174
rect 312102 348938 312134 349174
rect 311514 348854 312134 348938
rect 311514 348618 311546 348854
rect 311782 348618 311866 348854
rect 312102 348618 312134 348854
rect 311514 313174 312134 348618
rect 311514 312938 311546 313174
rect 311782 312938 311866 313174
rect 312102 312938 312134 313174
rect 311514 312854 312134 312938
rect 311514 312618 311546 312854
rect 311782 312618 311866 312854
rect 312102 312618 312134 312854
rect 311514 277174 312134 312618
rect 311514 276938 311546 277174
rect 311782 276938 311866 277174
rect 312102 276938 312134 277174
rect 311514 276854 312134 276938
rect 311514 276618 311546 276854
rect 311782 276618 311866 276854
rect 312102 276618 312134 276854
rect 311514 241174 312134 276618
rect 311514 240938 311546 241174
rect 311782 240938 311866 241174
rect 312102 240938 312134 241174
rect 311514 240854 312134 240938
rect 311514 240618 311546 240854
rect 311782 240618 311866 240854
rect 312102 240618 312134 240854
rect 311514 205174 312134 240618
rect 311514 204938 311546 205174
rect 311782 204938 311866 205174
rect 312102 204938 312134 205174
rect 311514 204854 312134 204938
rect 311514 204618 311546 204854
rect 311782 204618 311866 204854
rect 312102 204618 312134 204854
rect 311514 169174 312134 204618
rect 311514 168938 311546 169174
rect 311782 168938 311866 169174
rect 312102 168938 312134 169174
rect 311514 168854 312134 168938
rect 311514 168618 311546 168854
rect 311782 168618 311866 168854
rect 312102 168618 312134 168854
rect 311514 133174 312134 168618
rect 311514 132938 311546 133174
rect 311782 132938 311866 133174
rect 312102 132938 312134 133174
rect 311514 132854 312134 132938
rect 311514 132618 311546 132854
rect 311782 132618 311866 132854
rect 312102 132618 312134 132854
rect 311514 97174 312134 132618
rect 311514 96938 311546 97174
rect 311782 96938 311866 97174
rect 312102 96938 312134 97174
rect 311514 96854 312134 96938
rect 311514 96618 311546 96854
rect 311782 96618 311866 96854
rect 312102 96618 312134 96854
rect 311514 61174 312134 96618
rect 311514 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 312134 61174
rect 311514 60854 312134 60938
rect 311514 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 312134 60854
rect 311514 25174 312134 60618
rect 311514 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 312134 25174
rect 311514 24854 312134 24938
rect 311514 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 312134 24854
rect 311514 -3226 312134 24618
rect 311514 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 312134 -3226
rect 311514 -3546 312134 -3462
rect 311514 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 312134 -3546
rect 311514 -3814 312134 -3782
rect 315234 388894 315854 398000
rect 318382 396813 318442 399470
rect 318379 396812 318445 396813
rect 318379 396748 318380 396812
rect 318444 396748 318445 396812
rect 318379 396747 318445 396748
rect 315234 388658 315266 388894
rect 315502 388658 315586 388894
rect 315822 388658 315854 388894
rect 315234 388574 315854 388658
rect 315234 388338 315266 388574
rect 315502 388338 315586 388574
rect 315822 388338 315854 388574
rect 315234 352894 315854 388338
rect 315234 352658 315266 352894
rect 315502 352658 315586 352894
rect 315822 352658 315854 352894
rect 315234 352574 315854 352658
rect 315234 352338 315266 352574
rect 315502 352338 315586 352574
rect 315822 352338 315854 352574
rect 315234 316894 315854 352338
rect 315234 316658 315266 316894
rect 315502 316658 315586 316894
rect 315822 316658 315854 316894
rect 315234 316574 315854 316658
rect 315234 316338 315266 316574
rect 315502 316338 315586 316574
rect 315822 316338 315854 316574
rect 315234 280894 315854 316338
rect 315234 280658 315266 280894
rect 315502 280658 315586 280894
rect 315822 280658 315854 280894
rect 315234 280574 315854 280658
rect 315234 280338 315266 280574
rect 315502 280338 315586 280574
rect 315822 280338 315854 280574
rect 315234 244894 315854 280338
rect 315234 244658 315266 244894
rect 315502 244658 315586 244894
rect 315822 244658 315854 244894
rect 315234 244574 315854 244658
rect 315234 244338 315266 244574
rect 315502 244338 315586 244574
rect 315822 244338 315854 244574
rect 315234 208894 315854 244338
rect 315234 208658 315266 208894
rect 315502 208658 315586 208894
rect 315822 208658 315854 208894
rect 315234 208574 315854 208658
rect 315234 208338 315266 208574
rect 315502 208338 315586 208574
rect 315822 208338 315854 208574
rect 315234 172894 315854 208338
rect 315234 172658 315266 172894
rect 315502 172658 315586 172894
rect 315822 172658 315854 172894
rect 315234 172574 315854 172658
rect 315234 172338 315266 172574
rect 315502 172338 315586 172574
rect 315822 172338 315854 172574
rect 315234 136894 315854 172338
rect 315234 136658 315266 136894
rect 315502 136658 315586 136894
rect 315822 136658 315854 136894
rect 315234 136574 315854 136658
rect 315234 136338 315266 136574
rect 315502 136338 315586 136574
rect 315822 136338 315854 136574
rect 315234 100894 315854 136338
rect 315234 100658 315266 100894
rect 315502 100658 315586 100894
rect 315822 100658 315854 100894
rect 315234 100574 315854 100658
rect 315234 100338 315266 100574
rect 315502 100338 315586 100574
rect 315822 100338 315854 100574
rect 315234 64894 315854 100338
rect 315234 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 315854 64894
rect 315234 64574 315854 64658
rect 315234 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 315854 64574
rect 315234 28894 315854 64338
rect 315234 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 315854 28894
rect 315234 28574 315854 28658
rect 315234 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 315854 28574
rect 315234 -5146 315854 28338
rect 315234 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 315854 -5146
rect 315234 -5466 315854 -5382
rect 315234 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 315854 -5466
rect 315234 -5734 315854 -5702
rect 318954 392614 319574 398000
rect 320958 396813 321018 399470
rect 323350 399470 323428 399530
rect 325926 399470 326012 399530
rect 343222 399470 343284 399530
rect 343360 399530 343420 400106
rect 343360 399470 343466 399530
rect 323350 396813 323410 399470
rect 325926 398173 325986 399470
rect 325923 398172 325989 398173
rect 325923 398108 325924 398172
rect 325988 398108 325989 398172
rect 325923 398107 325989 398108
rect 320955 396812 321021 396813
rect 320955 396748 320956 396812
rect 321020 396748 321021 396812
rect 320955 396747 321021 396748
rect 323347 396812 323413 396813
rect 323347 396748 323348 396812
rect 323412 396748 323413 396812
rect 323347 396747 323413 396748
rect 318954 392378 318986 392614
rect 319222 392378 319306 392614
rect 319542 392378 319574 392614
rect 318954 392294 319574 392378
rect 318954 392058 318986 392294
rect 319222 392058 319306 392294
rect 319542 392058 319574 392294
rect 318954 356614 319574 392058
rect 318954 356378 318986 356614
rect 319222 356378 319306 356614
rect 319542 356378 319574 356614
rect 318954 356294 319574 356378
rect 318954 356058 318986 356294
rect 319222 356058 319306 356294
rect 319542 356058 319574 356294
rect 318954 320614 319574 356058
rect 318954 320378 318986 320614
rect 319222 320378 319306 320614
rect 319542 320378 319574 320614
rect 318954 320294 319574 320378
rect 318954 320058 318986 320294
rect 319222 320058 319306 320294
rect 319542 320058 319574 320294
rect 318954 284614 319574 320058
rect 318954 284378 318986 284614
rect 319222 284378 319306 284614
rect 319542 284378 319574 284614
rect 318954 284294 319574 284378
rect 318954 284058 318986 284294
rect 319222 284058 319306 284294
rect 319542 284058 319574 284294
rect 318954 248614 319574 284058
rect 318954 248378 318986 248614
rect 319222 248378 319306 248614
rect 319542 248378 319574 248614
rect 318954 248294 319574 248378
rect 318954 248058 318986 248294
rect 319222 248058 319306 248294
rect 319542 248058 319574 248294
rect 318954 212614 319574 248058
rect 318954 212378 318986 212614
rect 319222 212378 319306 212614
rect 319542 212378 319574 212614
rect 318954 212294 319574 212378
rect 318954 212058 318986 212294
rect 319222 212058 319306 212294
rect 319542 212058 319574 212294
rect 318954 176614 319574 212058
rect 318954 176378 318986 176614
rect 319222 176378 319306 176614
rect 319542 176378 319574 176614
rect 318954 176294 319574 176378
rect 318954 176058 318986 176294
rect 319222 176058 319306 176294
rect 319542 176058 319574 176294
rect 318954 140614 319574 176058
rect 318954 140378 318986 140614
rect 319222 140378 319306 140614
rect 319542 140378 319574 140614
rect 318954 140294 319574 140378
rect 318954 140058 318986 140294
rect 319222 140058 319306 140294
rect 319542 140058 319574 140294
rect 318954 104614 319574 140058
rect 318954 104378 318986 104614
rect 319222 104378 319306 104614
rect 319542 104378 319574 104614
rect 318954 104294 319574 104378
rect 318954 104058 318986 104294
rect 319222 104058 319306 104294
rect 319542 104058 319574 104294
rect 318954 68614 319574 104058
rect 318954 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 319574 68614
rect 318954 68294 319574 68378
rect 318954 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 319574 68294
rect 318954 32614 319574 68058
rect 318954 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 319574 32614
rect 318954 32294 319574 32378
rect 318954 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 319574 32294
rect 300954 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 301574 -6106
rect 300954 -6426 301574 -6342
rect 300954 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 301574 -6426
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 32058
rect 325794 363454 326414 398000
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325794 327454 326414 362898
rect 325794 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 326414 327454
rect 325794 327134 326414 327218
rect 325794 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 326414 327134
rect 325794 291454 326414 326898
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 219454 326414 254898
rect 325794 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 326414 219454
rect 325794 219134 326414 219218
rect 325794 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 326414 219134
rect 325794 183454 326414 218898
rect 325794 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 326414 183454
rect 325794 183134 326414 183218
rect 325794 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 326414 183134
rect 325794 147454 326414 182898
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 329514 367174 330134 398000
rect 329514 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 330134 367174
rect 329514 366854 330134 366938
rect 329514 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 330134 366854
rect 329514 331174 330134 366618
rect 329514 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 330134 331174
rect 329514 330854 330134 330938
rect 329514 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 330134 330854
rect 329514 295174 330134 330618
rect 329514 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 330134 295174
rect 329514 294854 330134 294938
rect 329514 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 330134 294854
rect 329514 259174 330134 294618
rect 329514 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 330134 259174
rect 329514 258854 330134 258938
rect 329514 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 330134 258854
rect 329514 223174 330134 258618
rect 329514 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 330134 223174
rect 329514 222854 330134 222938
rect 329514 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 330134 222854
rect 329514 187174 330134 222618
rect 329514 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 330134 187174
rect 329514 186854 330134 186938
rect 329514 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 330134 186854
rect 329514 151174 330134 186618
rect 329514 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 330134 151174
rect 329514 150854 330134 150938
rect 329514 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 330134 150854
rect 329514 115174 330134 150618
rect 329514 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 330134 115174
rect 329514 114854 330134 114938
rect 329514 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 330134 114854
rect 329514 79174 330134 114618
rect 329514 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 330134 79174
rect 329514 78854 330134 78938
rect 329514 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 330134 78854
rect 329514 43174 330134 78618
rect 329514 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 330134 43174
rect 329514 42854 330134 42938
rect 329514 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 330134 42854
rect 329514 7174 330134 42618
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -2266 330134 6618
rect 329514 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 330134 -2266
rect 329514 -2586 330134 -2502
rect 329514 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 330134 -2586
rect 329514 -3814 330134 -2822
rect 333234 370894 333854 398000
rect 333234 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 333854 370894
rect 333234 370574 333854 370658
rect 333234 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 333854 370574
rect 333234 334894 333854 370338
rect 333234 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 333854 334894
rect 333234 334574 333854 334658
rect 333234 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 333854 334574
rect 333234 298894 333854 334338
rect 333234 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 333854 298894
rect 333234 298574 333854 298658
rect 333234 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 333854 298574
rect 333234 262894 333854 298338
rect 333234 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 333854 262894
rect 333234 262574 333854 262658
rect 333234 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 333854 262574
rect 333234 226894 333854 262338
rect 333234 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 333854 226894
rect 333234 226574 333854 226658
rect 333234 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 333854 226574
rect 333234 190894 333854 226338
rect 333234 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 333854 190894
rect 333234 190574 333854 190658
rect 333234 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 333854 190574
rect 333234 154894 333854 190338
rect 333234 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 333854 154894
rect 333234 154574 333854 154658
rect 333234 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 333854 154574
rect 333234 118894 333854 154338
rect 333234 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 333854 118894
rect 333234 118574 333854 118658
rect 333234 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 333854 118574
rect 333234 82894 333854 118338
rect 333234 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 333854 82894
rect 333234 82574 333854 82658
rect 333234 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 333854 82574
rect 333234 46894 333854 82338
rect 333234 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 333854 46894
rect 333234 46574 333854 46658
rect 333234 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 333854 46574
rect 333234 10894 333854 46338
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -4186 333854 10338
rect 333234 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 333854 -4186
rect 333234 -4506 333854 -4422
rect 333234 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 333854 -4506
rect 333234 -5734 333854 -4742
rect 336954 374614 337574 398000
rect 343222 396813 343282 399470
rect 343406 397357 343466 399470
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 343403 397356 343469 397357
rect 343403 397292 343404 397356
rect 343468 397292 343469 397356
rect 343403 397291 343469 397292
rect 343219 396812 343285 396813
rect 343219 396748 343220 396812
rect 343284 396748 343285 396812
rect 343219 396747 343285 396748
rect 336954 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 337574 374614
rect 336954 374294 337574 374378
rect 336954 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 337574 374294
rect 336954 338614 337574 374058
rect 336954 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 337574 338614
rect 336954 338294 337574 338378
rect 336954 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 337574 338294
rect 336954 302614 337574 338058
rect 336954 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 337574 302614
rect 336954 302294 337574 302378
rect 336954 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 337574 302294
rect 336954 266614 337574 302058
rect 336954 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 337574 266614
rect 336954 266294 337574 266378
rect 336954 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 337574 266294
rect 336954 230614 337574 266058
rect 336954 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 337574 230614
rect 336954 230294 337574 230378
rect 336954 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 337574 230294
rect 336954 194614 337574 230058
rect 336954 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 337574 194614
rect 336954 194294 337574 194378
rect 336954 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 337574 194294
rect 336954 158614 337574 194058
rect 336954 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 337574 158614
rect 336954 158294 337574 158378
rect 336954 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 337574 158294
rect 336954 122614 337574 158058
rect 336954 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 337574 122614
rect 336954 122294 337574 122378
rect 336954 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 337574 122294
rect 336954 86614 337574 122058
rect 336954 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 337574 86614
rect 336954 86294 337574 86378
rect 336954 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 337574 86294
rect 336954 50614 337574 86058
rect 336954 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 337574 50614
rect 336954 50294 337574 50378
rect 336954 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 337574 50294
rect 336954 14614 337574 50058
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 318954 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 319574 -7066
rect 318954 -7386 319574 -7302
rect 318954 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 319574 -7386
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 14058
rect 343794 381454 344414 398000
rect 343794 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 344414 381454
rect 343794 381134 344414 381218
rect 343794 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 344414 381134
rect 343794 345454 344414 380898
rect 343794 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 344414 345454
rect 343794 345134 344414 345218
rect 343794 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 344414 345134
rect 343794 309454 344414 344898
rect 343794 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 344414 309454
rect 343794 309134 344414 309218
rect 343794 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 344414 309134
rect 343794 273454 344414 308898
rect 343794 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 344414 273454
rect 343794 273134 344414 273218
rect 343794 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 344414 273134
rect 343794 237454 344414 272898
rect 343794 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 344414 237454
rect 343794 237134 344414 237218
rect 343794 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 344414 237134
rect 343794 201454 344414 236898
rect 343794 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 344414 201454
rect 343794 201134 344414 201218
rect 343794 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 344414 201134
rect 343794 165454 344414 200898
rect 343794 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 344414 165454
rect 343794 165134 344414 165218
rect 343794 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 344414 165134
rect 343794 129454 344414 164898
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 343794 93454 344414 128898
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -1306 344414 20898
rect 343794 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 344414 -1306
rect 343794 -1626 344414 -1542
rect 343794 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 344414 -1626
rect 343794 -1894 344414 -1862
rect 347514 385174 348134 398000
rect 347514 384938 347546 385174
rect 347782 384938 347866 385174
rect 348102 384938 348134 385174
rect 347514 384854 348134 384938
rect 347514 384618 347546 384854
rect 347782 384618 347866 384854
rect 348102 384618 348134 384854
rect 347514 349174 348134 384618
rect 347514 348938 347546 349174
rect 347782 348938 347866 349174
rect 348102 348938 348134 349174
rect 347514 348854 348134 348938
rect 347514 348618 347546 348854
rect 347782 348618 347866 348854
rect 348102 348618 348134 348854
rect 347514 313174 348134 348618
rect 347514 312938 347546 313174
rect 347782 312938 347866 313174
rect 348102 312938 348134 313174
rect 347514 312854 348134 312938
rect 347514 312618 347546 312854
rect 347782 312618 347866 312854
rect 348102 312618 348134 312854
rect 347514 277174 348134 312618
rect 347514 276938 347546 277174
rect 347782 276938 347866 277174
rect 348102 276938 348134 277174
rect 347514 276854 348134 276938
rect 347514 276618 347546 276854
rect 347782 276618 347866 276854
rect 348102 276618 348134 276854
rect 347514 241174 348134 276618
rect 347514 240938 347546 241174
rect 347782 240938 347866 241174
rect 348102 240938 348134 241174
rect 347514 240854 348134 240938
rect 347514 240618 347546 240854
rect 347782 240618 347866 240854
rect 348102 240618 348134 240854
rect 347514 205174 348134 240618
rect 347514 204938 347546 205174
rect 347782 204938 347866 205174
rect 348102 204938 348134 205174
rect 347514 204854 348134 204938
rect 347514 204618 347546 204854
rect 347782 204618 347866 204854
rect 348102 204618 348134 204854
rect 347514 169174 348134 204618
rect 347514 168938 347546 169174
rect 347782 168938 347866 169174
rect 348102 168938 348134 169174
rect 347514 168854 348134 168938
rect 347514 168618 347546 168854
rect 347782 168618 347866 168854
rect 348102 168618 348134 168854
rect 347514 133174 348134 168618
rect 347514 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 348134 133174
rect 347514 132854 348134 132938
rect 347514 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 348134 132854
rect 347514 97174 348134 132618
rect 347514 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 348134 97174
rect 347514 96854 348134 96938
rect 347514 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 348134 96854
rect 347514 61174 348134 96618
rect 347514 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 348134 61174
rect 347514 60854 348134 60938
rect 347514 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 348134 60854
rect 347514 25174 348134 60618
rect 347514 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 348134 25174
rect 347514 24854 348134 24938
rect 347514 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 348134 24854
rect 347514 -3226 348134 24618
rect 347514 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 348134 -3226
rect 347514 -3546 348134 -3462
rect 347514 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 348134 -3546
rect 347514 -3814 348134 -3782
rect 351234 388894 351854 398000
rect 351234 388658 351266 388894
rect 351502 388658 351586 388894
rect 351822 388658 351854 388894
rect 351234 388574 351854 388658
rect 351234 388338 351266 388574
rect 351502 388338 351586 388574
rect 351822 388338 351854 388574
rect 351234 352894 351854 388338
rect 351234 352658 351266 352894
rect 351502 352658 351586 352894
rect 351822 352658 351854 352894
rect 351234 352574 351854 352658
rect 351234 352338 351266 352574
rect 351502 352338 351586 352574
rect 351822 352338 351854 352574
rect 351234 316894 351854 352338
rect 351234 316658 351266 316894
rect 351502 316658 351586 316894
rect 351822 316658 351854 316894
rect 351234 316574 351854 316658
rect 351234 316338 351266 316574
rect 351502 316338 351586 316574
rect 351822 316338 351854 316574
rect 351234 280894 351854 316338
rect 351234 280658 351266 280894
rect 351502 280658 351586 280894
rect 351822 280658 351854 280894
rect 351234 280574 351854 280658
rect 351234 280338 351266 280574
rect 351502 280338 351586 280574
rect 351822 280338 351854 280574
rect 351234 244894 351854 280338
rect 351234 244658 351266 244894
rect 351502 244658 351586 244894
rect 351822 244658 351854 244894
rect 351234 244574 351854 244658
rect 351234 244338 351266 244574
rect 351502 244338 351586 244574
rect 351822 244338 351854 244574
rect 351234 208894 351854 244338
rect 351234 208658 351266 208894
rect 351502 208658 351586 208894
rect 351822 208658 351854 208894
rect 351234 208574 351854 208658
rect 351234 208338 351266 208574
rect 351502 208338 351586 208574
rect 351822 208338 351854 208574
rect 351234 172894 351854 208338
rect 351234 172658 351266 172894
rect 351502 172658 351586 172894
rect 351822 172658 351854 172894
rect 351234 172574 351854 172658
rect 351234 172338 351266 172574
rect 351502 172338 351586 172574
rect 351822 172338 351854 172574
rect 351234 136894 351854 172338
rect 351234 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 351854 136894
rect 351234 136574 351854 136658
rect 351234 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 351854 136574
rect 351234 100894 351854 136338
rect 351234 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 351854 100894
rect 351234 100574 351854 100658
rect 351234 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 351854 100574
rect 351234 64894 351854 100338
rect 351234 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 351854 64894
rect 351234 64574 351854 64658
rect 351234 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 351854 64574
rect 351234 28894 351854 64338
rect 351234 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 351854 28894
rect 351234 28574 351854 28658
rect 351234 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 351854 28574
rect 351234 -5146 351854 28338
rect 351234 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 351854 -5146
rect 351234 -5466 351854 -5382
rect 351234 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 351854 -5466
rect 351234 -5734 351854 -5702
rect 354954 392614 355574 398000
rect 354954 392378 354986 392614
rect 355222 392378 355306 392614
rect 355542 392378 355574 392614
rect 354954 392294 355574 392378
rect 354954 392058 354986 392294
rect 355222 392058 355306 392294
rect 355542 392058 355574 392294
rect 354954 356614 355574 392058
rect 354954 356378 354986 356614
rect 355222 356378 355306 356614
rect 355542 356378 355574 356614
rect 354954 356294 355574 356378
rect 354954 356058 354986 356294
rect 355222 356058 355306 356294
rect 355542 356058 355574 356294
rect 354954 320614 355574 356058
rect 354954 320378 354986 320614
rect 355222 320378 355306 320614
rect 355542 320378 355574 320614
rect 354954 320294 355574 320378
rect 354954 320058 354986 320294
rect 355222 320058 355306 320294
rect 355542 320058 355574 320294
rect 354954 284614 355574 320058
rect 354954 284378 354986 284614
rect 355222 284378 355306 284614
rect 355542 284378 355574 284614
rect 354954 284294 355574 284378
rect 354954 284058 354986 284294
rect 355222 284058 355306 284294
rect 355542 284058 355574 284294
rect 354954 248614 355574 284058
rect 354954 248378 354986 248614
rect 355222 248378 355306 248614
rect 355542 248378 355574 248614
rect 354954 248294 355574 248378
rect 354954 248058 354986 248294
rect 355222 248058 355306 248294
rect 355542 248058 355574 248294
rect 354954 212614 355574 248058
rect 354954 212378 354986 212614
rect 355222 212378 355306 212614
rect 355542 212378 355574 212614
rect 354954 212294 355574 212378
rect 354954 212058 354986 212294
rect 355222 212058 355306 212294
rect 355542 212058 355574 212294
rect 354954 176614 355574 212058
rect 354954 176378 354986 176614
rect 355222 176378 355306 176614
rect 355542 176378 355574 176614
rect 354954 176294 355574 176378
rect 354954 176058 354986 176294
rect 355222 176058 355306 176294
rect 355542 176058 355574 176294
rect 354954 140614 355574 176058
rect 354954 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 355574 140614
rect 354954 140294 355574 140378
rect 354954 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 355574 140294
rect 354954 104614 355574 140058
rect 354954 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 355574 104614
rect 354954 104294 355574 104378
rect 354954 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 355574 104294
rect 354954 68614 355574 104058
rect 354954 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 355574 68614
rect 354954 68294 355574 68378
rect 354954 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 355574 68294
rect 354954 32614 355574 68058
rect 354954 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 355574 32614
rect 354954 32294 355574 32378
rect 354954 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 355574 32294
rect 336954 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 337574 -6106
rect 336954 -6426 337574 -6342
rect 336954 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 337574 -6426
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 32058
rect 361794 363454 362414 398898
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 365514 691174 366134 706202
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 619174 366134 654618
rect 365514 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 366134 619174
rect 365514 618854 366134 618938
rect 365514 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 366134 618854
rect 365514 583174 366134 618618
rect 365514 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 366134 583174
rect 365514 582854 366134 582938
rect 365514 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 366134 582854
rect 365514 547174 366134 582618
rect 365514 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 366134 547174
rect 365514 546854 366134 546938
rect 365514 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 366134 546854
rect 365514 511174 366134 546618
rect 365514 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 366134 511174
rect 365514 510854 366134 510938
rect 365514 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 366134 510854
rect 365514 475174 366134 510618
rect 365514 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 366134 475174
rect 365514 474854 366134 474938
rect 365514 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 366134 474854
rect 365514 439174 366134 474618
rect 365514 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 366134 439174
rect 365514 438854 366134 438938
rect 365514 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 366134 438854
rect 365514 403174 366134 438618
rect 365514 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 366134 403174
rect 365514 402854 366134 402938
rect 365514 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 366134 402854
rect 365514 367174 366134 402618
rect 365514 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 366134 367174
rect 365514 366854 366134 366938
rect 365514 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 366134 366854
rect 365514 331174 366134 366618
rect 365514 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 366134 331174
rect 365514 330854 366134 330938
rect 365514 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 366134 330854
rect 365514 295174 366134 330618
rect 365514 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 366134 295174
rect 365514 294854 366134 294938
rect 365514 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 366134 294854
rect 365514 259174 366134 294618
rect 365514 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 366134 259174
rect 365514 258854 366134 258938
rect 365514 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 366134 258854
rect 365514 223174 366134 258618
rect 365514 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 366134 223174
rect 365514 222854 366134 222938
rect 365514 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 366134 222854
rect 365514 187174 366134 222618
rect 365514 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 366134 187174
rect 365514 186854 366134 186938
rect 365514 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 366134 186854
rect 365514 151174 366134 186618
rect 365514 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 366134 151174
rect 365514 150854 366134 150938
rect 365514 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 366134 150854
rect 365514 115174 366134 150618
rect 365514 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 366134 115174
rect 365514 114854 366134 114938
rect 365514 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 366134 114854
rect 365514 79174 366134 114618
rect 365514 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 366134 79174
rect 365514 78854 366134 78938
rect 365514 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 366134 78854
rect 365514 43174 366134 78618
rect 365514 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 366134 43174
rect 365514 42854 366134 42938
rect 365514 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 366134 42854
rect 365514 7174 366134 42618
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -2266 366134 6618
rect 365514 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 366134 -2266
rect 365514 -2586 366134 -2502
rect 365514 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 366134 -2586
rect 365514 -3814 366134 -2822
rect 369234 694894 369854 708122
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 622894 369854 658338
rect 369234 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 369854 622894
rect 369234 622574 369854 622658
rect 369234 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 369854 622574
rect 369234 586894 369854 622338
rect 369234 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 369854 586894
rect 369234 586574 369854 586658
rect 369234 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 369854 586574
rect 369234 550894 369854 586338
rect 369234 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 369854 550894
rect 369234 550574 369854 550658
rect 369234 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 369854 550574
rect 369234 514894 369854 550338
rect 369234 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 369854 514894
rect 369234 514574 369854 514658
rect 369234 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 369854 514574
rect 369234 478894 369854 514338
rect 369234 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 369854 478894
rect 369234 478574 369854 478658
rect 369234 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 369854 478574
rect 369234 442894 369854 478338
rect 369234 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 369854 442894
rect 369234 442574 369854 442658
rect 369234 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 369854 442574
rect 369234 406894 369854 442338
rect 369234 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 369854 406894
rect 369234 406574 369854 406658
rect 369234 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 369854 406574
rect 369234 370894 369854 406338
rect 369234 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 369854 370894
rect 369234 370574 369854 370658
rect 369234 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 369854 370574
rect 369234 334894 369854 370338
rect 369234 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 369854 334894
rect 369234 334574 369854 334658
rect 369234 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 369854 334574
rect 369234 298894 369854 334338
rect 369234 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 369854 298894
rect 369234 298574 369854 298658
rect 369234 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 369854 298574
rect 369234 262894 369854 298338
rect 369234 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 369854 262894
rect 369234 262574 369854 262658
rect 369234 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 369854 262574
rect 369234 226894 369854 262338
rect 369234 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 369854 226894
rect 369234 226574 369854 226658
rect 369234 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 369854 226574
rect 369234 190894 369854 226338
rect 369234 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 369854 190894
rect 369234 190574 369854 190658
rect 369234 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 369854 190574
rect 369234 154894 369854 190338
rect 369234 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 369854 154894
rect 369234 154574 369854 154658
rect 369234 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 369854 154574
rect 369234 118894 369854 154338
rect 369234 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 369854 118894
rect 369234 118574 369854 118658
rect 369234 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 369854 118574
rect 369234 82894 369854 118338
rect 369234 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 369854 82894
rect 369234 82574 369854 82658
rect 369234 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 369854 82574
rect 369234 46894 369854 82338
rect 369234 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 369854 46894
rect 369234 46574 369854 46658
rect 369234 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 369854 46574
rect 369234 10894 369854 46338
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -4186 369854 10338
rect 369234 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 369854 -4186
rect 369234 -4506 369854 -4422
rect 369234 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 369854 -4506
rect 369234 -5734 369854 -4742
rect 372954 698614 373574 710042
rect 390954 711558 391574 711590
rect 390954 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 391574 711558
rect 390954 711238 391574 711322
rect 390954 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 391574 711238
rect 387234 709638 387854 709670
rect 387234 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 387854 709638
rect 387234 709318 387854 709402
rect 387234 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 387854 709318
rect 383514 707718 384134 707750
rect 383514 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 384134 707718
rect 383514 707398 384134 707482
rect 383514 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 384134 707398
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 626614 373574 662058
rect 372954 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 373574 626614
rect 372954 626294 373574 626378
rect 372954 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 373574 626294
rect 372954 590614 373574 626058
rect 372954 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 373574 590614
rect 372954 590294 373574 590378
rect 372954 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 373574 590294
rect 372954 554614 373574 590058
rect 372954 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 373574 554614
rect 372954 554294 373574 554378
rect 372954 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 373574 554294
rect 372954 518614 373574 554058
rect 372954 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 373574 518614
rect 372954 518294 373574 518378
rect 372954 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 373574 518294
rect 372954 482614 373574 518058
rect 372954 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 373574 482614
rect 372954 482294 373574 482378
rect 372954 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 373574 482294
rect 372954 446614 373574 482058
rect 372954 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 373574 446614
rect 372954 446294 373574 446378
rect 372954 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 373574 446294
rect 372954 410614 373574 446058
rect 372954 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 373574 410614
rect 372954 410294 373574 410378
rect 372954 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 373574 410294
rect 372954 374614 373574 410058
rect 372954 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 373574 374614
rect 372954 374294 373574 374378
rect 372954 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 373574 374294
rect 372954 338614 373574 374058
rect 372954 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 373574 338614
rect 372954 338294 373574 338378
rect 372954 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 373574 338294
rect 372954 302614 373574 338058
rect 372954 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 373574 302614
rect 372954 302294 373574 302378
rect 372954 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 373574 302294
rect 372954 266614 373574 302058
rect 372954 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 373574 266614
rect 372954 266294 373574 266378
rect 372954 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 373574 266294
rect 372954 230614 373574 266058
rect 372954 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 373574 230614
rect 372954 230294 373574 230378
rect 372954 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 373574 230294
rect 372954 194614 373574 230058
rect 372954 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 373574 194614
rect 372954 194294 373574 194378
rect 372954 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 373574 194294
rect 372954 158614 373574 194058
rect 372954 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 373574 158614
rect 372954 158294 373574 158378
rect 372954 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 373574 158294
rect 372954 122614 373574 158058
rect 372954 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 373574 122614
rect 372954 122294 373574 122378
rect 372954 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 373574 122294
rect 372954 86614 373574 122058
rect 372954 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 373574 86614
rect 372954 86294 373574 86378
rect 372954 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 373574 86294
rect 372954 50614 373574 86058
rect 372954 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 373574 50614
rect 372954 50294 373574 50378
rect 372954 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 373574 50294
rect 372954 14614 373574 50058
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 354954 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 355574 -7066
rect 354954 -7386 355574 -7302
rect 354954 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 355574 -7386
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 14058
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 379794 669454 380414 705242
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 417454 380414 452898
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 379794 381454 380414 416898
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 379794 345454 380414 380898
rect 379794 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 380414 345454
rect 379794 345134 380414 345218
rect 379794 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 380414 345134
rect 379794 309454 380414 344898
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 273454 380414 308898
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 237454 380414 272898
rect 379794 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 380414 237454
rect 379794 237134 380414 237218
rect 379794 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 380414 237134
rect 379794 201454 380414 236898
rect 379794 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 380414 201454
rect 379794 201134 380414 201218
rect 379794 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 380414 201134
rect 379794 165454 380414 200898
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 129454 380414 164898
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -1306 380414 20898
rect 379794 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 380414 -1306
rect 379794 -1626 380414 -1542
rect 379794 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 380414 -1626
rect 379794 -1894 380414 -1862
rect 383514 673174 384134 707162
rect 383514 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 384134 673174
rect 383514 672854 384134 672938
rect 383514 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 384134 672854
rect 383514 637174 384134 672618
rect 383514 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 384134 637174
rect 383514 636854 384134 636938
rect 383514 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 384134 636854
rect 383514 601174 384134 636618
rect 383514 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 384134 601174
rect 383514 600854 384134 600938
rect 383514 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 384134 600854
rect 383514 565174 384134 600618
rect 383514 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 384134 565174
rect 383514 564854 384134 564938
rect 383514 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 384134 564854
rect 383514 529174 384134 564618
rect 383514 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 384134 529174
rect 383514 528854 384134 528938
rect 383514 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 384134 528854
rect 383514 493174 384134 528618
rect 383514 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 384134 493174
rect 383514 492854 384134 492938
rect 383514 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 384134 492854
rect 383514 457174 384134 492618
rect 383514 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 384134 457174
rect 383514 456854 384134 456938
rect 383514 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 384134 456854
rect 383514 421174 384134 456618
rect 383514 420938 383546 421174
rect 383782 420938 383866 421174
rect 384102 420938 384134 421174
rect 383514 420854 384134 420938
rect 383514 420618 383546 420854
rect 383782 420618 383866 420854
rect 384102 420618 384134 420854
rect 383514 385174 384134 420618
rect 383514 384938 383546 385174
rect 383782 384938 383866 385174
rect 384102 384938 384134 385174
rect 383514 384854 384134 384938
rect 383514 384618 383546 384854
rect 383782 384618 383866 384854
rect 384102 384618 384134 384854
rect 383514 349174 384134 384618
rect 383514 348938 383546 349174
rect 383782 348938 383866 349174
rect 384102 348938 384134 349174
rect 383514 348854 384134 348938
rect 383514 348618 383546 348854
rect 383782 348618 383866 348854
rect 384102 348618 384134 348854
rect 383514 313174 384134 348618
rect 383514 312938 383546 313174
rect 383782 312938 383866 313174
rect 384102 312938 384134 313174
rect 383514 312854 384134 312938
rect 383514 312618 383546 312854
rect 383782 312618 383866 312854
rect 384102 312618 384134 312854
rect 383514 277174 384134 312618
rect 383514 276938 383546 277174
rect 383782 276938 383866 277174
rect 384102 276938 384134 277174
rect 383514 276854 384134 276938
rect 383514 276618 383546 276854
rect 383782 276618 383866 276854
rect 384102 276618 384134 276854
rect 383514 241174 384134 276618
rect 383514 240938 383546 241174
rect 383782 240938 383866 241174
rect 384102 240938 384134 241174
rect 383514 240854 384134 240938
rect 383514 240618 383546 240854
rect 383782 240618 383866 240854
rect 384102 240618 384134 240854
rect 383514 205174 384134 240618
rect 383514 204938 383546 205174
rect 383782 204938 383866 205174
rect 384102 204938 384134 205174
rect 383514 204854 384134 204938
rect 383514 204618 383546 204854
rect 383782 204618 383866 204854
rect 384102 204618 384134 204854
rect 383514 169174 384134 204618
rect 383514 168938 383546 169174
rect 383782 168938 383866 169174
rect 384102 168938 384134 169174
rect 383514 168854 384134 168938
rect 383514 168618 383546 168854
rect 383782 168618 383866 168854
rect 384102 168618 384134 168854
rect 383514 133174 384134 168618
rect 383514 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 384134 133174
rect 383514 132854 384134 132938
rect 383514 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 384134 132854
rect 383514 97174 384134 132618
rect 383514 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 384134 97174
rect 383514 96854 384134 96938
rect 383514 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 384134 96854
rect 383514 61174 384134 96618
rect 383514 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 384134 61174
rect 383514 60854 384134 60938
rect 383514 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 384134 60854
rect 383514 25174 384134 60618
rect 383514 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 384134 25174
rect 383514 24854 384134 24938
rect 383514 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 384134 24854
rect 383514 -3226 384134 24618
rect 383514 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 384134 -3226
rect 383514 -3546 384134 -3462
rect 383514 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 384134 -3546
rect 383514 -3814 384134 -3782
rect 387234 676894 387854 709082
rect 387234 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 387854 676894
rect 387234 676574 387854 676658
rect 387234 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 387854 676574
rect 387234 640894 387854 676338
rect 387234 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 387854 640894
rect 387234 640574 387854 640658
rect 387234 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 387854 640574
rect 387234 604894 387854 640338
rect 387234 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 387854 604894
rect 387234 604574 387854 604658
rect 387234 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 387854 604574
rect 387234 568894 387854 604338
rect 387234 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 387854 568894
rect 387234 568574 387854 568658
rect 387234 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 387854 568574
rect 387234 532894 387854 568338
rect 387234 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 387854 532894
rect 387234 532574 387854 532658
rect 387234 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 387854 532574
rect 387234 496894 387854 532338
rect 387234 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 387854 496894
rect 387234 496574 387854 496658
rect 387234 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 387854 496574
rect 387234 460894 387854 496338
rect 387234 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 387854 460894
rect 387234 460574 387854 460658
rect 387234 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 387854 460574
rect 387234 424894 387854 460338
rect 387234 424658 387266 424894
rect 387502 424658 387586 424894
rect 387822 424658 387854 424894
rect 387234 424574 387854 424658
rect 387234 424338 387266 424574
rect 387502 424338 387586 424574
rect 387822 424338 387854 424574
rect 387234 388894 387854 424338
rect 387234 388658 387266 388894
rect 387502 388658 387586 388894
rect 387822 388658 387854 388894
rect 387234 388574 387854 388658
rect 387234 388338 387266 388574
rect 387502 388338 387586 388574
rect 387822 388338 387854 388574
rect 387234 352894 387854 388338
rect 387234 352658 387266 352894
rect 387502 352658 387586 352894
rect 387822 352658 387854 352894
rect 387234 352574 387854 352658
rect 387234 352338 387266 352574
rect 387502 352338 387586 352574
rect 387822 352338 387854 352574
rect 387234 316894 387854 352338
rect 387234 316658 387266 316894
rect 387502 316658 387586 316894
rect 387822 316658 387854 316894
rect 387234 316574 387854 316658
rect 387234 316338 387266 316574
rect 387502 316338 387586 316574
rect 387822 316338 387854 316574
rect 387234 280894 387854 316338
rect 387234 280658 387266 280894
rect 387502 280658 387586 280894
rect 387822 280658 387854 280894
rect 387234 280574 387854 280658
rect 387234 280338 387266 280574
rect 387502 280338 387586 280574
rect 387822 280338 387854 280574
rect 387234 244894 387854 280338
rect 387234 244658 387266 244894
rect 387502 244658 387586 244894
rect 387822 244658 387854 244894
rect 387234 244574 387854 244658
rect 387234 244338 387266 244574
rect 387502 244338 387586 244574
rect 387822 244338 387854 244574
rect 387234 208894 387854 244338
rect 387234 208658 387266 208894
rect 387502 208658 387586 208894
rect 387822 208658 387854 208894
rect 387234 208574 387854 208658
rect 387234 208338 387266 208574
rect 387502 208338 387586 208574
rect 387822 208338 387854 208574
rect 387234 172894 387854 208338
rect 387234 172658 387266 172894
rect 387502 172658 387586 172894
rect 387822 172658 387854 172894
rect 387234 172574 387854 172658
rect 387234 172338 387266 172574
rect 387502 172338 387586 172574
rect 387822 172338 387854 172574
rect 387234 136894 387854 172338
rect 387234 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 387854 136894
rect 387234 136574 387854 136658
rect 387234 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 387854 136574
rect 387234 100894 387854 136338
rect 387234 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 387854 100894
rect 387234 100574 387854 100658
rect 387234 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 387854 100574
rect 387234 64894 387854 100338
rect 387234 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 387854 64894
rect 387234 64574 387854 64658
rect 387234 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 387854 64574
rect 387234 28894 387854 64338
rect 387234 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 387854 28894
rect 387234 28574 387854 28658
rect 387234 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 387854 28574
rect 387234 -5146 387854 28338
rect 387234 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 387854 -5146
rect 387234 -5466 387854 -5382
rect 387234 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 387854 -5466
rect 387234 -5734 387854 -5702
rect 390954 680614 391574 711002
rect 408954 710598 409574 711590
rect 408954 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 409574 710598
rect 408954 710278 409574 710362
rect 408954 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 409574 710278
rect 405234 708678 405854 709670
rect 405234 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 405854 708678
rect 405234 708358 405854 708442
rect 405234 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 405854 708358
rect 401514 706758 402134 707750
rect 401514 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 402134 706758
rect 401514 706438 402134 706522
rect 401514 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 402134 706438
rect 390954 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 391574 680614
rect 390954 680294 391574 680378
rect 390954 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 391574 680294
rect 390954 644614 391574 680058
rect 390954 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 391574 644614
rect 390954 644294 391574 644378
rect 390954 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 391574 644294
rect 390954 608614 391574 644058
rect 390954 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 391574 608614
rect 390954 608294 391574 608378
rect 390954 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 391574 608294
rect 390954 572614 391574 608058
rect 390954 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 391574 572614
rect 390954 572294 391574 572378
rect 390954 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 391574 572294
rect 390954 536614 391574 572058
rect 390954 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 391574 536614
rect 390954 536294 391574 536378
rect 390954 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 391574 536294
rect 390954 500614 391574 536058
rect 390954 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 391574 500614
rect 390954 500294 391574 500378
rect 390954 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 391574 500294
rect 390954 464614 391574 500058
rect 390954 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 391574 464614
rect 390954 464294 391574 464378
rect 390954 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 391574 464294
rect 390954 428614 391574 464058
rect 390954 428378 390986 428614
rect 391222 428378 391306 428614
rect 391542 428378 391574 428614
rect 390954 428294 391574 428378
rect 390954 428058 390986 428294
rect 391222 428058 391306 428294
rect 391542 428058 391574 428294
rect 390954 392614 391574 428058
rect 390954 392378 390986 392614
rect 391222 392378 391306 392614
rect 391542 392378 391574 392614
rect 390954 392294 391574 392378
rect 390954 392058 390986 392294
rect 391222 392058 391306 392294
rect 391542 392058 391574 392294
rect 390954 356614 391574 392058
rect 390954 356378 390986 356614
rect 391222 356378 391306 356614
rect 391542 356378 391574 356614
rect 390954 356294 391574 356378
rect 390954 356058 390986 356294
rect 391222 356058 391306 356294
rect 391542 356058 391574 356294
rect 390954 320614 391574 356058
rect 390954 320378 390986 320614
rect 391222 320378 391306 320614
rect 391542 320378 391574 320614
rect 390954 320294 391574 320378
rect 390954 320058 390986 320294
rect 391222 320058 391306 320294
rect 391542 320058 391574 320294
rect 390954 284614 391574 320058
rect 390954 284378 390986 284614
rect 391222 284378 391306 284614
rect 391542 284378 391574 284614
rect 390954 284294 391574 284378
rect 390954 284058 390986 284294
rect 391222 284058 391306 284294
rect 391542 284058 391574 284294
rect 390954 248614 391574 284058
rect 390954 248378 390986 248614
rect 391222 248378 391306 248614
rect 391542 248378 391574 248614
rect 390954 248294 391574 248378
rect 390954 248058 390986 248294
rect 391222 248058 391306 248294
rect 391542 248058 391574 248294
rect 390954 212614 391574 248058
rect 390954 212378 390986 212614
rect 391222 212378 391306 212614
rect 391542 212378 391574 212614
rect 390954 212294 391574 212378
rect 390954 212058 390986 212294
rect 391222 212058 391306 212294
rect 391542 212058 391574 212294
rect 390954 176614 391574 212058
rect 390954 176378 390986 176614
rect 391222 176378 391306 176614
rect 391542 176378 391574 176614
rect 390954 176294 391574 176378
rect 390954 176058 390986 176294
rect 391222 176058 391306 176294
rect 391542 176058 391574 176294
rect 390954 140614 391574 176058
rect 390954 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 391574 140614
rect 390954 140294 391574 140378
rect 390954 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 391574 140294
rect 390954 104614 391574 140058
rect 390954 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 391574 104614
rect 390954 104294 391574 104378
rect 390954 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 391574 104294
rect 390954 68614 391574 104058
rect 390954 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 391574 68614
rect 390954 68294 391574 68378
rect 390954 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 391574 68294
rect 390954 32614 391574 68058
rect 390954 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 391574 32614
rect 390954 32294 391574 32378
rect 390954 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 391574 32294
rect 372954 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 373574 -6106
rect 372954 -6426 373574 -6342
rect 372954 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 373574 -6426
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 32058
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 401514 691174 402134 706202
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 619174 402134 654618
rect 401514 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 402134 619174
rect 401514 618854 402134 618938
rect 401514 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 402134 618854
rect 401514 583174 402134 618618
rect 401514 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 402134 583174
rect 401514 582854 402134 582938
rect 401514 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 402134 582854
rect 401514 547174 402134 582618
rect 401514 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 402134 547174
rect 401514 546854 402134 546938
rect 401514 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 402134 546854
rect 401514 511174 402134 546618
rect 401514 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 402134 511174
rect 401514 510854 402134 510938
rect 401514 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 402134 510854
rect 401514 475174 402134 510618
rect 401514 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 402134 475174
rect 401514 474854 402134 474938
rect 401514 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 402134 474854
rect 401514 439174 402134 474618
rect 401514 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 402134 439174
rect 401514 438854 402134 438938
rect 401514 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 402134 438854
rect 401514 403174 402134 438618
rect 401514 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 402134 403174
rect 401514 402854 402134 402938
rect 401514 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 402134 402854
rect 401514 367174 402134 402618
rect 401514 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 402134 367174
rect 401514 366854 402134 366938
rect 401514 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 402134 366854
rect 401514 331174 402134 366618
rect 401514 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 402134 331174
rect 401514 330854 402134 330938
rect 401514 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 402134 330854
rect 401514 295174 402134 330618
rect 401514 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 402134 295174
rect 401514 294854 402134 294938
rect 401514 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 402134 294854
rect 401514 259174 402134 294618
rect 401514 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 402134 259174
rect 401514 258854 402134 258938
rect 401514 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 402134 258854
rect 401514 223174 402134 258618
rect 401514 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 402134 223174
rect 401514 222854 402134 222938
rect 401514 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 402134 222854
rect 401514 187174 402134 222618
rect 401514 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 402134 187174
rect 401514 186854 402134 186938
rect 401514 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 402134 186854
rect 401514 151174 402134 186618
rect 401514 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 402134 151174
rect 401514 150854 402134 150938
rect 401514 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 402134 150854
rect 401514 115174 402134 150618
rect 401514 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 402134 115174
rect 401514 114854 402134 114938
rect 401514 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 402134 114854
rect 401514 79174 402134 114618
rect 401514 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 402134 79174
rect 401514 78854 402134 78938
rect 401514 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 402134 78854
rect 401514 43174 402134 78618
rect 401514 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 402134 43174
rect 401514 42854 402134 42938
rect 401514 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 402134 42854
rect 401514 7174 402134 42618
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -2266 402134 6618
rect 401514 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 402134 -2266
rect 401514 -2586 402134 -2502
rect 401514 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 402134 -2586
rect 401514 -3814 402134 -2822
rect 405234 694894 405854 708122
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 658894 405854 694338
rect 405234 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 405854 658894
rect 405234 658574 405854 658658
rect 405234 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 405854 658574
rect 405234 622894 405854 658338
rect 405234 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 405854 622894
rect 405234 622574 405854 622658
rect 405234 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 405854 622574
rect 405234 586894 405854 622338
rect 405234 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 405854 586894
rect 405234 586574 405854 586658
rect 405234 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 405854 586574
rect 405234 550894 405854 586338
rect 405234 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 405854 550894
rect 405234 550574 405854 550658
rect 405234 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 405854 550574
rect 405234 514894 405854 550338
rect 405234 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 405854 514894
rect 405234 514574 405854 514658
rect 405234 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 405854 514574
rect 405234 478894 405854 514338
rect 405234 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 405854 478894
rect 405234 478574 405854 478658
rect 405234 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 405854 478574
rect 405234 442894 405854 478338
rect 405234 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 405854 442894
rect 405234 442574 405854 442658
rect 405234 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 405854 442574
rect 405234 406894 405854 442338
rect 405234 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 405854 406894
rect 405234 406574 405854 406658
rect 405234 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 405854 406574
rect 405234 370894 405854 406338
rect 405234 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 405854 370894
rect 405234 370574 405854 370658
rect 405234 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 405854 370574
rect 405234 334894 405854 370338
rect 405234 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 405854 334894
rect 405234 334574 405854 334658
rect 405234 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 405854 334574
rect 405234 298894 405854 334338
rect 405234 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 405854 298894
rect 405234 298574 405854 298658
rect 405234 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 405854 298574
rect 405234 262894 405854 298338
rect 405234 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 405854 262894
rect 405234 262574 405854 262658
rect 405234 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 405854 262574
rect 405234 226894 405854 262338
rect 405234 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 405854 226894
rect 405234 226574 405854 226658
rect 405234 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 405854 226574
rect 405234 190894 405854 226338
rect 405234 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 405854 190894
rect 405234 190574 405854 190658
rect 405234 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 405854 190574
rect 405234 154894 405854 190338
rect 405234 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 405854 154894
rect 405234 154574 405854 154658
rect 405234 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 405854 154574
rect 405234 118894 405854 154338
rect 405234 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 405854 118894
rect 405234 118574 405854 118658
rect 405234 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 405854 118574
rect 405234 82894 405854 118338
rect 405234 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 405854 82894
rect 405234 82574 405854 82658
rect 405234 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 405854 82574
rect 405234 46894 405854 82338
rect 405234 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 405854 46894
rect 405234 46574 405854 46658
rect 405234 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 405854 46574
rect 405234 10894 405854 46338
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -4186 405854 10338
rect 405234 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 405854 -4186
rect 405234 -4506 405854 -4422
rect 405234 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 405854 -4506
rect 405234 -5734 405854 -4742
rect 408954 698614 409574 710042
rect 426954 711558 427574 711590
rect 426954 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 427574 711558
rect 426954 711238 427574 711322
rect 426954 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 427574 711238
rect 423234 709638 423854 709670
rect 423234 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 423854 709638
rect 423234 709318 423854 709402
rect 423234 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 423854 709318
rect 419514 707718 420134 707750
rect 419514 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 420134 707718
rect 419514 707398 420134 707482
rect 419514 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 420134 707398
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 626614 409574 662058
rect 408954 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 409574 626614
rect 408954 626294 409574 626378
rect 408954 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 409574 626294
rect 408954 590614 409574 626058
rect 408954 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 409574 590614
rect 408954 590294 409574 590378
rect 408954 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 409574 590294
rect 408954 554614 409574 590058
rect 408954 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 409574 554614
rect 408954 554294 409574 554378
rect 408954 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 409574 554294
rect 408954 518614 409574 554058
rect 408954 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 409574 518614
rect 408954 518294 409574 518378
rect 408954 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 409574 518294
rect 408954 482614 409574 518058
rect 408954 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 409574 482614
rect 408954 482294 409574 482378
rect 408954 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 409574 482294
rect 408954 446614 409574 482058
rect 408954 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 409574 446614
rect 408954 446294 409574 446378
rect 408954 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 409574 446294
rect 408954 410614 409574 446058
rect 408954 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 409574 410614
rect 408954 410294 409574 410378
rect 408954 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 409574 410294
rect 408954 374614 409574 410058
rect 408954 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 409574 374614
rect 408954 374294 409574 374378
rect 408954 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 409574 374294
rect 408954 338614 409574 374058
rect 408954 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 409574 338614
rect 408954 338294 409574 338378
rect 408954 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 409574 338294
rect 408954 302614 409574 338058
rect 408954 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 409574 302614
rect 408954 302294 409574 302378
rect 408954 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 409574 302294
rect 408954 266614 409574 302058
rect 408954 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 409574 266614
rect 408954 266294 409574 266378
rect 408954 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 409574 266294
rect 408954 230614 409574 266058
rect 408954 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 409574 230614
rect 408954 230294 409574 230378
rect 408954 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 409574 230294
rect 408954 194614 409574 230058
rect 408954 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 409574 194614
rect 408954 194294 409574 194378
rect 408954 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 409574 194294
rect 408954 158614 409574 194058
rect 408954 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 409574 158614
rect 408954 158294 409574 158378
rect 408954 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 409574 158294
rect 408954 122614 409574 158058
rect 408954 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 409574 122614
rect 408954 122294 409574 122378
rect 408954 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 409574 122294
rect 408954 86614 409574 122058
rect 408954 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 409574 86614
rect 408954 86294 409574 86378
rect 408954 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 409574 86294
rect 408954 50614 409574 86058
rect 408954 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 409574 50614
rect 408954 50294 409574 50378
rect 408954 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 409574 50294
rect 408954 14614 409574 50058
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 390954 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 391574 -7066
rect 390954 -7386 391574 -7302
rect 390954 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 391574 -7386
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 14058
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 415794 669454 416414 705242
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 381454 416414 416898
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 273454 416414 308898
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 415794 237454 416414 272898
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 129454 416414 164898
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -1306 416414 20898
rect 415794 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 416414 -1306
rect 415794 -1626 416414 -1542
rect 415794 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 416414 -1626
rect 415794 -1894 416414 -1862
rect 419514 673174 420134 707162
rect 419514 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 420134 673174
rect 419514 672854 420134 672938
rect 419514 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 420134 672854
rect 419514 637174 420134 672618
rect 419514 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 420134 637174
rect 419514 636854 420134 636938
rect 419514 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 420134 636854
rect 419514 601174 420134 636618
rect 419514 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 420134 601174
rect 419514 600854 420134 600938
rect 419514 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 420134 600854
rect 419514 565174 420134 600618
rect 419514 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 420134 565174
rect 419514 564854 420134 564938
rect 419514 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 420134 564854
rect 419514 529174 420134 564618
rect 419514 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 420134 529174
rect 419514 528854 420134 528938
rect 419514 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 420134 528854
rect 419514 493174 420134 528618
rect 419514 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 420134 493174
rect 419514 492854 420134 492938
rect 419514 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 420134 492854
rect 419514 457174 420134 492618
rect 419514 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 420134 457174
rect 419514 456854 420134 456938
rect 419514 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 420134 456854
rect 419514 421174 420134 456618
rect 419514 420938 419546 421174
rect 419782 420938 419866 421174
rect 420102 420938 420134 421174
rect 419514 420854 420134 420938
rect 419514 420618 419546 420854
rect 419782 420618 419866 420854
rect 420102 420618 420134 420854
rect 419514 385174 420134 420618
rect 419514 384938 419546 385174
rect 419782 384938 419866 385174
rect 420102 384938 420134 385174
rect 419514 384854 420134 384938
rect 419514 384618 419546 384854
rect 419782 384618 419866 384854
rect 420102 384618 420134 384854
rect 419514 349174 420134 384618
rect 419514 348938 419546 349174
rect 419782 348938 419866 349174
rect 420102 348938 420134 349174
rect 419514 348854 420134 348938
rect 419514 348618 419546 348854
rect 419782 348618 419866 348854
rect 420102 348618 420134 348854
rect 419514 313174 420134 348618
rect 419514 312938 419546 313174
rect 419782 312938 419866 313174
rect 420102 312938 420134 313174
rect 419514 312854 420134 312938
rect 419514 312618 419546 312854
rect 419782 312618 419866 312854
rect 420102 312618 420134 312854
rect 419514 277174 420134 312618
rect 419514 276938 419546 277174
rect 419782 276938 419866 277174
rect 420102 276938 420134 277174
rect 419514 276854 420134 276938
rect 419514 276618 419546 276854
rect 419782 276618 419866 276854
rect 420102 276618 420134 276854
rect 419514 241174 420134 276618
rect 419514 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 420134 241174
rect 419514 240854 420134 240938
rect 419514 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 420134 240854
rect 419514 205174 420134 240618
rect 419514 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 420134 205174
rect 419514 204854 420134 204938
rect 419514 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 420134 204854
rect 419514 169174 420134 204618
rect 419514 168938 419546 169174
rect 419782 168938 419866 169174
rect 420102 168938 420134 169174
rect 419514 168854 420134 168938
rect 419514 168618 419546 168854
rect 419782 168618 419866 168854
rect 420102 168618 420134 168854
rect 419514 133174 420134 168618
rect 419514 132938 419546 133174
rect 419782 132938 419866 133174
rect 420102 132938 420134 133174
rect 419514 132854 420134 132938
rect 419514 132618 419546 132854
rect 419782 132618 419866 132854
rect 420102 132618 420134 132854
rect 419514 97174 420134 132618
rect 419514 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 420134 97174
rect 419514 96854 420134 96938
rect 419514 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 420134 96854
rect 419514 61174 420134 96618
rect 419514 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 420134 61174
rect 419514 60854 420134 60938
rect 419514 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 420134 60854
rect 419514 25174 420134 60618
rect 419514 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 420134 25174
rect 419514 24854 420134 24938
rect 419514 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 420134 24854
rect 419514 -3226 420134 24618
rect 419514 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 420134 -3226
rect 419514 -3546 420134 -3462
rect 419514 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 420134 -3546
rect 419514 -3814 420134 -3782
rect 423234 676894 423854 709082
rect 423234 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 423854 676894
rect 423234 676574 423854 676658
rect 423234 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 423854 676574
rect 423234 640894 423854 676338
rect 423234 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 423854 640894
rect 423234 640574 423854 640658
rect 423234 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 423854 640574
rect 423234 604894 423854 640338
rect 423234 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 423854 604894
rect 423234 604574 423854 604658
rect 423234 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 423854 604574
rect 423234 568894 423854 604338
rect 423234 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 423854 568894
rect 423234 568574 423854 568658
rect 423234 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 423854 568574
rect 423234 532894 423854 568338
rect 423234 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 423854 532894
rect 423234 532574 423854 532658
rect 423234 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 423854 532574
rect 423234 496894 423854 532338
rect 423234 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 423854 496894
rect 423234 496574 423854 496658
rect 423234 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 423854 496574
rect 423234 460894 423854 496338
rect 423234 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 423854 460894
rect 423234 460574 423854 460658
rect 423234 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 423854 460574
rect 423234 424894 423854 460338
rect 423234 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 423854 424894
rect 423234 424574 423854 424658
rect 423234 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 423854 424574
rect 423234 388894 423854 424338
rect 423234 388658 423266 388894
rect 423502 388658 423586 388894
rect 423822 388658 423854 388894
rect 423234 388574 423854 388658
rect 423234 388338 423266 388574
rect 423502 388338 423586 388574
rect 423822 388338 423854 388574
rect 423234 352894 423854 388338
rect 423234 352658 423266 352894
rect 423502 352658 423586 352894
rect 423822 352658 423854 352894
rect 423234 352574 423854 352658
rect 423234 352338 423266 352574
rect 423502 352338 423586 352574
rect 423822 352338 423854 352574
rect 423234 316894 423854 352338
rect 423234 316658 423266 316894
rect 423502 316658 423586 316894
rect 423822 316658 423854 316894
rect 423234 316574 423854 316658
rect 423234 316338 423266 316574
rect 423502 316338 423586 316574
rect 423822 316338 423854 316574
rect 423234 280894 423854 316338
rect 423234 280658 423266 280894
rect 423502 280658 423586 280894
rect 423822 280658 423854 280894
rect 423234 280574 423854 280658
rect 423234 280338 423266 280574
rect 423502 280338 423586 280574
rect 423822 280338 423854 280574
rect 423234 244894 423854 280338
rect 423234 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 423854 244894
rect 423234 244574 423854 244658
rect 423234 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 423854 244574
rect 423234 208894 423854 244338
rect 423234 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 423854 208894
rect 423234 208574 423854 208658
rect 423234 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 423854 208574
rect 423234 172894 423854 208338
rect 423234 172658 423266 172894
rect 423502 172658 423586 172894
rect 423822 172658 423854 172894
rect 423234 172574 423854 172658
rect 423234 172338 423266 172574
rect 423502 172338 423586 172574
rect 423822 172338 423854 172574
rect 423234 136894 423854 172338
rect 423234 136658 423266 136894
rect 423502 136658 423586 136894
rect 423822 136658 423854 136894
rect 423234 136574 423854 136658
rect 423234 136338 423266 136574
rect 423502 136338 423586 136574
rect 423822 136338 423854 136574
rect 423234 100894 423854 136338
rect 423234 100658 423266 100894
rect 423502 100658 423586 100894
rect 423822 100658 423854 100894
rect 423234 100574 423854 100658
rect 423234 100338 423266 100574
rect 423502 100338 423586 100574
rect 423822 100338 423854 100574
rect 423234 64894 423854 100338
rect 423234 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 423854 64894
rect 423234 64574 423854 64658
rect 423234 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 423854 64574
rect 423234 28894 423854 64338
rect 423234 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 423854 28894
rect 423234 28574 423854 28658
rect 423234 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 423854 28574
rect 423234 -5146 423854 28338
rect 423234 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 423854 -5146
rect 423234 -5466 423854 -5382
rect 423234 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 423854 -5466
rect 423234 -5734 423854 -5702
rect 426954 680614 427574 711002
rect 444954 710598 445574 711590
rect 444954 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 445574 710598
rect 444954 710278 445574 710362
rect 444954 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 445574 710278
rect 441234 708678 441854 709670
rect 441234 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 441854 708678
rect 441234 708358 441854 708442
rect 441234 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 441854 708358
rect 437514 706758 438134 707750
rect 437514 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 438134 706758
rect 437514 706438 438134 706522
rect 437514 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 438134 706438
rect 426954 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 427574 680614
rect 426954 680294 427574 680378
rect 426954 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 427574 680294
rect 426954 644614 427574 680058
rect 426954 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 427574 644614
rect 426954 644294 427574 644378
rect 426954 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 427574 644294
rect 426954 608614 427574 644058
rect 426954 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 427574 608614
rect 426954 608294 427574 608378
rect 426954 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 427574 608294
rect 426954 572614 427574 608058
rect 426954 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 427574 572614
rect 426954 572294 427574 572378
rect 426954 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 427574 572294
rect 426954 536614 427574 572058
rect 426954 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 427574 536614
rect 426954 536294 427574 536378
rect 426954 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 427574 536294
rect 426954 500614 427574 536058
rect 426954 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 427574 500614
rect 426954 500294 427574 500378
rect 426954 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 427574 500294
rect 426954 464614 427574 500058
rect 426954 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 427574 464614
rect 426954 464294 427574 464378
rect 426954 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 427574 464294
rect 426954 428614 427574 464058
rect 426954 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 427574 428614
rect 426954 428294 427574 428378
rect 426954 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 427574 428294
rect 426954 392614 427574 428058
rect 426954 392378 426986 392614
rect 427222 392378 427306 392614
rect 427542 392378 427574 392614
rect 426954 392294 427574 392378
rect 426954 392058 426986 392294
rect 427222 392058 427306 392294
rect 427542 392058 427574 392294
rect 426954 356614 427574 392058
rect 426954 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 427574 356614
rect 426954 356294 427574 356378
rect 426954 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 427574 356294
rect 426954 320614 427574 356058
rect 426954 320378 426986 320614
rect 427222 320378 427306 320614
rect 427542 320378 427574 320614
rect 426954 320294 427574 320378
rect 426954 320058 426986 320294
rect 427222 320058 427306 320294
rect 427542 320058 427574 320294
rect 426954 284614 427574 320058
rect 426954 284378 426986 284614
rect 427222 284378 427306 284614
rect 427542 284378 427574 284614
rect 426954 284294 427574 284378
rect 426954 284058 426986 284294
rect 427222 284058 427306 284294
rect 427542 284058 427574 284294
rect 426954 248614 427574 284058
rect 426954 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 427574 248614
rect 426954 248294 427574 248378
rect 426954 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 427574 248294
rect 426954 212614 427574 248058
rect 426954 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 427574 212614
rect 426954 212294 427574 212378
rect 426954 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 427574 212294
rect 426954 176614 427574 212058
rect 426954 176378 426986 176614
rect 427222 176378 427306 176614
rect 427542 176378 427574 176614
rect 426954 176294 427574 176378
rect 426954 176058 426986 176294
rect 427222 176058 427306 176294
rect 427542 176058 427574 176294
rect 426954 140614 427574 176058
rect 426954 140378 426986 140614
rect 427222 140378 427306 140614
rect 427542 140378 427574 140614
rect 426954 140294 427574 140378
rect 426954 140058 426986 140294
rect 427222 140058 427306 140294
rect 427542 140058 427574 140294
rect 426954 104614 427574 140058
rect 426954 104378 426986 104614
rect 427222 104378 427306 104614
rect 427542 104378 427574 104614
rect 426954 104294 427574 104378
rect 426954 104058 426986 104294
rect 427222 104058 427306 104294
rect 427542 104058 427574 104294
rect 426954 68614 427574 104058
rect 426954 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 427574 68614
rect 426954 68294 427574 68378
rect 426954 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 427574 68294
rect 426954 32614 427574 68058
rect 426954 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 427574 32614
rect 426954 32294 427574 32378
rect 426954 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 427574 32294
rect 408954 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 409574 -6106
rect 408954 -6426 409574 -6342
rect 408954 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 409574 -6426
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 32058
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 437514 691174 438134 706202
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 655174 438134 690618
rect 437514 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 438134 655174
rect 437514 654854 438134 654938
rect 437514 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 438134 654854
rect 437514 619174 438134 654618
rect 437514 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 438134 619174
rect 437514 618854 438134 618938
rect 437514 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 438134 618854
rect 437514 583174 438134 618618
rect 437514 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 438134 583174
rect 437514 582854 438134 582938
rect 437514 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 438134 582854
rect 437514 547174 438134 582618
rect 437514 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 438134 547174
rect 437514 546854 438134 546938
rect 437514 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 438134 546854
rect 437514 511174 438134 546618
rect 437514 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 438134 511174
rect 437514 510854 438134 510938
rect 437514 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 438134 510854
rect 437514 475174 438134 510618
rect 437514 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 438134 475174
rect 437514 474854 438134 474938
rect 437514 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 438134 474854
rect 437514 439174 438134 474618
rect 437514 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 438134 439174
rect 437514 438854 438134 438938
rect 437514 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 438134 438854
rect 437514 403174 438134 438618
rect 437514 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 438134 403174
rect 437514 402854 438134 402938
rect 437514 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 438134 402854
rect 437514 367174 438134 402618
rect 437514 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 438134 367174
rect 437514 366854 438134 366938
rect 437514 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 438134 366854
rect 437514 331174 438134 366618
rect 437514 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 438134 331174
rect 437514 330854 438134 330938
rect 437514 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 438134 330854
rect 437514 295174 438134 330618
rect 437514 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 438134 295174
rect 437514 294854 438134 294938
rect 437514 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 438134 294854
rect 437514 259174 438134 294618
rect 437514 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 438134 259174
rect 437514 258854 438134 258938
rect 437514 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 438134 258854
rect 437514 223174 438134 258618
rect 437514 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 438134 223174
rect 437514 222854 438134 222938
rect 437514 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 438134 222854
rect 437514 187174 438134 222618
rect 437514 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 438134 187174
rect 437514 186854 438134 186938
rect 437514 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 438134 186854
rect 437514 151174 438134 186618
rect 437514 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 438134 151174
rect 437514 150854 438134 150938
rect 437514 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 438134 150854
rect 437514 115174 438134 150618
rect 437514 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 438134 115174
rect 437514 114854 438134 114938
rect 437514 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 438134 114854
rect 437514 79174 438134 114618
rect 437514 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 438134 79174
rect 437514 78854 438134 78938
rect 437514 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 438134 78854
rect 437514 43174 438134 78618
rect 437514 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 438134 43174
rect 437514 42854 438134 42938
rect 437514 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 438134 42854
rect 437514 7174 438134 42618
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -2266 438134 6618
rect 437514 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 438134 -2266
rect 437514 -2586 438134 -2502
rect 437514 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 438134 -2586
rect 437514 -3814 438134 -2822
rect 441234 694894 441854 708122
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 658894 441854 694338
rect 441234 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 441854 658894
rect 441234 658574 441854 658658
rect 441234 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 441854 658574
rect 441234 622894 441854 658338
rect 441234 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 441854 622894
rect 441234 622574 441854 622658
rect 441234 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 441854 622574
rect 441234 586894 441854 622338
rect 441234 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 441854 586894
rect 441234 586574 441854 586658
rect 441234 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 441854 586574
rect 441234 550894 441854 586338
rect 441234 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 441854 550894
rect 441234 550574 441854 550658
rect 441234 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 441854 550574
rect 441234 514894 441854 550338
rect 441234 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 441854 514894
rect 441234 514574 441854 514658
rect 441234 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 441854 514574
rect 441234 478894 441854 514338
rect 441234 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 441854 478894
rect 441234 478574 441854 478658
rect 441234 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 441854 478574
rect 441234 442894 441854 478338
rect 441234 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 441854 442894
rect 441234 442574 441854 442658
rect 441234 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 441854 442574
rect 441234 406894 441854 442338
rect 441234 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 441854 406894
rect 441234 406574 441854 406658
rect 441234 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 441854 406574
rect 441234 370894 441854 406338
rect 441234 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 441854 370894
rect 441234 370574 441854 370658
rect 441234 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 441854 370574
rect 441234 334894 441854 370338
rect 441234 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 441854 334894
rect 441234 334574 441854 334658
rect 441234 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 441854 334574
rect 441234 298894 441854 334338
rect 441234 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 441854 298894
rect 441234 298574 441854 298658
rect 441234 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 441854 298574
rect 441234 262894 441854 298338
rect 441234 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 441854 262894
rect 441234 262574 441854 262658
rect 441234 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 441854 262574
rect 441234 226894 441854 262338
rect 441234 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 441854 226894
rect 441234 226574 441854 226658
rect 441234 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 441854 226574
rect 441234 190894 441854 226338
rect 441234 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 441854 190894
rect 441234 190574 441854 190658
rect 441234 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 441854 190574
rect 441234 154894 441854 190338
rect 441234 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 441854 154894
rect 441234 154574 441854 154658
rect 441234 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 441854 154574
rect 441234 118894 441854 154338
rect 441234 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 441854 118894
rect 441234 118574 441854 118658
rect 441234 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 441854 118574
rect 441234 82894 441854 118338
rect 441234 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 441854 82894
rect 441234 82574 441854 82658
rect 441234 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 441854 82574
rect 441234 46894 441854 82338
rect 441234 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 441854 46894
rect 441234 46574 441854 46658
rect 441234 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 441854 46574
rect 441234 10894 441854 46338
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -4186 441854 10338
rect 441234 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 441854 -4186
rect 441234 -4506 441854 -4422
rect 441234 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 441854 -4506
rect 441234 -5734 441854 -4742
rect 444954 698614 445574 710042
rect 462954 711558 463574 711590
rect 462954 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 463574 711558
rect 462954 711238 463574 711322
rect 462954 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 463574 711238
rect 459234 709638 459854 709670
rect 459234 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 459854 709638
rect 459234 709318 459854 709402
rect 459234 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 459854 709318
rect 455514 707718 456134 707750
rect 455514 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 456134 707718
rect 455514 707398 456134 707482
rect 455514 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 456134 707398
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 662614 445574 698058
rect 444954 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 445574 662614
rect 444954 662294 445574 662378
rect 444954 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 445574 662294
rect 444954 626614 445574 662058
rect 444954 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 445574 626614
rect 444954 626294 445574 626378
rect 444954 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 445574 626294
rect 444954 590614 445574 626058
rect 444954 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 445574 590614
rect 444954 590294 445574 590378
rect 444954 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 445574 590294
rect 444954 554614 445574 590058
rect 444954 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 445574 554614
rect 444954 554294 445574 554378
rect 444954 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 445574 554294
rect 444954 518614 445574 554058
rect 444954 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 445574 518614
rect 444954 518294 445574 518378
rect 444954 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 445574 518294
rect 444954 482614 445574 518058
rect 444954 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 445574 482614
rect 444954 482294 445574 482378
rect 444954 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 445574 482294
rect 444954 446614 445574 482058
rect 444954 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 445574 446614
rect 444954 446294 445574 446378
rect 444954 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 445574 446294
rect 444954 410614 445574 446058
rect 444954 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 445574 410614
rect 444954 410294 445574 410378
rect 444954 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 445574 410294
rect 444954 374614 445574 410058
rect 444954 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 445574 374614
rect 444954 374294 445574 374378
rect 444954 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 445574 374294
rect 444954 338614 445574 374058
rect 444954 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 445574 338614
rect 444954 338294 445574 338378
rect 444954 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 445574 338294
rect 444954 302614 445574 338058
rect 444954 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 445574 302614
rect 444954 302294 445574 302378
rect 444954 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 445574 302294
rect 444954 266614 445574 302058
rect 444954 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 445574 266614
rect 444954 266294 445574 266378
rect 444954 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 445574 266294
rect 444954 230614 445574 266058
rect 444954 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 445574 230614
rect 444954 230294 445574 230378
rect 444954 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 445574 230294
rect 444954 194614 445574 230058
rect 444954 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 445574 194614
rect 444954 194294 445574 194378
rect 444954 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 445574 194294
rect 444954 158614 445574 194058
rect 444954 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 445574 158614
rect 444954 158294 445574 158378
rect 444954 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 445574 158294
rect 444954 122614 445574 158058
rect 444954 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 445574 122614
rect 444954 122294 445574 122378
rect 444954 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 445574 122294
rect 444954 86614 445574 122058
rect 444954 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 445574 86614
rect 444954 86294 445574 86378
rect 444954 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 445574 86294
rect 444954 50614 445574 86058
rect 444954 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 445574 50614
rect 444954 50294 445574 50378
rect 444954 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 445574 50294
rect 444954 14614 445574 50058
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 426954 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 427574 -7066
rect 426954 -7386 427574 -7302
rect 426954 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 427574 -7386
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 14058
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 669454 452414 705242
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 273454 452414 308898
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -1306 452414 20898
rect 451794 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 452414 -1306
rect 451794 -1626 452414 -1542
rect 451794 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 452414 -1626
rect 451794 -1894 452414 -1862
rect 455514 673174 456134 707162
rect 455514 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 456134 673174
rect 455514 672854 456134 672938
rect 455514 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 456134 672854
rect 455514 637174 456134 672618
rect 455514 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 456134 637174
rect 455514 636854 456134 636938
rect 455514 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 456134 636854
rect 455514 601174 456134 636618
rect 455514 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 456134 601174
rect 455514 600854 456134 600938
rect 455514 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 456134 600854
rect 455514 565174 456134 600618
rect 455514 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 456134 565174
rect 455514 564854 456134 564938
rect 455514 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 456134 564854
rect 455514 529174 456134 564618
rect 455514 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 456134 529174
rect 455514 528854 456134 528938
rect 455514 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 456134 528854
rect 455514 493174 456134 528618
rect 455514 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 456134 493174
rect 455514 492854 456134 492938
rect 455514 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 456134 492854
rect 455514 457174 456134 492618
rect 455514 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 456134 457174
rect 455514 456854 456134 456938
rect 455514 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 456134 456854
rect 455514 421174 456134 456618
rect 455514 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 456134 421174
rect 455514 420854 456134 420938
rect 455514 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 456134 420854
rect 455514 385174 456134 420618
rect 455514 384938 455546 385174
rect 455782 384938 455866 385174
rect 456102 384938 456134 385174
rect 455514 384854 456134 384938
rect 455514 384618 455546 384854
rect 455782 384618 455866 384854
rect 456102 384618 456134 384854
rect 455514 349174 456134 384618
rect 455514 348938 455546 349174
rect 455782 348938 455866 349174
rect 456102 348938 456134 349174
rect 455514 348854 456134 348938
rect 455514 348618 455546 348854
rect 455782 348618 455866 348854
rect 456102 348618 456134 348854
rect 455514 313174 456134 348618
rect 455514 312938 455546 313174
rect 455782 312938 455866 313174
rect 456102 312938 456134 313174
rect 455514 312854 456134 312938
rect 455514 312618 455546 312854
rect 455782 312618 455866 312854
rect 456102 312618 456134 312854
rect 455514 277174 456134 312618
rect 455514 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 456134 277174
rect 455514 276854 456134 276938
rect 455514 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 456134 276854
rect 455514 241174 456134 276618
rect 455514 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 456134 241174
rect 455514 240854 456134 240938
rect 455514 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 456134 240854
rect 455514 205174 456134 240618
rect 455514 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 456134 205174
rect 455514 204854 456134 204938
rect 455514 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 456134 204854
rect 455514 169174 456134 204618
rect 455514 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 456134 169174
rect 455514 168854 456134 168938
rect 455514 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 456134 168854
rect 455514 133174 456134 168618
rect 455514 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 456134 133174
rect 455514 132854 456134 132938
rect 455514 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 456134 132854
rect 455514 97174 456134 132618
rect 455514 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 456134 97174
rect 455514 96854 456134 96938
rect 455514 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 456134 96854
rect 455514 61174 456134 96618
rect 455514 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 456134 61174
rect 455514 60854 456134 60938
rect 455514 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 456134 60854
rect 455514 25174 456134 60618
rect 455514 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 456134 25174
rect 455514 24854 456134 24938
rect 455514 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 456134 24854
rect 455514 -3226 456134 24618
rect 455514 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 456134 -3226
rect 455514 -3546 456134 -3462
rect 455514 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 456134 -3546
rect 455514 -3814 456134 -3782
rect 459234 676894 459854 709082
rect 459234 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 459854 676894
rect 459234 676574 459854 676658
rect 459234 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 459854 676574
rect 459234 640894 459854 676338
rect 459234 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 459854 640894
rect 459234 640574 459854 640658
rect 459234 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 459854 640574
rect 459234 604894 459854 640338
rect 459234 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 459854 604894
rect 459234 604574 459854 604658
rect 459234 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 459854 604574
rect 459234 568894 459854 604338
rect 459234 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 459854 568894
rect 459234 568574 459854 568658
rect 459234 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 459854 568574
rect 459234 532894 459854 568338
rect 459234 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 459854 532894
rect 459234 532574 459854 532658
rect 459234 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 459854 532574
rect 459234 496894 459854 532338
rect 459234 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 459854 496894
rect 459234 496574 459854 496658
rect 459234 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 459854 496574
rect 459234 460894 459854 496338
rect 459234 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 459854 460894
rect 459234 460574 459854 460658
rect 459234 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 459854 460574
rect 459234 424894 459854 460338
rect 459234 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 459854 424894
rect 459234 424574 459854 424658
rect 459234 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 459854 424574
rect 459234 388894 459854 424338
rect 459234 388658 459266 388894
rect 459502 388658 459586 388894
rect 459822 388658 459854 388894
rect 459234 388574 459854 388658
rect 459234 388338 459266 388574
rect 459502 388338 459586 388574
rect 459822 388338 459854 388574
rect 459234 352894 459854 388338
rect 459234 352658 459266 352894
rect 459502 352658 459586 352894
rect 459822 352658 459854 352894
rect 459234 352574 459854 352658
rect 459234 352338 459266 352574
rect 459502 352338 459586 352574
rect 459822 352338 459854 352574
rect 459234 316894 459854 352338
rect 459234 316658 459266 316894
rect 459502 316658 459586 316894
rect 459822 316658 459854 316894
rect 459234 316574 459854 316658
rect 459234 316338 459266 316574
rect 459502 316338 459586 316574
rect 459822 316338 459854 316574
rect 459234 280894 459854 316338
rect 459234 280658 459266 280894
rect 459502 280658 459586 280894
rect 459822 280658 459854 280894
rect 459234 280574 459854 280658
rect 459234 280338 459266 280574
rect 459502 280338 459586 280574
rect 459822 280338 459854 280574
rect 459234 244894 459854 280338
rect 459234 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 459854 244894
rect 459234 244574 459854 244658
rect 459234 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 459854 244574
rect 459234 208894 459854 244338
rect 459234 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 459854 208894
rect 459234 208574 459854 208658
rect 459234 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 459854 208574
rect 459234 172894 459854 208338
rect 459234 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 459854 172894
rect 459234 172574 459854 172658
rect 459234 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 459854 172574
rect 459234 136894 459854 172338
rect 459234 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 459854 136894
rect 459234 136574 459854 136658
rect 459234 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 459854 136574
rect 459234 100894 459854 136338
rect 459234 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 459854 100894
rect 459234 100574 459854 100658
rect 459234 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 459854 100574
rect 459234 64894 459854 100338
rect 459234 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 459854 64894
rect 459234 64574 459854 64658
rect 459234 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 459854 64574
rect 459234 28894 459854 64338
rect 459234 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 459854 28894
rect 459234 28574 459854 28658
rect 459234 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 459854 28574
rect 459234 -5146 459854 28338
rect 459234 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 459854 -5146
rect 459234 -5466 459854 -5382
rect 459234 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 459854 -5466
rect 459234 -5734 459854 -5702
rect 462954 680614 463574 711002
rect 480954 710598 481574 711590
rect 480954 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 481574 710598
rect 480954 710278 481574 710362
rect 480954 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 481574 710278
rect 477234 708678 477854 709670
rect 477234 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 477854 708678
rect 477234 708358 477854 708442
rect 477234 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 477854 708358
rect 473514 706758 474134 707750
rect 473514 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 474134 706758
rect 473514 706438 474134 706522
rect 473514 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 474134 706438
rect 462954 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 463574 680614
rect 462954 680294 463574 680378
rect 462954 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 463574 680294
rect 462954 644614 463574 680058
rect 462954 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 463574 644614
rect 462954 644294 463574 644378
rect 462954 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 463574 644294
rect 462954 608614 463574 644058
rect 462954 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 463574 608614
rect 462954 608294 463574 608378
rect 462954 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 463574 608294
rect 462954 572614 463574 608058
rect 462954 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 463574 572614
rect 462954 572294 463574 572378
rect 462954 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 463574 572294
rect 462954 536614 463574 572058
rect 462954 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 463574 536614
rect 462954 536294 463574 536378
rect 462954 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 463574 536294
rect 462954 500614 463574 536058
rect 462954 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 463574 500614
rect 462954 500294 463574 500378
rect 462954 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 463574 500294
rect 462954 464614 463574 500058
rect 462954 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 463574 464614
rect 462954 464294 463574 464378
rect 462954 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 463574 464294
rect 462954 428614 463574 464058
rect 462954 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 463574 428614
rect 462954 428294 463574 428378
rect 462954 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 463574 428294
rect 462954 392614 463574 428058
rect 462954 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 463574 392614
rect 462954 392294 463574 392378
rect 462954 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 463574 392294
rect 462954 356614 463574 392058
rect 462954 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 463574 356614
rect 462954 356294 463574 356378
rect 462954 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 463574 356294
rect 462954 320614 463574 356058
rect 462954 320378 462986 320614
rect 463222 320378 463306 320614
rect 463542 320378 463574 320614
rect 462954 320294 463574 320378
rect 462954 320058 462986 320294
rect 463222 320058 463306 320294
rect 463542 320058 463574 320294
rect 462954 284614 463574 320058
rect 462954 284378 462986 284614
rect 463222 284378 463306 284614
rect 463542 284378 463574 284614
rect 462954 284294 463574 284378
rect 462954 284058 462986 284294
rect 463222 284058 463306 284294
rect 463542 284058 463574 284294
rect 462954 248614 463574 284058
rect 462954 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 463574 248614
rect 462954 248294 463574 248378
rect 462954 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 463574 248294
rect 462954 212614 463574 248058
rect 462954 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 463574 212614
rect 462954 212294 463574 212378
rect 462954 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 463574 212294
rect 462954 176614 463574 212058
rect 462954 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 463574 176614
rect 462954 176294 463574 176378
rect 462954 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 463574 176294
rect 462954 140614 463574 176058
rect 462954 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 463574 140614
rect 462954 140294 463574 140378
rect 462954 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 463574 140294
rect 462954 104614 463574 140058
rect 462954 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 463574 104614
rect 462954 104294 463574 104378
rect 462954 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 463574 104294
rect 462954 68614 463574 104058
rect 462954 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 463574 68614
rect 462954 68294 463574 68378
rect 462954 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 463574 68294
rect 462954 32614 463574 68058
rect 462954 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 463574 32614
rect 462954 32294 463574 32378
rect 462954 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 463574 32294
rect 444954 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 445574 -6106
rect 444954 -6426 445574 -6342
rect 444954 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 445574 -6426
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 32058
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 473514 691174 474134 706202
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 655174 474134 690618
rect 473514 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 474134 655174
rect 473514 654854 474134 654938
rect 473514 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 474134 654854
rect 473514 619174 474134 654618
rect 473514 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 474134 619174
rect 473514 618854 474134 618938
rect 473514 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 474134 618854
rect 473514 583174 474134 618618
rect 473514 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 474134 583174
rect 473514 582854 474134 582938
rect 473514 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 474134 582854
rect 473514 547174 474134 582618
rect 473514 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 474134 547174
rect 473514 546854 474134 546938
rect 473514 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 474134 546854
rect 473514 511174 474134 546618
rect 473514 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 474134 511174
rect 473514 510854 474134 510938
rect 473514 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 474134 510854
rect 473514 475174 474134 510618
rect 473514 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 474134 475174
rect 473514 474854 474134 474938
rect 473514 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 474134 474854
rect 473514 439174 474134 474618
rect 473514 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 474134 439174
rect 473514 438854 474134 438938
rect 473514 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 474134 438854
rect 473514 403174 474134 438618
rect 473514 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 474134 403174
rect 473514 402854 474134 402938
rect 473514 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 474134 402854
rect 473514 367174 474134 402618
rect 473514 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 474134 367174
rect 473514 366854 474134 366938
rect 473514 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 474134 366854
rect 473514 331174 474134 366618
rect 473514 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 474134 331174
rect 473514 330854 474134 330938
rect 473514 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 474134 330854
rect 473514 295174 474134 330618
rect 473514 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 474134 295174
rect 473514 294854 474134 294938
rect 473514 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 474134 294854
rect 473514 259174 474134 294618
rect 473514 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 474134 259174
rect 473514 258854 474134 258938
rect 473514 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 474134 258854
rect 473514 223174 474134 258618
rect 473514 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 474134 223174
rect 473514 222854 474134 222938
rect 473514 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 474134 222854
rect 473514 187174 474134 222618
rect 473514 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 474134 187174
rect 473514 186854 474134 186938
rect 473514 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 474134 186854
rect 473514 151174 474134 186618
rect 473514 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 474134 151174
rect 473514 150854 474134 150938
rect 473514 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 474134 150854
rect 473514 115174 474134 150618
rect 473514 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 474134 115174
rect 473514 114854 474134 114938
rect 473514 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 474134 114854
rect 473514 79174 474134 114618
rect 473514 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 474134 79174
rect 473514 78854 474134 78938
rect 473514 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 474134 78854
rect 473514 43174 474134 78618
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 473514 7174 474134 42618
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -2266 474134 6618
rect 473514 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 474134 -2266
rect 473514 -2586 474134 -2502
rect 473514 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 474134 -2586
rect 473514 -3814 474134 -2822
rect 477234 694894 477854 708122
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 658894 477854 694338
rect 477234 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 477854 658894
rect 477234 658574 477854 658658
rect 477234 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 477854 658574
rect 477234 622894 477854 658338
rect 477234 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 477854 622894
rect 477234 622574 477854 622658
rect 477234 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 477854 622574
rect 477234 586894 477854 622338
rect 477234 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 477854 586894
rect 477234 586574 477854 586658
rect 477234 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 477854 586574
rect 477234 550894 477854 586338
rect 477234 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 477854 550894
rect 477234 550574 477854 550658
rect 477234 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 477854 550574
rect 477234 514894 477854 550338
rect 477234 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 477854 514894
rect 477234 514574 477854 514658
rect 477234 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 477854 514574
rect 477234 478894 477854 514338
rect 477234 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 477854 478894
rect 477234 478574 477854 478658
rect 477234 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 477854 478574
rect 477234 442894 477854 478338
rect 477234 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 477854 442894
rect 477234 442574 477854 442658
rect 477234 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 477854 442574
rect 477234 406894 477854 442338
rect 477234 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 477854 406894
rect 477234 406574 477854 406658
rect 477234 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 477854 406574
rect 477234 370894 477854 406338
rect 477234 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 477854 370894
rect 477234 370574 477854 370658
rect 477234 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 477854 370574
rect 477234 334894 477854 370338
rect 477234 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 477854 334894
rect 477234 334574 477854 334658
rect 477234 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 477854 334574
rect 477234 298894 477854 334338
rect 477234 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 477854 298894
rect 477234 298574 477854 298658
rect 477234 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 477854 298574
rect 477234 262894 477854 298338
rect 477234 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 477854 262894
rect 477234 262574 477854 262658
rect 477234 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 477854 262574
rect 477234 226894 477854 262338
rect 477234 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 477854 226894
rect 477234 226574 477854 226658
rect 477234 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 477854 226574
rect 477234 190894 477854 226338
rect 477234 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 477854 190894
rect 477234 190574 477854 190658
rect 477234 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 477854 190574
rect 477234 154894 477854 190338
rect 477234 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 477854 154894
rect 477234 154574 477854 154658
rect 477234 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 477854 154574
rect 477234 118894 477854 154338
rect 477234 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 477854 118894
rect 477234 118574 477854 118658
rect 477234 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 477854 118574
rect 477234 82894 477854 118338
rect 477234 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 477854 82894
rect 477234 82574 477854 82658
rect 477234 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 477854 82574
rect 477234 46894 477854 82338
rect 477234 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 477854 46894
rect 477234 46574 477854 46658
rect 477234 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 477854 46574
rect 477234 10894 477854 46338
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -4186 477854 10338
rect 477234 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 477854 -4186
rect 477234 -4506 477854 -4422
rect 477234 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 477854 -4506
rect 477234 -5734 477854 -4742
rect 480954 698614 481574 710042
rect 498954 711558 499574 711590
rect 498954 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 499574 711558
rect 498954 711238 499574 711322
rect 498954 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 499574 711238
rect 495234 709638 495854 709670
rect 495234 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 495854 709638
rect 495234 709318 495854 709402
rect 495234 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 495854 709318
rect 491514 707718 492134 707750
rect 491514 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 492134 707718
rect 491514 707398 492134 707482
rect 491514 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 492134 707398
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 662614 481574 698058
rect 480954 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 481574 662614
rect 480954 662294 481574 662378
rect 480954 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 481574 662294
rect 480954 626614 481574 662058
rect 480954 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 481574 626614
rect 480954 626294 481574 626378
rect 480954 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 481574 626294
rect 480954 590614 481574 626058
rect 480954 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 481574 590614
rect 480954 590294 481574 590378
rect 480954 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 481574 590294
rect 480954 554614 481574 590058
rect 480954 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 481574 554614
rect 480954 554294 481574 554378
rect 480954 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 481574 554294
rect 480954 518614 481574 554058
rect 480954 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 481574 518614
rect 480954 518294 481574 518378
rect 480954 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 481574 518294
rect 480954 482614 481574 518058
rect 480954 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 481574 482614
rect 480954 482294 481574 482378
rect 480954 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 481574 482294
rect 480954 446614 481574 482058
rect 480954 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 481574 446614
rect 480954 446294 481574 446378
rect 480954 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 481574 446294
rect 480954 410614 481574 446058
rect 480954 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 481574 410614
rect 480954 410294 481574 410378
rect 480954 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 481574 410294
rect 480954 374614 481574 410058
rect 480954 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 481574 374614
rect 480954 374294 481574 374378
rect 480954 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 481574 374294
rect 480954 338614 481574 374058
rect 480954 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 481574 338614
rect 480954 338294 481574 338378
rect 480954 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 481574 338294
rect 480954 302614 481574 338058
rect 480954 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 481574 302614
rect 480954 302294 481574 302378
rect 480954 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 481574 302294
rect 480954 266614 481574 302058
rect 480954 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 481574 266614
rect 480954 266294 481574 266378
rect 480954 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 481574 266294
rect 480954 230614 481574 266058
rect 480954 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 481574 230614
rect 480954 230294 481574 230378
rect 480954 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 481574 230294
rect 480954 194614 481574 230058
rect 480954 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 481574 194614
rect 480954 194294 481574 194378
rect 480954 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 481574 194294
rect 480954 158614 481574 194058
rect 480954 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 481574 158614
rect 480954 158294 481574 158378
rect 480954 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 481574 158294
rect 480954 122614 481574 158058
rect 480954 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 481574 122614
rect 480954 122294 481574 122378
rect 480954 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 481574 122294
rect 480954 86614 481574 122058
rect 480954 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 481574 86614
rect 480954 86294 481574 86378
rect 480954 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 481574 86294
rect 480954 50614 481574 86058
rect 480954 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 481574 50614
rect 480954 50294 481574 50378
rect 480954 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 481574 50294
rect 480954 14614 481574 50058
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 462954 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 463574 -7066
rect 462954 -7386 463574 -7302
rect 462954 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 463574 -7386
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 14058
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 487794 669454 488414 705242
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -1306 488414 20898
rect 487794 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 488414 -1306
rect 487794 -1626 488414 -1542
rect 487794 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 488414 -1626
rect 487794 -1894 488414 -1862
rect 491514 673174 492134 707162
rect 491514 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 492134 673174
rect 491514 672854 492134 672938
rect 491514 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 492134 672854
rect 491514 637174 492134 672618
rect 491514 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 492134 637174
rect 491514 636854 492134 636938
rect 491514 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 492134 636854
rect 491514 601174 492134 636618
rect 491514 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 492134 601174
rect 491514 600854 492134 600938
rect 491514 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 492134 600854
rect 491514 565174 492134 600618
rect 491514 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 492134 565174
rect 491514 564854 492134 564938
rect 491514 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 492134 564854
rect 491514 529174 492134 564618
rect 491514 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 492134 529174
rect 491514 528854 492134 528938
rect 491514 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 492134 528854
rect 491514 493174 492134 528618
rect 491514 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 492134 493174
rect 491514 492854 492134 492938
rect 491514 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 492134 492854
rect 491514 457174 492134 492618
rect 491514 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 492134 457174
rect 491514 456854 492134 456938
rect 491514 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 492134 456854
rect 491514 421174 492134 456618
rect 491514 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 492134 421174
rect 491514 420854 492134 420938
rect 491514 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 492134 420854
rect 491514 385174 492134 420618
rect 491514 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 492134 385174
rect 491514 384854 492134 384938
rect 491514 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 492134 384854
rect 491514 349174 492134 384618
rect 491514 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 492134 349174
rect 491514 348854 492134 348938
rect 491514 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 492134 348854
rect 491514 313174 492134 348618
rect 491514 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 492134 313174
rect 491514 312854 492134 312938
rect 491514 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 492134 312854
rect 491514 277174 492134 312618
rect 491514 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 492134 277174
rect 491514 276854 492134 276938
rect 491514 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 492134 276854
rect 491514 241174 492134 276618
rect 491514 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 492134 241174
rect 491514 240854 492134 240938
rect 491514 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 492134 240854
rect 491514 205174 492134 240618
rect 491514 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 492134 205174
rect 491514 204854 492134 204938
rect 491514 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 492134 204854
rect 491514 169174 492134 204618
rect 491514 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 492134 169174
rect 491514 168854 492134 168938
rect 491514 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 492134 168854
rect 491514 133174 492134 168618
rect 491514 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 492134 133174
rect 491514 132854 492134 132938
rect 491514 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 492134 132854
rect 491514 97174 492134 132618
rect 491514 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 492134 97174
rect 491514 96854 492134 96938
rect 491514 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 492134 96854
rect 491514 61174 492134 96618
rect 491514 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 492134 61174
rect 491514 60854 492134 60938
rect 491514 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 492134 60854
rect 491514 25174 492134 60618
rect 491514 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 492134 25174
rect 491514 24854 492134 24938
rect 491514 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 492134 24854
rect 491514 -3226 492134 24618
rect 491514 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 492134 -3226
rect 491514 -3546 492134 -3462
rect 491514 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 492134 -3546
rect 491514 -3814 492134 -3782
rect 495234 676894 495854 709082
rect 495234 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 495854 676894
rect 495234 676574 495854 676658
rect 495234 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 495854 676574
rect 495234 640894 495854 676338
rect 495234 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 495854 640894
rect 495234 640574 495854 640658
rect 495234 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 495854 640574
rect 495234 604894 495854 640338
rect 495234 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 495854 604894
rect 495234 604574 495854 604658
rect 495234 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 495854 604574
rect 495234 568894 495854 604338
rect 495234 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 495854 568894
rect 495234 568574 495854 568658
rect 495234 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 495854 568574
rect 495234 532894 495854 568338
rect 495234 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 495854 532894
rect 495234 532574 495854 532658
rect 495234 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 495854 532574
rect 495234 496894 495854 532338
rect 495234 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 495854 496894
rect 495234 496574 495854 496658
rect 495234 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 495854 496574
rect 495234 460894 495854 496338
rect 495234 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 495854 460894
rect 495234 460574 495854 460658
rect 495234 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 495854 460574
rect 495234 424894 495854 460338
rect 495234 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 495854 424894
rect 495234 424574 495854 424658
rect 495234 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 495854 424574
rect 495234 388894 495854 424338
rect 495234 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 495854 388894
rect 495234 388574 495854 388658
rect 495234 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 495854 388574
rect 495234 352894 495854 388338
rect 495234 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 495854 352894
rect 495234 352574 495854 352658
rect 495234 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 495854 352574
rect 495234 316894 495854 352338
rect 495234 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 495854 316894
rect 495234 316574 495854 316658
rect 495234 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 495854 316574
rect 495234 280894 495854 316338
rect 495234 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 495854 280894
rect 495234 280574 495854 280658
rect 495234 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 495854 280574
rect 495234 244894 495854 280338
rect 495234 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 495854 244894
rect 495234 244574 495854 244658
rect 495234 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 495854 244574
rect 495234 208894 495854 244338
rect 495234 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 495854 208894
rect 495234 208574 495854 208658
rect 495234 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 495854 208574
rect 495234 172894 495854 208338
rect 495234 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 495854 172894
rect 495234 172574 495854 172658
rect 495234 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 495854 172574
rect 495234 136894 495854 172338
rect 495234 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 495854 136894
rect 495234 136574 495854 136658
rect 495234 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 495854 136574
rect 495234 100894 495854 136338
rect 495234 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 495854 100894
rect 495234 100574 495854 100658
rect 495234 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 495854 100574
rect 495234 64894 495854 100338
rect 495234 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 495854 64894
rect 495234 64574 495854 64658
rect 495234 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 495854 64574
rect 495234 28894 495854 64338
rect 495234 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 495854 28894
rect 495234 28574 495854 28658
rect 495234 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 495854 28574
rect 495234 -5146 495854 28338
rect 495234 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 495854 -5146
rect 495234 -5466 495854 -5382
rect 495234 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 495854 -5466
rect 495234 -5734 495854 -5702
rect 498954 680614 499574 711002
rect 516954 710598 517574 711590
rect 516954 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 517574 710598
rect 516954 710278 517574 710362
rect 516954 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 517574 710278
rect 513234 708678 513854 709670
rect 513234 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 513854 708678
rect 513234 708358 513854 708442
rect 513234 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 513854 708358
rect 509514 706758 510134 707750
rect 509514 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 510134 706758
rect 509514 706438 510134 706522
rect 509514 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 510134 706438
rect 498954 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 499574 680614
rect 498954 680294 499574 680378
rect 498954 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 499574 680294
rect 498954 644614 499574 680058
rect 498954 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 499574 644614
rect 498954 644294 499574 644378
rect 498954 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 499574 644294
rect 498954 608614 499574 644058
rect 498954 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 499574 608614
rect 498954 608294 499574 608378
rect 498954 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 499574 608294
rect 498954 572614 499574 608058
rect 498954 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 499574 572614
rect 498954 572294 499574 572378
rect 498954 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 499574 572294
rect 498954 536614 499574 572058
rect 498954 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 499574 536614
rect 498954 536294 499574 536378
rect 498954 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 499574 536294
rect 498954 500614 499574 536058
rect 498954 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 499574 500614
rect 498954 500294 499574 500378
rect 498954 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 499574 500294
rect 498954 464614 499574 500058
rect 498954 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 499574 464614
rect 498954 464294 499574 464378
rect 498954 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 499574 464294
rect 498954 428614 499574 464058
rect 498954 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 499574 428614
rect 498954 428294 499574 428378
rect 498954 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 499574 428294
rect 498954 392614 499574 428058
rect 498954 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 499574 392614
rect 498954 392294 499574 392378
rect 498954 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 499574 392294
rect 498954 356614 499574 392058
rect 498954 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 499574 356614
rect 498954 356294 499574 356378
rect 498954 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 499574 356294
rect 498954 320614 499574 356058
rect 498954 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 499574 320614
rect 498954 320294 499574 320378
rect 498954 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 499574 320294
rect 498954 284614 499574 320058
rect 498954 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 499574 284614
rect 498954 284294 499574 284378
rect 498954 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 499574 284294
rect 498954 248614 499574 284058
rect 498954 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 499574 248614
rect 498954 248294 499574 248378
rect 498954 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 499574 248294
rect 498954 212614 499574 248058
rect 498954 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 499574 212614
rect 498954 212294 499574 212378
rect 498954 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 499574 212294
rect 498954 176614 499574 212058
rect 498954 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 499574 176614
rect 498954 176294 499574 176378
rect 498954 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 499574 176294
rect 498954 140614 499574 176058
rect 498954 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 499574 140614
rect 498954 140294 499574 140378
rect 498954 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 499574 140294
rect 498954 104614 499574 140058
rect 498954 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 499574 104614
rect 498954 104294 499574 104378
rect 498954 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 499574 104294
rect 498954 68614 499574 104058
rect 498954 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 499574 68614
rect 498954 68294 499574 68378
rect 498954 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 499574 68294
rect 498954 32614 499574 68058
rect 498954 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 499574 32614
rect 498954 32294 499574 32378
rect 498954 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 499574 32294
rect 480954 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 481574 -6106
rect 480954 -6426 481574 -6342
rect 480954 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 481574 -6426
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 32058
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 509514 691174 510134 706202
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 655174 510134 690618
rect 509514 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 510134 655174
rect 509514 654854 510134 654938
rect 509514 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 510134 654854
rect 509514 619174 510134 654618
rect 509514 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 510134 619174
rect 509514 618854 510134 618938
rect 509514 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 510134 618854
rect 509514 583174 510134 618618
rect 509514 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 510134 583174
rect 509514 582854 510134 582938
rect 509514 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 510134 582854
rect 509514 547174 510134 582618
rect 509514 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 510134 547174
rect 509514 546854 510134 546938
rect 509514 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 510134 546854
rect 509514 511174 510134 546618
rect 509514 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 510134 511174
rect 509514 510854 510134 510938
rect 509514 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 510134 510854
rect 509514 475174 510134 510618
rect 509514 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 510134 475174
rect 509514 474854 510134 474938
rect 509514 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 510134 474854
rect 509514 439174 510134 474618
rect 509514 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 510134 439174
rect 509514 438854 510134 438938
rect 509514 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 510134 438854
rect 509514 403174 510134 438618
rect 509514 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 510134 403174
rect 509514 402854 510134 402938
rect 509514 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 510134 402854
rect 509514 367174 510134 402618
rect 509514 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 510134 367174
rect 509514 366854 510134 366938
rect 509514 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 510134 366854
rect 509514 331174 510134 366618
rect 509514 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 510134 331174
rect 509514 330854 510134 330938
rect 509514 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 510134 330854
rect 509514 295174 510134 330618
rect 509514 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 510134 295174
rect 509514 294854 510134 294938
rect 509514 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 510134 294854
rect 509514 259174 510134 294618
rect 509514 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 510134 259174
rect 509514 258854 510134 258938
rect 509514 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 510134 258854
rect 509514 223174 510134 258618
rect 509514 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 510134 223174
rect 509514 222854 510134 222938
rect 509514 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 510134 222854
rect 509514 187174 510134 222618
rect 509514 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 510134 187174
rect 509514 186854 510134 186938
rect 509514 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 510134 186854
rect 509514 151174 510134 186618
rect 509514 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 510134 151174
rect 509514 150854 510134 150938
rect 509514 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 510134 150854
rect 509514 115174 510134 150618
rect 509514 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 510134 115174
rect 509514 114854 510134 114938
rect 509514 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 510134 114854
rect 509514 79174 510134 114618
rect 509514 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 510134 79174
rect 509514 78854 510134 78938
rect 509514 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 510134 78854
rect 509514 43174 510134 78618
rect 509514 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 510134 43174
rect 509514 42854 510134 42938
rect 509514 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 510134 42854
rect 509514 7174 510134 42618
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -2266 510134 6618
rect 509514 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 510134 -2266
rect 509514 -2586 510134 -2502
rect 509514 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 510134 -2586
rect 509514 -3814 510134 -2822
rect 513234 694894 513854 708122
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 658894 513854 694338
rect 513234 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 513854 658894
rect 513234 658574 513854 658658
rect 513234 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 513854 658574
rect 513234 622894 513854 658338
rect 513234 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 513854 622894
rect 513234 622574 513854 622658
rect 513234 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 513854 622574
rect 513234 586894 513854 622338
rect 513234 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 513854 586894
rect 513234 586574 513854 586658
rect 513234 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 513854 586574
rect 513234 550894 513854 586338
rect 513234 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 513854 550894
rect 513234 550574 513854 550658
rect 513234 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 513854 550574
rect 513234 514894 513854 550338
rect 513234 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 513854 514894
rect 513234 514574 513854 514658
rect 513234 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 513854 514574
rect 513234 478894 513854 514338
rect 513234 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 513854 478894
rect 513234 478574 513854 478658
rect 513234 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 513854 478574
rect 513234 442894 513854 478338
rect 513234 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 513854 442894
rect 513234 442574 513854 442658
rect 513234 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 513854 442574
rect 513234 406894 513854 442338
rect 513234 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 513854 406894
rect 513234 406574 513854 406658
rect 513234 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 513854 406574
rect 513234 370894 513854 406338
rect 513234 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 513854 370894
rect 513234 370574 513854 370658
rect 513234 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 513854 370574
rect 513234 334894 513854 370338
rect 513234 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 513854 334894
rect 513234 334574 513854 334658
rect 513234 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 513854 334574
rect 513234 298894 513854 334338
rect 513234 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 513854 298894
rect 513234 298574 513854 298658
rect 513234 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 513854 298574
rect 513234 262894 513854 298338
rect 513234 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 513854 262894
rect 513234 262574 513854 262658
rect 513234 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 513854 262574
rect 513234 226894 513854 262338
rect 513234 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 513854 226894
rect 513234 226574 513854 226658
rect 513234 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 513854 226574
rect 513234 190894 513854 226338
rect 513234 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 513854 190894
rect 513234 190574 513854 190658
rect 513234 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 513854 190574
rect 513234 154894 513854 190338
rect 513234 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 513854 154894
rect 513234 154574 513854 154658
rect 513234 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 513854 154574
rect 513234 118894 513854 154338
rect 513234 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 513854 118894
rect 513234 118574 513854 118658
rect 513234 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 513854 118574
rect 513234 82894 513854 118338
rect 513234 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 513854 82894
rect 513234 82574 513854 82658
rect 513234 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 513854 82574
rect 513234 46894 513854 82338
rect 513234 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 513854 46894
rect 513234 46574 513854 46658
rect 513234 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 513854 46574
rect 513234 10894 513854 46338
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -4186 513854 10338
rect 513234 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 513854 -4186
rect 513234 -4506 513854 -4422
rect 513234 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 513854 -4506
rect 513234 -5734 513854 -4742
rect 516954 698614 517574 710042
rect 534954 711558 535574 711590
rect 534954 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 535574 711558
rect 534954 711238 535574 711322
rect 534954 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 535574 711238
rect 531234 709638 531854 709670
rect 531234 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 531854 709638
rect 531234 709318 531854 709402
rect 531234 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 531854 709318
rect 527514 707718 528134 707750
rect 527514 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 528134 707718
rect 527514 707398 528134 707482
rect 527514 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 528134 707398
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 662614 517574 698058
rect 516954 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 517574 662614
rect 516954 662294 517574 662378
rect 516954 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 517574 662294
rect 516954 626614 517574 662058
rect 516954 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 517574 626614
rect 516954 626294 517574 626378
rect 516954 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 517574 626294
rect 516954 590614 517574 626058
rect 516954 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 517574 590614
rect 516954 590294 517574 590378
rect 516954 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 517574 590294
rect 516954 554614 517574 590058
rect 516954 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 517574 554614
rect 516954 554294 517574 554378
rect 516954 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 517574 554294
rect 516954 518614 517574 554058
rect 516954 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 517574 518614
rect 516954 518294 517574 518378
rect 516954 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 517574 518294
rect 516954 482614 517574 518058
rect 516954 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 517574 482614
rect 516954 482294 517574 482378
rect 516954 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 517574 482294
rect 516954 446614 517574 482058
rect 516954 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 517574 446614
rect 516954 446294 517574 446378
rect 516954 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 517574 446294
rect 516954 410614 517574 446058
rect 516954 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 517574 410614
rect 516954 410294 517574 410378
rect 516954 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 517574 410294
rect 516954 374614 517574 410058
rect 516954 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 517574 374614
rect 516954 374294 517574 374378
rect 516954 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 517574 374294
rect 516954 338614 517574 374058
rect 516954 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 517574 338614
rect 516954 338294 517574 338378
rect 516954 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 517574 338294
rect 516954 302614 517574 338058
rect 516954 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 517574 302614
rect 516954 302294 517574 302378
rect 516954 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 517574 302294
rect 516954 266614 517574 302058
rect 516954 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 517574 266614
rect 516954 266294 517574 266378
rect 516954 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 517574 266294
rect 516954 230614 517574 266058
rect 516954 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 517574 230614
rect 516954 230294 517574 230378
rect 516954 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 517574 230294
rect 516954 194614 517574 230058
rect 516954 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 517574 194614
rect 516954 194294 517574 194378
rect 516954 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 517574 194294
rect 516954 158614 517574 194058
rect 516954 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 517574 158614
rect 516954 158294 517574 158378
rect 516954 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 517574 158294
rect 516954 122614 517574 158058
rect 516954 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 517574 122614
rect 516954 122294 517574 122378
rect 516954 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 517574 122294
rect 516954 86614 517574 122058
rect 516954 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 517574 86614
rect 516954 86294 517574 86378
rect 516954 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 517574 86294
rect 516954 50614 517574 86058
rect 516954 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 517574 50614
rect 516954 50294 517574 50378
rect 516954 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 517574 50294
rect 516954 14614 517574 50058
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 498954 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 499574 -7066
rect 498954 -7386 499574 -7302
rect 498954 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 499574 -7386
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 14058
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 669454 524414 705242
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -1306 524414 20898
rect 523794 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 524414 -1306
rect 523794 -1626 524414 -1542
rect 523794 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 524414 -1626
rect 523794 -1894 524414 -1862
rect 527514 673174 528134 707162
rect 527514 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 528134 673174
rect 527514 672854 528134 672938
rect 527514 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 528134 672854
rect 527514 637174 528134 672618
rect 527514 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 528134 637174
rect 527514 636854 528134 636938
rect 527514 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 528134 636854
rect 527514 601174 528134 636618
rect 527514 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 528134 601174
rect 527514 600854 528134 600938
rect 527514 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 528134 600854
rect 527514 565174 528134 600618
rect 527514 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 528134 565174
rect 527514 564854 528134 564938
rect 527514 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 528134 564854
rect 527514 529174 528134 564618
rect 527514 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 528134 529174
rect 527514 528854 528134 528938
rect 527514 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 528134 528854
rect 527514 493174 528134 528618
rect 527514 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 528134 493174
rect 527514 492854 528134 492938
rect 527514 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 528134 492854
rect 527514 457174 528134 492618
rect 527514 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 528134 457174
rect 527514 456854 528134 456938
rect 527514 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 528134 456854
rect 527514 421174 528134 456618
rect 527514 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 528134 421174
rect 527514 420854 528134 420938
rect 527514 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 528134 420854
rect 527514 385174 528134 420618
rect 527514 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 528134 385174
rect 527514 384854 528134 384938
rect 527514 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 528134 384854
rect 527514 349174 528134 384618
rect 527514 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 528134 349174
rect 527514 348854 528134 348938
rect 527514 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 528134 348854
rect 527514 313174 528134 348618
rect 527514 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 528134 313174
rect 527514 312854 528134 312938
rect 527514 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 528134 312854
rect 527514 277174 528134 312618
rect 527514 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 528134 277174
rect 527514 276854 528134 276938
rect 527514 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 528134 276854
rect 527514 241174 528134 276618
rect 527514 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 528134 241174
rect 527514 240854 528134 240938
rect 527514 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 528134 240854
rect 527514 205174 528134 240618
rect 527514 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 528134 205174
rect 527514 204854 528134 204938
rect 527514 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 528134 204854
rect 527514 169174 528134 204618
rect 527514 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 528134 169174
rect 527514 168854 528134 168938
rect 527514 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 528134 168854
rect 527514 133174 528134 168618
rect 527514 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 528134 133174
rect 527514 132854 528134 132938
rect 527514 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 528134 132854
rect 527514 97174 528134 132618
rect 527514 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 528134 97174
rect 527514 96854 528134 96938
rect 527514 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 528134 96854
rect 527514 61174 528134 96618
rect 527514 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 528134 61174
rect 527514 60854 528134 60938
rect 527514 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 528134 60854
rect 527514 25174 528134 60618
rect 527514 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 528134 25174
rect 527514 24854 528134 24938
rect 527514 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 528134 24854
rect 527514 -3226 528134 24618
rect 527514 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 528134 -3226
rect 527514 -3546 528134 -3462
rect 527514 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 528134 -3546
rect 527514 -3814 528134 -3782
rect 531234 676894 531854 709082
rect 531234 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 531854 676894
rect 531234 676574 531854 676658
rect 531234 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 531854 676574
rect 531234 640894 531854 676338
rect 531234 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 531854 640894
rect 531234 640574 531854 640658
rect 531234 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 531854 640574
rect 531234 604894 531854 640338
rect 531234 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 531854 604894
rect 531234 604574 531854 604658
rect 531234 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 531854 604574
rect 531234 568894 531854 604338
rect 531234 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 531854 568894
rect 531234 568574 531854 568658
rect 531234 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 531854 568574
rect 531234 532894 531854 568338
rect 531234 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 531854 532894
rect 531234 532574 531854 532658
rect 531234 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 531854 532574
rect 531234 496894 531854 532338
rect 531234 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 531854 496894
rect 531234 496574 531854 496658
rect 531234 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 531854 496574
rect 531234 460894 531854 496338
rect 531234 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 531854 460894
rect 531234 460574 531854 460658
rect 531234 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 531854 460574
rect 531234 424894 531854 460338
rect 531234 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 531854 424894
rect 531234 424574 531854 424658
rect 531234 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 531854 424574
rect 531234 388894 531854 424338
rect 531234 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 531854 388894
rect 531234 388574 531854 388658
rect 531234 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 531854 388574
rect 531234 352894 531854 388338
rect 531234 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 531854 352894
rect 531234 352574 531854 352658
rect 531234 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 531854 352574
rect 531234 316894 531854 352338
rect 531234 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 531854 316894
rect 531234 316574 531854 316658
rect 531234 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 531854 316574
rect 531234 280894 531854 316338
rect 531234 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 531854 280894
rect 531234 280574 531854 280658
rect 531234 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 531854 280574
rect 531234 244894 531854 280338
rect 531234 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 531854 244894
rect 531234 244574 531854 244658
rect 531234 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 531854 244574
rect 531234 208894 531854 244338
rect 531234 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 531854 208894
rect 531234 208574 531854 208658
rect 531234 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 531854 208574
rect 531234 172894 531854 208338
rect 531234 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 531854 172894
rect 531234 172574 531854 172658
rect 531234 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 531854 172574
rect 531234 136894 531854 172338
rect 531234 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 531854 136894
rect 531234 136574 531854 136658
rect 531234 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 531854 136574
rect 531234 100894 531854 136338
rect 531234 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 531854 100894
rect 531234 100574 531854 100658
rect 531234 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 531854 100574
rect 531234 64894 531854 100338
rect 531234 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 531854 64894
rect 531234 64574 531854 64658
rect 531234 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 531854 64574
rect 531234 28894 531854 64338
rect 531234 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 531854 28894
rect 531234 28574 531854 28658
rect 531234 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 531854 28574
rect 531234 -5146 531854 28338
rect 531234 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 531854 -5146
rect 531234 -5466 531854 -5382
rect 531234 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 531854 -5466
rect 531234 -5734 531854 -5702
rect 534954 680614 535574 711002
rect 552954 710598 553574 711590
rect 552954 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 553574 710598
rect 552954 710278 553574 710362
rect 552954 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 553574 710278
rect 549234 708678 549854 709670
rect 549234 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 549854 708678
rect 549234 708358 549854 708442
rect 549234 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 549854 708358
rect 545514 706758 546134 707750
rect 545514 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 546134 706758
rect 545514 706438 546134 706522
rect 545514 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 546134 706438
rect 534954 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 535574 680614
rect 534954 680294 535574 680378
rect 534954 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 535574 680294
rect 534954 644614 535574 680058
rect 534954 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 535574 644614
rect 534954 644294 535574 644378
rect 534954 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 535574 644294
rect 534954 608614 535574 644058
rect 534954 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 535574 608614
rect 534954 608294 535574 608378
rect 534954 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 535574 608294
rect 534954 572614 535574 608058
rect 534954 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 535574 572614
rect 534954 572294 535574 572378
rect 534954 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 535574 572294
rect 534954 536614 535574 572058
rect 534954 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 535574 536614
rect 534954 536294 535574 536378
rect 534954 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 535574 536294
rect 534954 500614 535574 536058
rect 534954 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 535574 500614
rect 534954 500294 535574 500378
rect 534954 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 535574 500294
rect 534954 464614 535574 500058
rect 534954 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 535574 464614
rect 534954 464294 535574 464378
rect 534954 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 535574 464294
rect 534954 428614 535574 464058
rect 534954 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 535574 428614
rect 534954 428294 535574 428378
rect 534954 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 535574 428294
rect 534954 392614 535574 428058
rect 534954 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 535574 392614
rect 534954 392294 535574 392378
rect 534954 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 535574 392294
rect 534954 356614 535574 392058
rect 534954 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 535574 356614
rect 534954 356294 535574 356378
rect 534954 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 535574 356294
rect 534954 320614 535574 356058
rect 534954 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 535574 320614
rect 534954 320294 535574 320378
rect 534954 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 535574 320294
rect 534954 284614 535574 320058
rect 534954 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 535574 284614
rect 534954 284294 535574 284378
rect 534954 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 535574 284294
rect 534954 248614 535574 284058
rect 534954 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 535574 248614
rect 534954 248294 535574 248378
rect 534954 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 535574 248294
rect 534954 212614 535574 248058
rect 534954 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 535574 212614
rect 534954 212294 535574 212378
rect 534954 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 535574 212294
rect 534954 176614 535574 212058
rect 534954 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 535574 176614
rect 534954 176294 535574 176378
rect 534954 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 535574 176294
rect 534954 140614 535574 176058
rect 534954 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 535574 140614
rect 534954 140294 535574 140378
rect 534954 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 535574 140294
rect 534954 104614 535574 140058
rect 534954 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 535574 104614
rect 534954 104294 535574 104378
rect 534954 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 535574 104294
rect 534954 68614 535574 104058
rect 534954 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 535574 68614
rect 534954 68294 535574 68378
rect 534954 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 535574 68294
rect 534954 32614 535574 68058
rect 534954 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 535574 32614
rect 534954 32294 535574 32378
rect 534954 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 535574 32294
rect 516954 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 517574 -6106
rect 516954 -6426 517574 -6342
rect 516954 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 517574 -6426
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 32058
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 545514 691174 546134 706202
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 545514 619174 546134 654618
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545514 583174 546134 618618
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 547174 546134 582618
rect 545514 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 546134 547174
rect 545514 546854 546134 546938
rect 545514 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 546134 546854
rect 545514 511174 546134 546618
rect 545514 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 546134 511174
rect 545514 510854 546134 510938
rect 545514 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 546134 510854
rect 545514 475174 546134 510618
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 545514 439174 546134 474618
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 545514 403174 546134 438618
rect 545514 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 546134 403174
rect 545514 402854 546134 402938
rect 545514 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 546134 402854
rect 545514 367174 546134 402618
rect 545514 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 546134 367174
rect 545514 366854 546134 366938
rect 545514 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 546134 366854
rect 545514 331174 546134 366618
rect 545514 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 546134 331174
rect 545514 330854 546134 330938
rect 545514 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 546134 330854
rect 545514 295174 546134 330618
rect 545514 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 546134 295174
rect 545514 294854 546134 294938
rect 545514 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 546134 294854
rect 545514 259174 546134 294618
rect 545514 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 546134 259174
rect 545514 258854 546134 258938
rect 545514 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 546134 258854
rect 545514 223174 546134 258618
rect 545514 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 546134 223174
rect 545514 222854 546134 222938
rect 545514 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 546134 222854
rect 545514 187174 546134 222618
rect 545514 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 546134 187174
rect 545514 186854 546134 186938
rect 545514 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 546134 186854
rect 545514 151174 546134 186618
rect 545514 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 546134 151174
rect 545514 150854 546134 150938
rect 545514 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 546134 150854
rect 545514 115174 546134 150618
rect 545514 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 546134 115174
rect 545514 114854 546134 114938
rect 545514 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 546134 114854
rect 545514 79174 546134 114618
rect 545514 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 546134 79174
rect 545514 78854 546134 78938
rect 545514 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 546134 78854
rect 545514 43174 546134 78618
rect 545514 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546134 43174
rect 545514 42854 546134 42938
rect 545514 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546134 42854
rect 545514 7174 546134 42618
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -2266 546134 6618
rect 545514 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 546134 -2266
rect 545514 -2586 546134 -2502
rect 545514 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 546134 -2586
rect 545514 -3814 546134 -2822
rect 549234 694894 549854 708122
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 658894 549854 694338
rect 549234 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 549854 658894
rect 549234 658574 549854 658658
rect 549234 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 549854 658574
rect 549234 622894 549854 658338
rect 549234 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 549854 622894
rect 549234 622574 549854 622658
rect 549234 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 549854 622574
rect 549234 586894 549854 622338
rect 549234 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 549854 586894
rect 549234 586574 549854 586658
rect 549234 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 549854 586574
rect 549234 550894 549854 586338
rect 549234 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 549854 550894
rect 549234 550574 549854 550658
rect 549234 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 549854 550574
rect 549234 514894 549854 550338
rect 549234 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 549854 514894
rect 549234 514574 549854 514658
rect 549234 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 549854 514574
rect 549234 478894 549854 514338
rect 549234 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 549854 478894
rect 549234 478574 549854 478658
rect 549234 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 549854 478574
rect 549234 442894 549854 478338
rect 549234 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 549854 442894
rect 549234 442574 549854 442658
rect 549234 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 549854 442574
rect 549234 406894 549854 442338
rect 549234 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 549854 406894
rect 549234 406574 549854 406658
rect 549234 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 549854 406574
rect 549234 370894 549854 406338
rect 549234 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 549854 370894
rect 549234 370574 549854 370658
rect 549234 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 549854 370574
rect 549234 334894 549854 370338
rect 549234 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 549854 334894
rect 549234 334574 549854 334658
rect 549234 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 549854 334574
rect 549234 298894 549854 334338
rect 549234 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 549854 298894
rect 549234 298574 549854 298658
rect 549234 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 549854 298574
rect 549234 262894 549854 298338
rect 549234 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 549854 262894
rect 549234 262574 549854 262658
rect 549234 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 549854 262574
rect 549234 226894 549854 262338
rect 549234 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 549854 226894
rect 549234 226574 549854 226658
rect 549234 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 549854 226574
rect 549234 190894 549854 226338
rect 549234 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 549854 190894
rect 549234 190574 549854 190658
rect 549234 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 549854 190574
rect 549234 154894 549854 190338
rect 549234 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 549854 154894
rect 549234 154574 549854 154658
rect 549234 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 549854 154574
rect 549234 118894 549854 154338
rect 549234 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 549854 118894
rect 549234 118574 549854 118658
rect 549234 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 549854 118574
rect 549234 82894 549854 118338
rect 549234 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 549854 82894
rect 549234 82574 549854 82658
rect 549234 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 549854 82574
rect 549234 46894 549854 82338
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 549234 10894 549854 46338
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -4186 549854 10338
rect 549234 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 549854 -4186
rect 549234 -4506 549854 -4422
rect 549234 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 549854 -4506
rect 549234 -5734 549854 -4742
rect 552954 698614 553574 710042
rect 570954 711558 571574 711590
rect 570954 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 571574 711558
rect 570954 711238 571574 711322
rect 570954 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 571574 711238
rect 567234 709638 567854 709670
rect 567234 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 567854 709638
rect 567234 709318 567854 709402
rect 567234 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 567854 709318
rect 563514 707718 564134 707750
rect 563514 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 564134 707718
rect 563514 707398 564134 707482
rect 563514 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 564134 707398
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 552954 626614 553574 662058
rect 552954 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 553574 626614
rect 552954 626294 553574 626378
rect 552954 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 553574 626294
rect 552954 590614 553574 626058
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 552954 554614 553574 590058
rect 552954 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 553574 554614
rect 552954 554294 553574 554378
rect 552954 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 553574 554294
rect 552954 518614 553574 554058
rect 552954 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 553574 518614
rect 552954 518294 553574 518378
rect 552954 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 553574 518294
rect 552954 482614 553574 518058
rect 552954 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 553574 482614
rect 552954 482294 553574 482378
rect 552954 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 553574 482294
rect 552954 446614 553574 482058
rect 552954 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 553574 446614
rect 552954 446294 553574 446378
rect 552954 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 553574 446294
rect 552954 410614 553574 446058
rect 552954 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 553574 410614
rect 552954 410294 553574 410378
rect 552954 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 553574 410294
rect 552954 374614 553574 410058
rect 552954 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 553574 374614
rect 552954 374294 553574 374378
rect 552954 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 553574 374294
rect 552954 338614 553574 374058
rect 552954 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 553574 338614
rect 552954 338294 553574 338378
rect 552954 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 553574 338294
rect 552954 302614 553574 338058
rect 552954 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 553574 302614
rect 552954 302294 553574 302378
rect 552954 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 553574 302294
rect 552954 266614 553574 302058
rect 552954 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 553574 266614
rect 552954 266294 553574 266378
rect 552954 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 553574 266294
rect 552954 230614 553574 266058
rect 552954 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 553574 230614
rect 552954 230294 553574 230378
rect 552954 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 553574 230294
rect 552954 194614 553574 230058
rect 552954 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 553574 194614
rect 552954 194294 553574 194378
rect 552954 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 553574 194294
rect 552954 158614 553574 194058
rect 552954 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 553574 158614
rect 552954 158294 553574 158378
rect 552954 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 553574 158294
rect 552954 122614 553574 158058
rect 552954 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 553574 122614
rect 552954 122294 553574 122378
rect 552954 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 553574 122294
rect 552954 86614 553574 122058
rect 552954 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 553574 86614
rect 552954 86294 553574 86378
rect 552954 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 553574 86294
rect 552954 50614 553574 86058
rect 552954 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 553574 50614
rect 552954 50294 553574 50378
rect 552954 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 553574 50294
rect 552954 14614 553574 50058
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 534954 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 535574 -7066
rect 534954 -7386 535574 -7302
rect 534954 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 535574 -7386
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 14058
rect 559794 705798 560414 705830
rect 559794 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 560414 705798
rect 559794 705478 560414 705562
rect 559794 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 560414 705478
rect 559794 669454 560414 705242
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -1306 560414 20898
rect 559794 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 560414 -1306
rect 559794 -1626 560414 -1542
rect 559794 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 560414 -1626
rect 559794 -1894 560414 -1862
rect 563514 673174 564134 707162
rect 563514 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 564134 673174
rect 563514 672854 564134 672938
rect 563514 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 564134 672854
rect 563514 637174 564134 672618
rect 563514 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 564134 637174
rect 563514 636854 564134 636938
rect 563514 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 564134 636854
rect 563514 601174 564134 636618
rect 563514 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 564134 601174
rect 563514 600854 564134 600938
rect 563514 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 564134 600854
rect 563514 565174 564134 600618
rect 563514 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 564134 565174
rect 563514 564854 564134 564938
rect 563514 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 564134 564854
rect 563514 529174 564134 564618
rect 563514 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 564134 529174
rect 563514 528854 564134 528938
rect 563514 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 564134 528854
rect 563514 493174 564134 528618
rect 563514 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 564134 493174
rect 563514 492854 564134 492938
rect 563514 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 564134 492854
rect 563514 457174 564134 492618
rect 563514 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 564134 457174
rect 563514 456854 564134 456938
rect 563514 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 564134 456854
rect 563514 421174 564134 456618
rect 563514 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 564134 421174
rect 563514 420854 564134 420938
rect 563514 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 564134 420854
rect 563514 385174 564134 420618
rect 563514 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 564134 385174
rect 563514 384854 564134 384938
rect 563514 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 564134 384854
rect 563514 349174 564134 384618
rect 563514 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 564134 349174
rect 563514 348854 564134 348938
rect 563514 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 564134 348854
rect 563514 313174 564134 348618
rect 563514 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 564134 313174
rect 563514 312854 564134 312938
rect 563514 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 564134 312854
rect 563514 277174 564134 312618
rect 563514 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 564134 277174
rect 563514 276854 564134 276938
rect 563514 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 564134 276854
rect 563514 241174 564134 276618
rect 563514 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 564134 241174
rect 563514 240854 564134 240938
rect 563514 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 564134 240854
rect 563514 205174 564134 240618
rect 563514 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 564134 205174
rect 563514 204854 564134 204938
rect 563514 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 564134 204854
rect 563514 169174 564134 204618
rect 563514 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 564134 169174
rect 563514 168854 564134 168938
rect 563514 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 564134 168854
rect 563514 133174 564134 168618
rect 563514 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 564134 133174
rect 563514 132854 564134 132938
rect 563514 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 564134 132854
rect 563514 97174 564134 132618
rect 563514 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 564134 97174
rect 563514 96854 564134 96938
rect 563514 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 564134 96854
rect 563514 61174 564134 96618
rect 563514 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 564134 61174
rect 563514 60854 564134 60938
rect 563514 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 564134 60854
rect 563514 25174 564134 60618
rect 563514 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 564134 25174
rect 563514 24854 564134 24938
rect 563514 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 564134 24854
rect 563514 -3226 564134 24618
rect 563514 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 564134 -3226
rect 563514 -3546 564134 -3462
rect 563514 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 564134 -3546
rect 563514 -3814 564134 -3782
rect 567234 676894 567854 709082
rect 567234 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 567854 676894
rect 567234 676574 567854 676658
rect 567234 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 567854 676574
rect 567234 640894 567854 676338
rect 567234 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 567854 640894
rect 567234 640574 567854 640658
rect 567234 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 567854 640574
rect 567234 604894 567854 640338
rect 567234 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 567854 604894
rect 567234 604574 567854 604658
rect 567234 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 567854 604574
rect 567234 568894 567854 604338
rect 567234 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 567854 568894
rect 567234 568574 567854 568658
rect 567234 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 567854 568574
rect 567234 532894 567854 568338
rect 567234 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 567854 532894
rect 567234 532574 567854 532658
rect 567234 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 567854 532574
rect 567234 496894 567854 532338
rect 567234 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 567854 496894
rect 567234 496574 567854 496658
rect 567234 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 567854 496574
rect 567234 460894 567854 496338
rect 567234 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 567854 460894
rect 567234 460574 567854 460658
rect 567234 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 567854 460574
rect 567234 424894 567854 460338
rect 567234 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 567854 424894
rect 567234 424574 567854 424658
rect 567234 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 567854 424574
rect 567234 388894 567854 424338
rect 567234 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 567854 388894
rect 567234 388574 567854 388658
rect 567234 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 567854 388574
rect 567234 352894 567854 388338
rect 567234 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 567854 352894
rect 567234 352574 567854 352658
rect 567234 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 567854 352574
rect 567234 316894 567854 352338
rect 567234 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 567854 316894
rect 567234 316574 567854 316658
rect 567234 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 567854 316574
rect 567234 280894 567854 316338
rect 567234 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 567854 280894
rect 567234 280574 567854 280658
rect 567234 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 567854 280574
rect 567234 244894 567854 280338
rect 567234 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 567854 244894
rect 567234 244574 567854 244658
rect 567234 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 567854 244574
rect 567234 208894 567854 244338
rect 567234 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 567854 208894
rect 567234 208574 567854 208658
rect 567234 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 567854 208574
rect 567234 172894 567854 208338
rect 567234 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 567854 172894
rect 567234 172574 567854 172658
rect 567234 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 567854 172574
rect 567234 136894 567854 172338
rect 567234 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 567854 136894
rect 567234 136574 567854 136658
rect 567234 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 567854 136574
rect 567234 100894 567854 136338
rect 567234 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 567854 100894
rect 567234 100574 567854 100658
rect 567234 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 567854 100574
rect 567234 64894 567854 100338
rect 567234 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 567854 64894
rect 567234 64574 567854 64658
rect 567234 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 567854 64574
rect 567234 28894 567854 64338
rect 567234 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 567854 28894
rect 567234 28574 567854 28658
rect 567234 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 567854 28574
rect 567234 -5146 567854 28338
rect 567234 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 567854 -5146
rect 567234 -5466 567854 -5382
rect 567234 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 567854 -5466
rect 567234 -5734 567854 -5702
rect 570954 680614 571574 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 581514 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 582134 706758
rect 581514 706438 582134 706522
rect 581514 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 582134 706438
rect 570954 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 571574 680614
rect 570954 680294 571574 680378
rect 570954 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 571574 680294
rect 570954 644614 571574 680058
rect 570954 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 571574 644614
rect 570954 644294 571574 644378
rect 570954 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 571574 644294
rect 570954 608614 571574 644058
rect 570954 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 571574 608614
rect 570954 608294 571574 608378
rect 570954 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 571574 608294
rect 570954 572614 571574 608058
rect 570954 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 571574 572614
rect 570954 572294 571574 572378
rect 570954 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 571574 572294
rect 570954 536614 571574 572058
rect 570954 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 571574 536614
rect 570954 536294 571574 536378
rect 570954 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 571574 536294
rect 570954 500614 571574 536058
rect 570954 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 571574 500614
rect 570954 500294 571574 500378
rect 570954 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 571574 500294
rect 570954 464614 571574 500058
rect 570954 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 571574 464614
rect 570954 464294 571574 464378
rect 570954 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 571574 464294
rect 570954 428614 571574 464058
rect 570954 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 571574 428614
rect 570954 428294 571574 428378
rect 570954 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 571574 428294
rect 570954 392614 571574 428058
rect 570954 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 571574 392614
rect 570954 392294 571574 392378
rect 570954 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 571574 392294
rect 570954 356614 571574 392058
rect 570954 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 571574 356614
rect 570954 356294 571574 356378
rect 570954 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 571574 356294
rect 570954 320614 571574 356058
rect 570954 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 571574 320614
rect 570954 320294 571574 320378
rect 570954 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 571574 320294
rect 570954 284614 571574 320058
rect 570954 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 571574 284614
rect 570954 284294 571574 284378
rect 570954 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 571574 284294
rect 570954 248614 571574 284058
rect 570954 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 571574 248614
rect 570954 248294 571574 248378
rect 570954 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 571574 248294
rect 570954 212614 571574 248058
rect 570954 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 571574 212614
rect 570954 212294 571574 212378
rect 570954 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 571574 212294
rect 570954 176614 571574 212058
rect 570954 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 571574 176614
rect 570954 176294 571574 176378
rect 570954 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 571574 176294
rect 570954 140614 571574 176058
rect 570954 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 571574 140614
rect 570954 140294 571574 140378
rect 570954 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 571574 140294
rect 570954 104614 571574 140058
rect 570954 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 571574 104614
rect 570954 104294 571574 104378
rect 570954 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 571574 104294
rect 570954 68614 571574 104058
rect 570954 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 571574 68614
rect 570954 68294 571574 68378
rect 570954 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 571574 68294
rect 570954 32614 571574 68058
rect 570954 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 571574 32614
rect 570954 32294 571574 32378
rect 570954 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 571574 32294
rect 552954 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 553574 -6106
rect 552954 -6426 553574 -6342
rect 552954 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 553574 -6426
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 32058
rect 577794 704838 578414 705830
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 581514 691174 582134 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -2266 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 587850 691174
rect 587230 690854 587850 690938
rect 587230 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 587850 690854
rect 587230 655174 587850 690618
rect 587230 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 587850 655174
rect 587230 654854 587850 654938
rect 587230 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 587850 654854
rect 587230 619174 587850 654618
rect 587230 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 587850 619174
rect 587230 618854 587850 618938
rect 587230 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 587850 618854
rect 587230 583174 587850 618618
rect 587230 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 587850 583174
rect 587230 582854 587850 582938
rect 587230 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 587850 582854
rect 587230 547174 587850 582618
rect 587230 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 587850 547174
rect 587230 546854 587850 546938
rect 587230 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 587850 546854
rect 587230 511174 587850 546618
rect 587230 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 587850 511174
rect 587230 510854 587850 510938
rect 587230 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 587850 510854
rect 587230 475174 587850 510618
rect 587230 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 587850 475174
rect 587230 474854 587850 474938
rect 587230 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 587850 474854
rect 587230 439174 587850 474618
rect 587230 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 587850 439174
rect 587230 438854 587850 438938
rect 587230 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 587850 438854
rect 587230 403174 587850 438618
rect 587230 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 587850 403174
rect 587230 402854 587850 402938
rect 587230 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 587850 402854
rect 587230 367174 587850 402618
rect 587230 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 587850 367174
rect 587230 366854 587850 366938
rect 587230 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 587850 366854
rect 587230 331174 587850 366618
rect 587230 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 587850 331174
rect 587230 330854 587850 330938
rect 587230 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 587850 330854
rect 587230 295174 587850 330618
rect 587230 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 587850 295174
rect 587230 294854 587850 294938
rect 587230 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 587850 294854
rect 587230 259174 587850 294618
rect 587230 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 587850 259174
rect 587230 258854 587850 258938
rect 587230 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 587850 258854
rect 587230 223174 587850 258618
rect 587230 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 587850 223174
rect 587230 222854 587850 222938
rect 587230 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 587850 222854
rect 587230 187174 587850 222618
rect 587230 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 587850 187174
rect 587230 186854 587850 186938
rect 587230 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 587850 186854
rect 587230 151174 587850 186618
rect 587230 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 587850 151174
rect 587230 150854 587850 150938
rect 587230 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 587850 150854
rect 587230 115174 587850 150618
rect 587230 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 587850 115174
rect 587230 114854 587850 114938
rect 587230 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 587850 114854
rect 587230 79174 587850 114618
rect 587230 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 587850 79174
rect 587230 78854 587850 78938
rect 587230 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 587850 78854
rect 587230 43174 587850 78618
rect 587230 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 587850 43174
rect 587230 42854 587850 42938
rect 587230 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 587850 42854
rect 587230 7174 587850 42618
rect 587230 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 587850 7174
rect 587230 6854 587850 6938
rect 587230 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 587850 6854
rect 581514 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 582134 -2266
rect 581514 -2586 582134 -2502
rect 581514 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 582134 -2586
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect 588190 672854 588810 672938
rect 588190 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect 588190 637174 588810 672618
rect 588190 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect 588190 636854 588810 636938
rect 588190 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect 588190 601174 588810 636618
rect 588190 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect 588190 600854 588810 600938
rect 588190 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect 588190 565174 588810 600618
rect 588190 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect 588190 564854 588810 564938
rect 588190 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect 588190 529174 588810 564618
rect 588190 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect 588190 528854 588810 528938
rect 588190 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect 588190 493174 588810 528618
rect 588190 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect 588190 492854 588810 492938
rect 588190 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect 588190 457174 588810 492618
rect 588190 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect 588190 456854 588810 456938
rect 588190 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect 588190 421174 588810 456618
rect 588190 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 588190 420854 588810 420938
rect 588190 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 588190 385174 588810 420618
rect 588190 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 588190 384854 588810 384938
rect 588190 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 588190 349174 588810 384618
rect 588190 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 588190 348854 588810 348938
rect 588190 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 588190 313174 588810 348618
rect 588190 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 588190 312854 588810 312938
rect 588190 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 588190 277174 588810 312618
rect 588190 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 588190 276854 588810 276938
rect 588190 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 588190 241174 588810 276618
rect 588190 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 588190 240854 588810 240938
rect 588190 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 588190 205174 588810 240618
rect 588190 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 588190 204854 588810 204938
rect 588190 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 588190 169174 588810 204618
rect 588190 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 588190 168854 588810 168938
rect 588190 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 588190 133174 588810 168618
rect 588190 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 588190 132854 588810 132938
rect 588190 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 588190 97174 588810 132618
rect 588190 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 588190 96854 588810 96938
rect 588190 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 588190 61174 588810 96618
rect 588190 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 588190 60854 588810 60938
rect 588190 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 588190 25174 588810 60618
rect 588190 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect 588190 24854 588810 24938
rect 588190 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect 588190 -3226 588810 24618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 589770 694894
rect 589150 694574 589770 694658
rect 589150 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 589770 694574
rect 589150 658894 589770 694338
rect 589150 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 589770 658894
rect 589150 658574 589770 658658
rect 589150 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 589770 658574
rect 589150 622894 589770 658338
rect 589150 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 589770 622894
rect 589150 622574 589770 622658
rect 589150 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 589770 622574
rect 589150 586894 589770 622338
rect 589150 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 589770 586894
rect 589150 586574 589770 586658
rect 589150 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 589770 586574
rect 589150 550894 589770 586338
rect 589150 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 589770 550894
rect 589150 550574 589770 550658
rect 589150 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 589770 550574
rect 589150 514894 589770 550338
rect 589150 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 589770 514894
rect 589150 514574 589770 514658
rect 589150 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 589770 514574
rect 589150 478894 589770 514338
rect 589150 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 589770 478894
rect 589150 478574 589770 478658
rect 589150 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 589770 478574
rect 589150 442894 589770 478338
rect 589150 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 589770 442894
rect 589150 442574 589770 442658
rect 589150 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 589770 442574
rect 589150 406894 589770 442338
rect 589150 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 589770 406894
rect 589150 406574 589770 406658
rect 589150 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 589770 406574
rect 589150 370894 589770 406338
rect 589150 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 589770 370894
rect 589150 370574 589770 370658
rect 589150 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 589770 370574
rect 589150 334894 589770 370338
rect 589150 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 589770 334894
rect 589150 334574 589770 334658
rect 589150 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 589770 334574
rect 589150 298894 589770 334338
rect 589150 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 589770 298894
rect 589150 298574 589770 298658
rect 589150 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 589770 298574
rect 589150 262894 589770 298338
rect 589150 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 589770 262894
rect 589150 262574 589770 262658
rect 589150 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 589770 262574
rect 589150 226894 589770 262338
rect 589150 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 589770 226894
rect 589150 226574 589770 226658
rect 589150 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 589770 226574
rect 589150 190894 589770 226338
rect 589150 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 589770 190894
rect 589150 190574 589770 190658
rect 589150 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 589770 190574
rect 589150 154894 589770 190338
rect 589150 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 589770 154894
rect 589150 154574 589770 154658
rect 589150 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 589770 154574
rect 589150 118894 589770 154338
rect 589150 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 589770 118894
rect 589150 118574 589770 118658
rect 589150 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 589770 118574
rect 589150 82894 589770 118338
rect 589150 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 589770 82894
rect 589150 82574 589770 82658
rect 589150 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 589770 82574
rect 589150 46894 589770 82338
rect 589150 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 589770 46894
rect 589150 46574 589770 46658
rect 589150 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 589770 46574
rect 589150 10894 589770 46338
rect 589150 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 589770 10894
rect 589150 10574 589770 10658
rect 589150 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 589770 10574
rect 589150 -4186 589770 10338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect 590110 676574 590730 676658
rect 590110 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect 590110 640894 590730 676338
rect 590110 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect 590110 640574 590730 640658
rect 590110 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect 590110 604894 590730 640338
rect 590110 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect 590110 604574 590730 604658
rect 590110 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect 590110 568894 590730 604338
rect 590110 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect 590110 568574 590730 568658
rect 590110 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect 590110 532894 590730 568338
rect 590110 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect 590110 532574 590730 532658
rect 590110 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect 590110 496894 590730 532338
rect 590110 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect 590110 496574 590730 496658
rect 590110 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect 590110 460894 590730 496338
rect 590110 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect 590110 460574 590730 460658
rect 590110 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect 590110 424894 590730 460338
rect 590110 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 590110 424574 590730 424658
rect 590110 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 590110 388894 590730 424338
rect 590110 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 590110 388574 590730 388658
rect 590110 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 590110 352894 590730 388338
rect 590110 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 590110 352574 590730 352658
rect 590110 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 590110 316894 590730 352338
rect 590110 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 590110 316574 590730 316658
rect 590110 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 590110 280894 590730 316338
rect 590110 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 590110 280574 590730 280658
rect 590110 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 590110 244894 590730 280338
rect 590110 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 590110 244574 590730 244658
rect 590110 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 590110 208894 590730 244338
rect 590110 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 590110 208574 590730 208658
rect 590110 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 590110 172894 590730 208338
rect 590110 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 590110 172574 590730 172658
rect 590110 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 590110 136894 590730 172338
rect 590110 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 590110 136574 590730 136658
rect 590110 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 590110 100894 590730 136338
rect 590110 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 590110 100574 590730 100658
rect 590110 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 590110 64894 590730 100338
rect 590110 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 590110 64574 590730 64658
rect 590110 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 590110 28894 590730 64338
rect 590110 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect 590110 28574 590730 28658
rect 590110 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect 590110 -5146 590730 28338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 591690 698614
rect 591070 698294 591690 698378
rect 591070 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 591690 698294
rect 591070 662614 591690 698058
rect 591070 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 591690 662614
rect 591070 662294 591690 662378
rect 591070 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 591690 662294
rect 591070 626614 591690 662058
rect 591070 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 591690 626614
rect 591070 626294 591690 626378
rect 591070 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 591690 626294
rect 591070 590614 591690 626058
rect 591070 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 591690 590614
rect 591070 590294 591690 590378
rect 591070 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 591690 590294
rect 591070 554614 591690 590058
rect 591070 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 591690 554614
rect 591070 554294 591690 554378
rect 591070 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 591690 554294
rect 591070 518614 591690 554058
rect 591070 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 591690 518614
rect 591070 518294 591690 518378
rect 591070 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 591690 518294
rect 591070 482614 591690 518058
rect 591070 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 591690 482614
rect 591070 482294 591690 482378
rect 591070 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 591690 482294
rect 591070 446614 591690 482058
rect 591070 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 591690 446614
rect 591070 446294 591690 446378
rect 591070 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 591690 446294
rect 591070 410614 591690 446058
rect 591070 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 591690 410614
rect 591070 410294 591690 410378
rect 591070 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 591690 410294
rect 591070 374614 591690 410058
rect 591070 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 591690 374614
rect 591070 374294 591690 374378
rect 591070 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 591690 374294
rect 591070 338614 591690 374058
rect 591070 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 591690 338614
rect 591070 338294 591690 338378
rect 591070 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 591690 338294
rect 591070 302614 591690 338058
rect 591070 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 591690 302614
rect 591070 302294 591690 302378
rect 591070 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 591690 302294
rect 591070 266614 591690 302058
rect 591070 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 591690 266614
rect 591070 266294 591690 266378
rect 591070 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 591690 266294
rect 591070 230614 591690 266058
rect 591070 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 591690 230614
rect 591070 230294 591690 230378
rect 591070 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 591690 230294
rect 591070 194614 591690 230058
rect 591070 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 591690 194614
rect 591070 194294 591690 194378
rect 591070 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 591690 194294
rect 591070 158614 591690 194058
rect 591070 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 591690 158614
rect 591070 158294 591690 158378
rect 591070 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 591690 158294
rect 591070 122614 591690 158058
rect 591070 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 591690 122614
rect 591070 122294 591690 122378
rect 591070 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 591690 122294
rect 591070 86614 591690 122058
rect 591070 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 591690 86614
rect 591070 86294 591690 86378
rect 591070 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 591690 86294
rect 591070 50614 591690 86058
rect 591070 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 591690 50614
rect 591070 50294 591690 50378
rect 591070 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 591690 50294
rect 591070 14614 591690 50058
rect 591070 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 591690 14614
rect 591070 14294 591690 14378
rect 591070 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 591690 14294
rect 591070 -6106 591690 14058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect 592030 680294 592650 680378
rect 592030 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect 592030 644614 592650 680058
rect 592030 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect 592030 644294 592650 644378
rect 592030 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect 592030 608614 592650 644058
rect 592030 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect 592030 608294 592650 608378
rect 592030 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect 592030 572614 592650 608058
rect 592030 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect 592030 572294 592650 572378
rect 592030 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect 592030 536614 592650 572058
rect 592030 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect 592030 536294 592650 536378
rect 592030 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect 592030 500614 592650 536058
rect 592030 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect 592030 500294 592650 500378
rect 592030 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect 592030 464614 592650 500058
rect 592030 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect 592030 464294 592650 464378
rect 592030 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect 592030 428614 592650 464058
rect 592030 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 592030 428294 592650 428378
rect 592030 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 592030 392614 592650 428058
rect 592030 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 592030 392294 592650 392378
rect 592030 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 592030 356614 592650 392058
rect 592030 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 592030 356294 592650 356378
rect 592030 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 592030 320614 592650 356058
rect 592030 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 592030 320294 592650 320378
rect 592030 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 592030 284614 592650 320058
rect 592030 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 592030 284294 592650 284378
rect 592030 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 592030 248614 592650 284058
rect 592030 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 592030 248294 592650 248378
rect 592030 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 592030 212614 592650 248058
rect 592030 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 592030 212294 592650 212378
rect 592030 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 592030 176614 592650 212058
rect 592030 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 592030 176294 592650 176378
rect 592030 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 592030 140614 592650 176058
rect 592030 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 592030 140294 592650 140378
rect 592030 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 592030 104614 592650 140058
rect 592030 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 592030 104294 592650 104378
rect 592030 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 592030 68614 592650 104058
rect 592030 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 592030 68294 592650 68378
rect 592030 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 592030 32614 592650 68058
rect 592030 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect 592030 32294 592650 32378
rect 592030 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect 570954 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 571574 -7066
rect 570954 -7386 571574 -7302
rect 570954 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 571574 -7386
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 680378 -8458 680614
rect -8374 680378 -8138 680614
rect -8694 680058 -8458 680294
rect -8374 680058 -8138 680294
rect -8694 644378 -8458 644614
rect -8374 644378 -8138 644614
rect -8694 644058 -8458 644294
rect -8374 644058 -8138 644294
rect -8694 608378 -8458 608614
rect -8374 608378 -8138 608614
rect -8694 608058 -8458 608294
rect -8374 608058 -8138 608294
rect -8694 572378 -8458 572614
rect -8374 572378 -8138 572614
rect -8694 572058 -8458 572294
rect -8374 572058 -8138 572294
rect -8694 536378 -8458 536614
rect -8374 536378 -8138 536614
rect -8694 536058 -8458 536294
rect -8374 536058 -8138 536294
rect -8694 500378 -8458 500614
rect -8374 500378 -8138 500614
rect -8694 500058 -8458 500294
rect -8374 500058 -8138 500294
rect -8694 464378 -8458 464614
rect -8374 464378 -8138 464614
rect -8694 464058 -8458 464294
rect -8374 464058 -8138 464294
rect -8694 428378 -8458 428614
rect -8374 428378 -8138 428614
rect -8694 428058 -8458 428294
rect -8374 428058 -8138 428294
rect -8694 392378 -8458 392614
rect -8374 392378 -8138 392614
rect -8694 392058 -8458 392294
rect -8374 392058 -8138 392294
rect -8694 356378 -8458 356614
rect -8374 356378 -8138 356614
rect -8694 356058 -8458 356294
rect -8374 356058 -8138 356294
rect -8694 320378 -8458 320614
rect -8374 320378 -8138 320614
rect -8694 320058 -8458 320294
rect -8374 320058 -8138 320294
rect -8694 284378 -8458 284614
rect -8374 284378 -8138 284614
rect -8694 284058 -8458 284294
rect -8374 284058 -8138 284294
rect -8694 248378 -8458 248614
rect -8374 248378 -8138 248614
rect -8694 248058 -8458 248294
rect -8374 248058 -8138 248294
rect -8694 212378 -8458 212614
rect -8374 212378 -8138 212614
rect -8694 212058 -8458 212294
rect -8374 212058 -8138 212294
rect -8694 176378 -8458 176614
rect -8374 176378 -8138 176614
rect -8694 176058 -8458 176294
rect -8374 176058 -8138 176294
rect -8694 140378 -8458 140614
rect -8374 140378 -8138 140614
rect -8694 140058 -8458 140294
rect -8374 140058 -8138 140294
rect -8694 104378 -8458 104614
rect -8374 104378 -8138 104614
rect -8694 104058 -8458 104294
rect -8374 104058 -8138 104294
rect -8694 68378 -8458 68614
rect -8374 68378 -8138 68614
rect -8694 68058 -8458 68294
rect -8374 68058 -8138 68294
rect -8694 32378 -8458 32614
rect -8374 32378 -8138 32614
rect -8694 32058 -8458 32294
rect -8374 32058 -8138 32294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12986 710362 13222 710598
rect 13306 710362 13542 710598
rect 12986 710042 13222 710278
rect 13306 710042 13542 710278
rect -7734 698378 -7498 698614
rect -7414 698378 -7178 698614
rect -7734 698058 -7498 698294
rect -7414 698058 -7178 698294
rect -7734 662378 -7498 662614
rect -7414 662378 -7178 662614
rect -7734 662058 -7498 662294
rect -7414 662058 -7178 662294
rect -7734 626378 -7498 626614
rect -7414 626378 -7178 626614
rect -7734 626058 -7498 626294
rect -7414 626058 -7178 626294
rect -7734 590378 -7498 590614
rect -7414 590378 -7178 590614
rect -7734 590058 -7498 590294
rect -7414 590058 -7178 590294
rect -7734 554378 -7498 554614
rect -7414 554378 -7178 554614
rect -7734 554058 -7498 554294
rect -7414 554058 -7178 554294
rect -7734 518378 -7498 518614
rect -7414 518378 -7178 518614
rect -7734 518058 -7498 518294
rect -7414 518058 -7178 518294
rect -7734 482378 -7498 482614
rect -7414 482378 -7178 482614
rect -7734 482058 -7498 482294
rect -7414 482058 -7178 482294
rect -7734 446378 -7498 446614
rect -7414 446378 -7178 446614
rect -7734 446058 -7498 446294
rect -7414 446058 -7178 446294
rect -7734 410378 -7498 410614
rect -7414 410378 -7178 410614
rect -7734 410058 -7498 410294
rect -7414 410058 -7178 410294
rect -7734 374378 -7498 374614
rect -7414 374378 -7178 374614
rect -7734 374058 -7498 374294
rect -7414 374058 -7178 374294
rect -7734 338378 -7498 338614
rect -7414 338378 -7178 338614
rect -7734 338058 -7498 338294
rect -7414 338058 -7178 338294
rect -7734 302378 -7498 302614
rect -7414 302378 -7178 302614
rect -7734 302058 -7498 302294
rect -7414 302058 -7178 302294
rect -7734 266378 -7498 266614
rect -7414 266378 -7178 266614
rect -7734 266058 -7498 266294
rect -7414 266058 -7178 266294
rect -7734 230378 -7498 230614
rect -7414 230378 -7178 230614
rect -7734 230058 -7498 230294
rect -7414 230058 -7178 230294
rect -7734 194378 -7498 194614
rect -7414 194378 -7178 194614
rect -7734 194058 -7498 194294
rect -7414 194058 -7178 194294
rect -7734 158378 -7498 158614
rect -7414 158378 -7178 158614
rect -7734 158058 -7498 158294
rect -7414 158058 -7178 158294
rect -7734 122378 -7498 122614
rect -7414 122378 -7178 122614
rect -7734 122058 -7498 122294
rect -7414 122058 -7178 122294
rect -7734 86378 -7498 86614
rect -7414 86378 -7178 86614
rect -7734 86058 -7498 86294
rect -7414 86058 -7178 86294
rect -7734 50378 -7498 50614
rect -7414 50378 -7178 50614
rect -7734 50058 -7498 50294
rect -7414 50058 -7178 50294
rect -7734 14378 -7498 14614
rect -7414 14378 -7178 14614
rect -7734 14058 -7498 14294
rect -7414 14058 -7178 14294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 676658 -6538 676894
rect -6454 676658 -6218 676894
rect -6774 676338 -6538 676574
rect -6454 676338 -6218 676574
rect -6774 640658 -6538 640894
rect -6454 640658 -6218 640894
rect -6774 640338 -6538 640574
rect -6454 640338 -6218 640574
rect -6774 604658 -6538 604894
rect -6454 604658 -6218 604894
rect -6774 604338 -6538 604574
rect -6454 604338 -6218 604574
rect -6774 568658 -6538 568894
rect -6454 568658 -6218 568894
rect -6774 568338 -6538 568574
rect -6454 568338 -6218 568574
rect -6774 532658 -6538 532894
rect -6454 532658 -6218 532894
rect -6774 532338 -6538 532574
rect -6454 532338 -6218 532574
rect -6774 496658 -6538 496894
rect -6454 496658 -6218 496894
rect -6774 496338 -6538 496574
rect -6454 496338 -6218 496574
rect -6774 460658 -6538 460894
rect -6454 460658 -6218 460894
rect -6774 460338 -6538 460574
rect -6454 460338 -6218 460574
rect -6774 424658 -6538 424894
rect -6454 424658 -6218 424894
rect -6774 424338 -6538 424574
rect -6454 424338 -6218 424574
rect -6774 388658 -6538 388894
rect -6454 388658 -6218 388894
rect -6774 388338 -6538 388574
rect -6454 388338 -6218 388574
rect -6774 352658 -6538 352894
rect -6454 352658 -6218 352894
rect -6774 352338 -6538 352574
rect -6454 352338 -6218 352574
rect -6774 316658 -6538 316894
rect -6454 316658 -6218 316894
rect -6774 316338 -6538 316574
rect -6454 316338 -6218 316574
rect -6774 280658 -6538 280894
rect -6454 280658 -6218 280894
rect -6774 280338 -6538 280574
rect -6454 280338 -6218 280574
rect -6774 244658 -6538 244894
rect -6454 244658 -6218 244894
rect -6774 244338 -6538 244574
rect -6454 244338 -6218 244574
rect -6774 208658 -6538 208894
rect -6454 208658 -6218 208894
rect -6774 208338 -6538 208574
rect -6454 208338 -6218 208574
rect -6774 172658 -6538 172894
rect -6454 172658 -6218 172894
rect -6774 172338 -6538 172574
rect -6454 172338 -6218 172574
rect -6774 136658 -6538 136894
rect -6454 136658 -6218 136894
rect -6774 136338 -6538 136574
rect -6454 136338 -6218 136574
rect -6774 100658 -6538 100894
rect -6454 100658 -6218 100894
rect -6774 100338 -6538 100574
rect -6454 100338 -6218 100574
rect -6774 64658 -6538 64894
rect -6454 64658 -6218 64894
rect -6774 64338 -6538 64574
rect -6454 64338 -6218 64574
rect -6774 28658 -6538 28894
rect -6454 28658 -6218 28894
rect -6774 28338 -6538 28574
rect -6454 28338 -6218 28574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 9266 708442 9502 708678
rect 9586 708442 9822 708678
rect 9266 708122 9502 708358
rect 9586 708122 9822 708358
rect -5814 694658 -5578 694894
rect -5494 694658 -5258 694894
rect -5814 694338 -5578 694574
rect -5494 694338 -5258 694574
rect -5814 658658 -5578 658894
rect -5494 658658 -5258 658894
rect -5814 658338 -5578 658574
rect -5494 658338 -5258 658574
rect -5814 622658 -5578 622894
rect -5494 622658 -5258 622894
rect -5814 622338 -5578 622574
rect -5494 622338 -5258 622574
rect -5814 586658 -5578 586894
rect -5494 586658 -5258 586894
rect -5814 586338 -5578 586574
rect -5494 586338 -5258 586574
rect -5814 550658 -5578 550894
rect -5494 550658 -5258 550894
rect -5814 550338 -5578 550574
rect -5494 550338 -5258 550574
rect -5814 514658 -5578 514894
rect -5494 514658 -5258 514894
rect -5814 514338 -5578 514574
rect -5494 514338 -5258 514574
rect -5814 478658 -5578 478894
rect -5494 478658 -5258 478894
rect -5814 478338 -5578 478574
rect -5494 478338 -5258 478574
rect -5814 442658 -5578 442894
rect -5494 442658 -5258 442894
rect -5814 442338 -5578 442574
rect -5494 442338 -5258 442574
rect -5814 406658 -5578 406894
rect -5494 406658 -5258 406894
rect -5814 406338 -5578 406574
rect -5494 406338 -5258 406574
rect -5814 370658 -5578 370894
rect -5494 370658 -5258 370894
rect -5814 370338 -5578 370574
rect -5494 370338 -5258 370574
rect -5814 334658 -5578 334894
rect -5494 334658 -5258 334894
rect -5814 334338 -5578 334574
rect -5494 334338 -5258 334574
rect -5814 298658 -5578 298894
rect -5494 298658 -5258 298894
rect -5814 298338 -5578 298574
rect -5494 298338 -5258 298574
rect -5814 262658 -5578 262894
rect -5494 262658 -5258 262894
rect -5814 262338 -5578 262574
rect -5494 262338 -5258 262574
rect -5814 226658 -5578 226894
rect -5494 226658 -5258 226894
rect -5814 226338 -5578 226574
rect -5494 226338 -5258 226574
rect -5814 190658 -5578 190894
rect -5494 190658 -5258 190894
rect -5814 190338 -5578 190574
rect -5494 190338 -5258 190574
rect -5814 154658 -5578 154894
rect -5494 154658 -5258 154894
rect -5814 154338 -5578 154574
rect -5494 154338 -5258 154574
rect -5814 118658 -5578 118894
rect -5494 118658 -5258 118894
rect -5814 118338 -5578 118574
rect -5494 118338 -5258 118574
rect -5814 82658 -5578 82894
rect -5494 82658 -5258 82894
rect -5814 82338 -5578 82574
rect -5494 82338 -5258 82574
rect -5814 46658 -5578 46894
rect -5494 46658 -5258 46894
rect -5814 46338 -5578 46574
rect -5494 46338 -5258 46574
rect -5814 10658 -5578 10894
rect -5494 10658 -5258 10894
rect -5814 10338 -5578 10574
rect -5494 10338 -5258 10574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 672938 -4618 673174
rect -4534 672938 -4298 673174
rect -4854 672618 -4618 672854
rect -4534 672618 -4298 672854
rect -4854 636938 -4618 637174
rect -4534 636938 -4298 637174
rect -4854 636618 -4618 636854
rect -4534 636618 -4298 636854
rect -4854 600938 -4618 601174
rect -4534 600938 -4298 601174
rect -4854 600618 -4618 600854
rect -4534 600618 -4298 600854
rect -4854 564938 -4618 565174
rect -4534 564938 -4298 565174
rect -4854 564618 -4618 564854
rect -4534 564618 -4298 564854
rect -4854 528938 -4618 529174
rect -4534 528938 -4298 529174
rect -4854 528618 -4618 528854
rect -4534 528618 -4298 528854
rect -4854 492938 -4618 493174
rect -4534 492938 -4298 493174
rect -4854 492618 -4618 492854
rect -4534 492618 -4298 492854
rect -4854 456938 -4618 457174
rect -4534 456938 -4298 457174
rect -4854 456618 -4618 456854
rect -4534 456618 -4298 456854
rect -4854 420938 -4618 421174
rect -4534 420938 -4298 421174
rect -4854 420618 -4618 420854
rect -4534 420618 -4298 420854
rect -4854 384938 -4618 385174
rect -4534 384938 -4298 385174
rect -4854 384618 -4618 384854
rect -4534 384618 -4298 384854
rect -4854 348938 -4618 349174
rect -4534 348938 -4298 349174
rect -4854 348618 -4618 348854
rect -4534 348618 -4298 348854
rect -4854 312938 -4618 313174
rect -4534 312938 -4298 313174
rect -4854 312618 -4618 312854
rect -4534 312618 -4298 312854
rect -4854 276938 -4618 277174
rect -4534 276938 -4298 277174
rect -4854 276618 -4618 276854
rect -4534 276618 -4298 276854
rect -4854 240938 -4618 241174
rect -4534 240938 -4298 241174
rect -4854 240618 -4618 240854
rect -4534 240618 -4298 240854
rect -4854 204938 -4618 205174
rect -4534 204938 -4298 205174
rect -4854 204618 -4618 204854
rect -4534 204618 -4298 204854
rect -4854 168938 -4618 169174
rect -4534 168938 -4298 169174
rect -4854 168618 -4618 168854
rect -4534 168618 -4298 168854
rect -4854 132938 -4618 133174
rect -4534 132938 -4298 133174
rect -4854 132618 -4618 132854
rect -4534 132618 -4298 132854
rect -4854 96938 -4618 97174
rect -4534 96938 -4298 97174
rect -4854 96618 -4618 96854
rect -4534 96618 -4298 96854
rect -4854 60938 -4618 61174
rect -4534 60938 -4298 61174
rect -4854 60618 -4618 60854
rect -4534 60618 -4298 60854
rect -4854 24938 -4618 25174
rect -4534 24938 -4298 25174
rect -4854 24618 -4618 24854
rect -4534 24618 -4298 24854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 5546 706522 5782 706758
rect 5866 706522 6102 706758
rect 5546 706202 5782 706438
rect 5866 706202 6102 706438
rect -3894 690938 -3658 691174
rect -3574 690938 -3338 691174
rect -3894 690618 -3658 690854
rect -3574 690618 -3338 690854
rect -3894 654938 -3658 655174
rect -3574 654938 -3338 655174
rect -3894 654618 -3658 654854
rect -3574 654618 -3338 654854
rect -3894 618938 -3658 619174
rect -3574 618938 -3338 619174
rect -3894 618618 -3658 618854
rect -3574 618618 -3338 618854
rect -3894 582938 -3658 583174
rect -3574 582938 -3338 583174
rect -3894 582618 -3658 582854
rect -3574 582618 -3338 582854
rect -3894 546938 -3658 547174
rect -3574 546938 -3338 547174
rect -3894 546618 -3658 546854
rect -3574 546618 -3338 546854
rect -3894 510938 -3658 511174
rect -3574 510938 -3338 511174
rect -3894 510618 -3658 510854
rect -3574 510618 -3338 510854
rect -3894 474938 -3658 475174
rect -3574 474938 -3338 475174
rect -3894 474618 -3658 474854
rect -3574 474618 -3338 474854
rect -3894 438938 -3658 439174
rect -3574 438938 -3338 439174
rect -3894 438618 -3658 438854
rect -3574 438618 -3338 438854
rect -3894 402938 -3658 403174
rect -3574 402938 -3338 403174
rect -3894 402618 -3658 402854
rect -3574 402618 -3338 402854
rect -3894 366938 -3658 367174
rect -3574 366938 -3338 367174
rect -3894 366618 -3658 366854
rect -3574 366618 -3338 366854
rect -3894 330938 -3658 331174
rect -3574 330938 -3338 331174
rect -3894 330618 -3658 330854
rect -3574 330618 -3338 330854
rect -3894 294938 -3658 295174
rect -3574 294938 -3338 295174
rect -3894 294618 -3658 294854
rect -3574 294618 -3338 294854
rect -3894 258938 -3658 259174
rect -3574 258938 -3338 259174
rect -3894 258618 -3658 258854
rect -3574 258618 -3338 258854
rect -3894 222938 -3658 223174
rect -3574 222938 -3338 223174
rect -3894 222618 -3658 222854
rect -3574 222618 -3338 222854
rect -3894 186938 -3658 187174
rect -3574 186938 -3338 187174
rect -3894 186618 -3658 186854
rect -3574 186618 -3338 186854
rect -3894 150938 -3658 151174
rect -3574 150938 -3338 151174
rect -3894 150618 -3658 150854
rect -3574 150618 -3338 150854
rect -3894 114938 -3658 115174
rect -3574 114938 -3338 115174
rect -3894 114618 -3658 114854
rect -3574 114618 -3338 114854
rect -3894 78938 -3658 79174
rect -3574 78938 -3338 79174
rect -3894 78618 -3658 78854
rect -3574 78618 -3338 78854
rect -3894 42938 -3658 43174
rect -3574 42938 -3338 43174
rect -3894 42618 -3658 42854
rect -3574 42618 -3338 42854
rect -3894 6938 -3658 7174
rect -3574 6938 -3338 7174
rect -3894 6618 -3658 6854
rect -3574 6618 -3338 6854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 5546 -2502 5782 -2266
rect 5866 -2502 6102 -2266
rect 5546 -2822 5782 -2586
rect 5866 -2822 6102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 9266 -4422 9502 -4186
rect 9586 -4422 9822 -4186
rect 9266 -4742 9502 -4506
rect 9586 -4742 9822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect 30986 711322 31222 711558
rect 31306 711322 31542 711558
rect 30986 711002 31222 711238
rect 31306 711002 31542 711238
rect 27266 709402 27502 709638
rect 27586 709402 27822 709638
rect 27266 709082 27502 709318
rect 27586 709082 27822 709318
rect 23546 707482 23782 707718
rect 23866 707482 24102 707718
rect 23546 707162 23782 707398
rect 23866 707162 24102 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -1542 20062 -1306
rect 20146 -1542 20382 -1306
rect 19826 -1862 20062 -1626
rect 20146 -1862 20382 -1626
rect 23546 672938 23782 673174
rect 23866 672938 24102 673174
rect 23546 672618 23782 672854
rect 23866 672618 24102 672854
rect 23546 636938 23782 637174
rect 23866 636938 24102 637174
rect 23546 636618 23782 636854
rect 23866 636618 24102 636854
rect 23546 600938 23782 601174
rect 23866 600938 24102 601174
rect 23546 600618 23782 600854
rect 23866 600618 24102 600854
rect 23546 564938 23782 565174
rect 23866 564938 24102 565174
rect 23546 564618 23782 564854
rect 23866 564618 24102 564854
rect 23546 528938 23782 529174
rect 23866 528938 24102 529174
rect 23546 528618 23782 528854
rect 23866 528618 24102 528854
rect 23546 492938 23782 493174
rect 23866 492938 24102 493174
rect 23546 492618 23782 492854
rect 23866 492618 24102 492854
rect 23546 456938 23782 457174
rect 23866 456938 24102 457174
rect 23546 456618 23782 456854
rect 23866 456618 24102 456854
rect 23546 420938 23782 421174
rect 23866 420938 24102 421174
rect 23546 420618 23782 420854
rect 23866 420618 24102 420854
rect 23546 384938 23782 385174
rect 23866 384938 24102 385174
rect 23546 384618 23782 384854
rect 23866 384618 24102 384854
rect 23546 348938 23782 349174
rect 23866 348938 24102 349174
rect 23546 348618 23782 348854
rect 23866 348618 24102 348854
rect 23546 312938 23782 313174
rect 23866 312938 24102 313174
rect 23546 312618 23782 312854
rect 23866 312618 24102 312854
rect 23546 276938 23782 277174
rect 23866 276938 24102 277174
rect 23546 276618 23782 276854
rect 23866 276618 24102 276854
rect 23546 240938 23782 241174
rect 23866 240938 24102 241174
rect 23546 240618 23782 240854
rect 23866 240618 24102 240854
rect 23546 204938 23782 205174
rect 23866 204938 24102 205174
rect 23546 204618 23782 204854
rect 23866 204618 24102 204854
rect 23546 168938 23782 169174
rect 23866 168938 24102 169174
rect 23546 168618 23782 168854
rect 23866 168618 24102 168854
rect 23546 132938 23782 133174
rect 23866 132938 24102 133174
rect 23546 132618 23782 132854
rect 23866 132618 24102 132854
rect 23546 96938 23782 97174
rect 23866 96938 24102 97174
rect 23546 96618 23782 96854
rect 23866 96618 24102 96854
rect 23546 60938 23782 61174
rect 23866 60938 24102 61174
rect 23546 60618 23782 60854
rect 23866 60618 24102 60854
rect 23546 24938 23782 25174
rect 23866 24938 24102 25174
rect 23546 24618 23782 24854
rect 23866 24618 24102 24854
rect 23546 -3462 23782 -3226
rect 23866 -3462 24102 -3226
rect 23546 -3782 23782 -3546
rect 23866 -3782 24102 -3546
rect 27266 676658 27502 676894
rect 27586 676658 27822 676894
rect 27266 676338 27502 676574
rect 27586 676338 27822 676574
rect 27266 640658 27502 640894
rect 27586 640658 27822 640894
rect 27266 640338 27502 640574
rect 27586 640338 27822 640574
rect 27266 604658 27502 604894
rect 27586 604658 27822 604894
rect 27266 604338 27502 604574
rect 27586 604338 27822 604574
rect 27266 568658 27502 568894
rect 27586 568658 27822 568894
rect 27266 568338 27502 568574
rect 27586 568338 27822 568574
rect 27266 532658 27502 532894
rect 27586 532658 27822 532894
rect 27266 532338 27502 532574
rect 27586 532338 27822 532574
rect 27266 496658 27502 496894
rect 27586 496658 27822 496894
rect 27266 496338 27502 496574
rect 27586 496338 27822 496574
rect 27266 460658 27502 460894
rect 27586 460658 27822 460894
rect 27266 460338 27502 460574
rect 27586 460338 27822 460574
rect 27266 424658 27502 424894
rect 27586 424658 27822 424894
rect 27266 424338 27502 424574
rect 27586 424338 27822 424574
rect 27266 388658 27502 388894
rect 27586 388658 27822 388894
rect 27266 388338 27502 388574
rect 27586 388338 27822 388574
rect 27266 352658 27502 352894
rect 27586 352658 27822 352894
rect 27266 352338 27502 352574
rect 27586 352338 27822 352574
rect 27266 316658 27502 316894
rect 27586 316658 27822 316894
rect 27266 316338 27502 316574
rect 27586 316338 27822 316574
rect 27266 280658 27502 280894
rect 27586 280658 27822 280894
rect 27266 280338 27502 280574
rect 27586 280338 27822 280574
rect 27266 244658 27502 244894
rect 27586 244658 27822 244894
rect 27266 244338 27502 244574
rect 27586 244338 27822 244574
rect 27266 208658 27502 208894
rect 27586 208658 27822 208894
rect 27266 208338 27502 208574
rect 27586 208338 27822 208574
rect 27266 172658 27502 172894
rect 27586 172658 27822 172894
rect 27266 172338 27502 172574
rect 27586 172338 27822 172574
rect 27266 136658 27502 136894
rect 27586 136658 27822 136894
rect 27266 136338 27502 136574
rect 27586 136338 27822 136574
rect 27266 100658 27502 100894
rect 27586 100658 27822 100894
rect 27266 100338 27502 100574
rect 27586 100338 27822 100574
rect 27266 64658 27502 64894
rect 27586 64658 27822 64894
rect 27266 64338 27502 64574
rect 27586 64338 27822 64574
rect 27266 28658 27502 28894
rect 27586 28658 27822 28894
rect 27266 28338 27502 28574
rect 27586 28338 27822 28574
rect 27266 -5382 27502 -5146
rect 27586 -5382 27822 -5146
rect 27266 -5702 27502 -5466
rect 27586 -5702 27822 -5466
rect 48986 710362 49222 710598
rect 49306 710362 49542 710598
rect 48986 710042 49222 710278
rect 49306 710042 49542 710278
rect 45266 708442 45502 708678
rect 45586 708442 45822 708678
rect 45266 708122 45502 708358
rect 45586 708122 45822 708358
rect 41546 706522 41782 706758
rect 41866 706522 42102 706758
rect 41546 706202 41782 706438
rect 41866 706202 42102 706438
rect 30986 680378 31222 680614
rect 31306 680378 31542 680614
rect 30986 680058 31222 680294
rect 31306 680058 31542 680294
rect 30986 644378 31222 644614
rect 31306 644378 31542 644614
rect 30986 644058 31222 644294
rect 31306 644058 31542 644294
rect 30986 608378 31222 608614
rect 31306 608378 31542 608614
rect 30986 608058 31222 608294
rect 31306 608058 31542 608294
rect 30986 572378 31222 572614
rect 31306 572378 31542 572614
rect 30986 572058 31222 572294
rect 31306 572058 31542 572294
rect 30986 536378 31222 536614
rect 31306 536378 31542 536614
rect 30986 536058 31222 536294
rect 31306 536058 31542 536294
rect 30986 500378 31222 500614
rect 31306 500378 31542 500614
rect 30986 500058 31222 500294
rect 31306 500058 31542 500294
rect 30986 464378 31222 464614
rect 31306 464378 31542 464614
rect 30986 464058 31222 464294
rect 31306 464058 31542 464294
rect 30986 428378 31222 428614
rect 31306 428378 31542 428614
rect 30986 428058 31222 428294
rect 31306 428058 31542 428294
rect 30986 392378 31222 392614
rect 31306 392378 31542 392614
rect 30986 392058 31222 392294
rect 31306 392058 31542 392294
rect 30986 356378 31222 356614
rect 31306 356378 31542 356614
rect 30986 356058 31222 356294
rect 31306 356058 31542 356294
rect 30986 320378 31222 320614
rect 31306 320378 31542 320614
rect 30986 320058 31222 320294
rect 31306 320058 31542 320294
rect 30986 284378 31222 284614
rect 31306 284378 31542 284614
rect 30986 284058 31222 284294
rect 31306 284058 31542 284294
rect 30986 248378 31222 248614
rect 31306 248378 31542 248614
rect 30986 248058 31222 248294
rect 31306 248058 31542 248294
rect 30986 212378 31222 212614
rect 31306 212378 31542 212614
rect 30986 212058 31222 212294
rect 31306 212058 31542 212294
rect 30986 176378 31222 176614
rect 31306 176378 31542 176614
rect 30986 176058 31222 176294
rect 31306 176058 31542 176294
rect 30986 140378 31222 140614
rect 31306 140378 31542 140614
rect 30986 140058 31222 140294
rect 31306 140058 31542 140294
rect 30986 104378 31222 104614
rect 31306 104378 31542 104614
rect 30986 104058 31222 104294
rect 31306 104058 31542 104294
rect 30986 68378 31222 68614
rect 31306 68378 31542 68614
rect 30986 68058 31222 68294
rect 31306 68058 31542 68294
rect 30986 32378 31222 32614
rect 31306 32378 31542 32614
rect 30986 32058 31222 32294
rect 31306 32058 31542 32294
rect 12986 -6342 13222 -6106
rect 13306 -6342 13542 -6106
rect 12986 -6662 13222 -6426
rect 13306 -6662 13542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 41546 654938 41782 655174
rect 41866 654938 42102 655174
rect 41546 654618 41782 654854
rect 41866 654618 42102 654854
rect 41546 618938 41782 619174
rect 41866 618938 42102 619174
rect 41546 618618 41782 618854
rect 41866 618618 42102 618854
rect 41546 582938 41782 583174
rect 41866 582938 42102 583174
rect 41546 582618 41782 582854
rect 41866 582618 42102 582854
rect 41546 546938 41782 547174
rect 41866 546938 42102 547174
rect 41546 546618 41782 546854
rect 41866 546618 42102 546854
rect 41546 510938 41782 511174
rect 41866 510938 42102 511174
rect 41546 510618 41782 510854
rect 41866 510618 42102 510854
rect 41546 474938 41782 475174
rect 41866 474938 42102 475174
rect 41546 474618 41782 474854
rect 41866 474618 42102 474854
rect 41546 438938 41782 439174
rect 41866 438938 42102 439174
rect 41546 438618 41782 438854
rect 41866 438618 42102 438854
rect 41546 402938 41782 403174
rect 41866 402938 42102 403174
rect 41546 402618 41782 402854
rect 41866 402618 42102 402854
rect 41546 366938 41782 367174
rect 41866 366938 42102 367174
rect 41546 366618 41782 366854
rect 41866 366618 42102 366854
rect 41546 330938 41782 331174
rect 41866 330938 42102 331174
rect 41546 330618 41782 330854
rect 41866 330618 42102 330854
rect 41546 294938 41782 295174
rect 41866 294938 42102 295174
rect 41546 294618 41782 294854
rect 41866 294618 42102 294854
rect 41546 258938 41782 259174
rect 41866 258938 42102 259174
rect 41546 258618 41782 258854
rect 41866 258618 42102 258854
rect 41546 222938 41782 223174
rect 41866 222938 42102 223174
rect 41546 222618 41782 222854
rect 41866 222618 42102 222854
rect 41546 186938 41782 187174
rect 41866 186938 42102 187174
rect 41546 186618 41782 186854
rect 41866 186618 42102 186854
rect 41546 150938 41782 151174
rect 41866 150938 42102 151174
rect 41546 150618 41782 150854
rect 41866 150618 42102 150854
rect 41546 114938 41782 115174
rect 41866 114938 42102 115174
rect 41546 114618 41782 114854
rect 41866 114618 42102 114854
rect 41546 78938 41782 79174
rect 41866 78938 42102 79174
rect 41546 78618 41782 78854
rect 41866 78618 42102 78854
rect 41546 42938 41782 43174
rect 41866 42938 42102 43174
rect 41546 42618 41782 42854
rect 41866 42618 42102 42854
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -2502 41782 -2266
rect 41866 -2502 42102 -2266
rect 41546 -2822 41782 -2586
rect 41866 -2822 42102 -2586
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 45266 658658 45502 658894
rect 45586 658658 45822 658894
rect 45266 658338 45502 658574
rect 45586 658338 45822 658574
rect 45266 622658 45502 622894
rect 45586 622658 45822 622894
rect 45266 622338 45502 622574
rect 45586 622338 45822 622574
rect 45266 586658 45502 586894
rect 45586 586658 45822 586894
rect 45266 586338 45502 586574
rect 45586 586338 45822 586574
rect 45266 550658 45502 550894
rect 45586 550658 45822 550894
rect 45266 550338 45502 550574
rect 45586 550338 45822 550574
rect 45266 514658 45502 514894
rect 45586 514658 45822 514894
rect 45266 514338 45502 514574
rect 45586 514338 45822 514574
rect 45266 478658 45502 478894
rect 45586 478658 45822 478894
rect 45266 478338 45502 478574
rect 45586 478338 45822 478574
rect 45266 442658 45502 442894
rect 45586 442658 45822 442894
rect 45266 442338 45502 442574
rect 45586 442338 45822 442574
rect 45266 406658 45502 406894
rect 45586 406658 45822 406894
rect 45266 406338 45502 406574
rect 45586 406338 45822 406574
rect 45266 370658 45502 370894
rect 45586 370658 45822 370894
rect 45266 370338 45502 370574
rect 45586 370338 45822 370574
rect 45266 334658 45502 334894
rect 45586 334658 45822 334894
rect 45266 334338 45502 334574
rect 45586 334338 45822 334574
rect 45266 298658 45502 298894
rect 45586 298658 45822 298894
rect 45266 298338 45502 298574
rect 45586 298338 45822 298574
rect 45266 262658 45502 262894
rect 45586 262658 45822 262894
rect 45266 262338 45502 262574
rect 45586 262338 45822 262574
rect 45266 226658 45502 226894
rect 45586 226658 45822 226894
rect 45266 226338 45502 226574
rect 45586 226338 45822 226574
rect 45266 190658 45502 190894
rect 45586 190658 45822 190894
rect 45266 190338 45502 190574
rect 45586 190338 45822 190574
rect 45266 154658 45502 154894
rect 45586 154658 45822 154894
rect 45266 154338 45502 154574
rect 45586 154338 45822 154574
rect 45266 118658 45502 118894
rect 45586 118658 45822 118894
rect 45266 118338 45502 118574
rect 45586 118338 45822 118574
rect 45266 82658 45502 82894
rect 45586 82658 45822 82894
rect 45266 82338 45502 82574
rect 45586 82338 45822 82574
rect 45266 46658 45502 46894
rect 45586 46658 45822 46894
rect 45266 46338 45502 46574
rect 45586 46338 45822 46574
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -4422 45502 -4186
rect 45586 -4422 45822 -4186
rect 45266 -4742 45502 -4506
rect 45586 -4742 45822 -4506
rect 66986 711322 67222 711558
rect 67306 711322 67542 711558
rect 66986 711002 67222 711238
rect 67306 711002 67542 711238
rect 63266 709402 63502 709638
rect 63586 709402 63822 709638
rect 63266 709082 63502 709318
rect 63586 709082 63822 709318
rect 59546 707482 59782 707718
rect 59866 707482 60102 707718
rect 59546 707162 59782 707398
rect 59866 707162 60102 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 48986 662378 49222 662614
rect 49306 662378 49542 662614
rect 48986 662058 49222 662294
rect 49306 662058 49542 662294
rect 48986 626378 49222 626614
rect 49306 626378 49542 626614
rect 48986 626058 49222 626294
rect 49306 626058 49542 626294
rect 48986 590378 49222 590614
rect 49306 590378 49542 590614
rect 48986 590058 49222 590294
rect 49306 590058 49542 590294
rect 48986 554378 49222 554614
rect 49306 554378 49542 554614
rect 48986 554058 49222 554294
rect 49306 554058 49542 554294
rect 48986 518378 49222 518614
rect 49306 518378 49542 518614
rect 48986 518058 49222 518294
rect 49306 518058 49542 518294
rect 48986 482378 49222 482614
rect 49306 482378 49542 482614
rect 48986 482058 49222 482294
rect 49306 482058 49542 482294
rect 48986 446378 49222 446614
rect 49306 446378 49542 446614
rect 48986 446058 49222 446294
rect 49306 446058 49542 446294
rect 48986 410378 49222 410614
rect 49306 410378 49542 410614
rect 48986 410058 49222 410294
rect 49306 410058 49542 410294
rect 48986 374378 49222 374614
rect 49306 374378 49542 374614
rect 48986 374058 49222 374294
rect 49306 374058 49542 374294
rect 48986 338378 49222 338614
rect 49306 338378 49542 338614
rect 48986 338058 49222 338294
rect 49306 338058 49542 338294
rect 48986 302378 49222 302614
rect 49306 302378 49542 302614
rect 48986 302058 49222 302294
rect 49306 302058 49542 302294
rect 48986 266378 49222 266614
rect 49306 266378 49542 266614
rect 48986 266058 49222 266294
rect 49306 266058 49542 266294
rect 48986 230378 49222 230614
rect 49306 230378 49542 230614
rect 48986 230058 49222 230294
rect 49306 230058 49542 230294
rect 48986 194378 49222 194614
rect 49306 194378 49542 194614
rect 48986 194058 49222 194294
rect 49306 194058 49542 194294
rect 48986 158378 49222 158614
rect 49306 158378 49542 158614
rect 48986 158058 49222 158294
rect 49306 158058 49542 158294
rect 48986 122378 49222 122614
rect 49306 122378 49542 122614
rect 48986 122058 49222 122294
rect 49306 122058 49542 122294
rect 48986 86378 49222 86614
rect 49306 86378 49542 86614
rect 48986 86058 49222 86294
rect 49306 86058 49542 86294
rect 48986 50378 49222 50614
rect 49306 50378 49542 50614
rect 48986 50058 49222 50294
rect 49306 50058 49542 50294
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 30986 -7302 31222 -7066
rect 31306 -7302 31542 -7066
rect 30986 -7622 31222 -7386
rect 31306 -7622 31542 -7386
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 59546 672938 59782 673174
rect 59866 672938 60102 673174
rect 59546 672618 59782 672854
rect 59866 672618 60102 672854
rect 59546 636938 59782 637174
rect 59866 636938 60102 637174
rect 59546 636618 59782 636854
rect 59866 636618 60102 636854
rect 59546 600938 59782 601174
rect 59866 600938 60102 601174
rect 59546 600618 59782 600854
rect 59866 600618 60102 600854
rect 59546 564938 59782 565174
rect 59866 564938 60102 565174
rect 59546 564618 59782 564854
rect 59866 564618 60102 564854
rect 59546 528938 59782 529174
rect 59866 528938 60102 529174
rect 59546 528618 59782 528854
rect 59866 528618 60102 528854
rect 59546 492938 59782 493174
rect 59866 492938 60102 493174
rect 59546 492618 59782 492854
rect 59866 492618 60102 492854
rect 63266 676658 63502 676894
rect 63586 676658 63822 676894
rect 63266 676338 63502 676574
rect 63586 676338 63822 676574
rect 63266 640658 63502 640894
rect 63586 640658 63822 640894
rect 63266 640338 63502 640574
rect 63586 640338 63822 640574
rect 63266 604658 63502 604894
rect 63586 604658 63822 604894
rect 63266 604338 63502 604574
rect 63586 604338 63822 604574
rect 63266 568658 63502 568894
rect 63586 568658 63822 568894
rect 63266 568338 63502 568574
rect 63586 568338 63822 568574
rect 63266 532658 63502 532894
rect 63586 532658 63822 532894
rect 63266 532338 63502 532574
rect 63586 532338 63822 532574
rect 63266 496658 63502 496894
rect 63586 496658 63822 496894
rect 63266 496338 63502 496574
rect 63586 496338 63822 496574
rect 84986 710362 85222 710598
rect 85306 710362 85542 710598
rect 84986 710042 85222 710278
rect 85306 710042 85542 710278
rect 81266 708442 81502 708678
rect 81586 708442 81822 708678
rect 81266 708122 81502 708358
rect 81586 708122 81822 708358
rect 77546 706522 77782 706758
rect 77866 706522 78102 706758
rect 77546 706202 77782 706438
rect 77866 706202 78102 706438
rect 66986 680378 67222 680614
rect 67306 680378 67542 680614
rect 66986 680058 67222 680294
rect 67306 680058 67542 680294
rect 66986 644378 67222 644614
rect 67306 644378 67542 644614
rect 66986 644058 67222 644294
rect 67306 644058 67542 644294
rect 66986 608378 67222 608614
rect 67306 608378 67542 608614
rect 66986 608058 67222 608294
rect 67306 608058 67542 608294
rect 66986 572378 67222 572614
rect 67306 572378 67542 572614
rect 66986 572058 67222 572294
rect 67306 572058 67542 572294
rect 66986 536378 67222 536614
rect 67306 536378 67542 536614
rect 66986 536058 67222 536294
rect 67306 536058 67542 536294
rect 66986 500378 67222 500614
rect 67306 500378 67542 500614
rect 66986 500058 67222 500294
rect 67306 500058 67542 500294
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 77546 654938 77782 655174
rect 77866 654938 78102 655174
rect 77546 654618 77782 654854
rect 77866 654618 78102 654854
rect 77546 618938 77782 619174
rect 77866 618938 78102 619174
rect 77546 618618 77782 618854
rect 77866 618618 78102 618854
rect 77546 582938 77782 583174
rect 77866 582938 78102 583174
rect 77546 582618 77782 582854
rect 77866 582618 78102 582854
rect 77546 546938 77782 547174
rect 77866 546938 78102 547174
rect 77546 546618 77782 546854
rect 77866 546618 78102 546854
rect 77546 510938 77782 511174
rect 77866 510938 78102 511174
rect 77546 510618 77782 510854
rect 77866 510618 78102 510854
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 81266 658658 81502 658894
rect 81586 658658 81822 658894
rect 81266 658338 81502 658574
rect 81586 658338 81822 658574
rect 81266 622658 81502 622894
rect 81586 622658 81822 622894
rect 81266 622338 81502 622574
rect 81586 622338 81822 622574
rect 81266 586658 81502 586894
rect 81586 586658 81822 586894
rect 81266 586338 81502 586574
rect 81586 586338 81822 586574
rect 81266 550658 81502 550894
rect 81586 550658 81822 550894
rect 81266 550338 81502 550574
rect 81586 550338 81822 550574
rect 81266 514658 81502 514894
rect 81586 514658 81822 514894
rect 81266 514338 81502 514574
rect 81586 514338 81822 514574
rect 102986 711322 103222 711558
rect 103306 711322 103542 711558
rect 102986 711002 103222 711238
rect 103306 711002 103542 711238
rect 99266 709402 99502 709638
rect 99586 709402 99822 709638
rect 99266 709082 99502 709318
rect 99586 709082 99822 709318
rect 95546 707482 95782 707718
rect 95866 707482 96102 707718
rect 95546 707162 95782 707398
rect 95866 707162 96102 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 84986 662378 85222 662614
rect 85306 662378 85542 662614
rect 84986 662058 85222 662294
rect 85306 662058 85542 662294
rect 84986 626378 85222 626614
rect 85306 626378 85542 626614
rect 84986 626058 85222 626294
rect 85306 626058 85542 626294
rect 84986 590378 85222 590614
rect 85306 590378 85542 590614
rect 84986 590058 85222 590294
rect 85306 590058 85542 590294
rect 84986 554378 85222 554614
rect 85306 554378 85542 554614
rect 84986 554058 85222 554294
rect 85306 554058 85542 554294
rect 84986 518378 85222 518614
rect 85306 518378 85542 518614
rect 84986 518058 85222 518294
rect 85306 518058 85542 518294
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 95546 672938 95782 673174
rect 95866 672938 96102 673174
rect 95546 672618 95782 672854
rect 95866 672618 96102 672854
rect 95546 636938 95782 637174
rect 95866 636938 96102 637174
rect 95546 636618 95782 636854
rect 95866 636618 96102 636854
rect 95546 600938 95782 601174
rect 95866 600938 96102 601174
rect 95546 600618 95782 600854
rect 95866 600618 96102 600854
rect 95546 564938 95782 565174
rect 95866 564938 96102 565174
rect 95546 564618 95782 564854
rect 95866 564618 96102 564854
rect 95546 528938 95782 529174
rect 95866 528938 96102 529174
rect 95546 528618 95782 528854
rect 95866 528618 96102 528854
rect 99266 676658 99502 676894
rect 99586 676658 99822 676894
rect 99266 676338 99502 676574
rect 99586 676338 99822 676574
rect 99266 640658 99502 640894
rect 99586 640658 99822 640894
rect 99266 640338 99502 640574
rect 99586 640338 99822 640574
rect 99266 604658 99502 604894
rect 99586 604658 99822 604894
rect 99266 604338 99502 604574
rect 99586 604338 99822 604574
rect 99266 568658 99502 568894
rect 99586 568658 99822 568894
rect 99266 568338 99502 568574
rect 99586 568338 99822 568574
rect 99266 532658 99502 532894
rect 99586 532658 99822 532894
rect 99266 532338 99502 532574
rect 99586 532338 99822 532574
rect 95546 492938 95782 493174
rect 95866 492938 96102 493174
rect 95546 492618 95782 492854
rect 95866 492618 96102 492854
rect 120986 710362 121222 710598
rect 121306 710362 121542 710598
rect 120986 710042 121222 710278
rect 121306 710042 121542 710278
rect 117266 708442 117502 708678
rect 117586 708442 117822 708678
rect 117266 708122 117502 708358
rect 117586 708122 117822 708358
rect 113546 706522 113782 706758
rect 113866 706522 114102 706758
rect 113546 706202 113782 706438
rect 113866 706202 114102 706438
rect 102986 680378 103222 680614
rect 103306 680378 103542 680614
rect 102986 680058 103222 680294
rect 103306 680058 103542 680294
rect 102986 644378 103222 644614
rect 103306 644378 103542 644614
rect 102986 644058 103222 644294
rect 103306 644058 103542 644294
rect 102986 608378 103222 608614
rect 103306 608378 103542 608614
rect 102986 608058 103222 608294
rect 103306 608058 103542 608294
rect 102986 572378 103222 572614
rect 103306 572378 103542 572614
rect 102986 572058 103222 572294
rect 103306 572058 103542 572294
rect 102986 536378 103222 536614
rect 103306 536378 103542 536614
rect 102986 536058 103222 536294
rect 103306 536058 103542 536294
rect 99266 496658 99502 496894
rect 99586 496658 99822 496894
rect 99266 496338 99502 496574
rect 99586 496338 99822 496574
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 102986 500378 103222 500614
rect 103306 500378 103542 500614
rect 102986 500058 103222 500294
rect 103306 500058 103542 500294
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 113546 654938 113782 655174
rect 113866 654938 114102 655174
rect 113546 654618 113782 654854
rect 113866 654618 114102 654854
rect 113546 618938 113782 619174
rect 113866 618938 114102 619174
rect 113546 618618 113782 618854
rect 113866 618618 114102 618854
rect 113546 582938 113782 583174
rect 113866 582938 114102 583174
rect 113546 582618 113782 582854
rect 113866 582618 114102 582854
rect 113546 546938 113782 547174
rect 113866 546938 114102 547174
rect 113546 546618 113782 546854
rect 113866 546618 114102 546854
rect 113546 510938 113782 511174
rect 113866 510938 114102 511174
rect 113546 510618 113782 510854
rect 113866 510618 114102 510854
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 117266 658658 117502 658894
rect 117586 658658 117822 658894
rect 117266 658338 117502 658574
rect 117586 658338 117822 658574
rect 117266 622658 117502 622894
rect 117586 622658 117822 622894
rect 117266 622338 117502 622574
rect 117586 622338 117822 622574
rect 117266 586658 117502 586894
rect 117586 586658 117822 586894
rect 117266 586338 117502 586574
rect 117586 586338 117822 586574
rect 117266 550658 117502 550894
rect 117586 550658 117822 550894
rect 117266 550338 117502 550574
rect 117586 550338 117822 550574
rect 117266 514658 117502 514894
rect 117586 514658 117822 514894
rect 117266 514338 117502 514574
rect 117586 514338 117822 514574
rect 138986 711322 139222 711558
rect 139306 711322 139542 711558
rect 138986 711002 139222 711238
rect 139306 711002 139542 711238
rect 135266 709402 135502 709638
rect 135586 709402 135822 709638
rect 135266 709082 135502 709318
rect 135586 709082 135822 709318
rect 131546 707482 131782 707718
rect 131866 707482 132102 707718
rect 131546 707162 131782 707398
rect 131866 707162 132102 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 120986 662378 121222 662614
rect 121306 662378 121542 662614
rect 120986 662058 121222 662294
rect 121306 662058 121542 662294
rect 120986 626378 121222 626614
rect 121306 626378 121542 626614
rect 120986 626058 121222 626294
rect 121306 626058 121542 626294
rect 120986 590378 121222 590614
rect 121306 590378 121542 590614
rect 120986 590058 121222 590294
rect 121306 590058 121542 590294
rect 120986 554378 121222 554614
rect 121306 554378 121542 554614
rect 120986 554058 121222 554294
rect 121306 554058 121542 554294
rect 120986 518378 121222 518614
rect 121306 518378 121542 518614
rect 120986 518058 121222 518294
rect 121306 518058 121542 518294
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 131546 672938 131782 673174
rect 131866 672938 132102 673174
rect 131546 672618 131782 672854
rect 131866 672618 132102 672854
rect 131546 636938 131782 637174
rect 131866 636938 132102 637174
rect 131546 636618 131782 636854
rect 131866 636618 132102 636854
rect 131546 600938 131782 601174
rect 131866 600938 132102 601174
rect 131546 600618 131782 600854
rect 131866 600618 132102 600854
rect 131546 564938 131782 565174
rect 131866 564938 132102 565174
rect 131546 564618 131782 564854
rect 131866 564618 132102 564854
rect 131546 528938 131782 529174
rect 131866 528938 132102 529174
rect 131546 528618 131782 528854
rect 131866 528618 132102 528854
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 135266 676658 135502 676894
rect 135586 676658 135822 676894
rect 135266 676338 135502 676574
rect 135586 676338 135822 676574
rect 135266 640658 135502 640894
rect 135586 640658 135822 640894
rect 135266 640338 135502 640574
rect 135586 640338 135822 640574
rect 135266 604658 135502 604894
rect 135586 604658 135822 604894
rect 135266 604338 135502 604574
rect 135586 604338 135822 604574
rect 135266 568658 135502 568894
rect 135586 568658 135822 568894
rect 135266 568338 135502 568574
rect 135586 568338 135822 568574
rect 135266 532658 135502 532894
rect 135586 532658 135822 532894
rect 135266 532338 135502 532574
rect 135586 532338 135822 532574
rect 131546 492938 131782 493174
rect 131866 492938 132102 493174
rect 131546 492618 131782 492854
rect 131866 492618 132102 492854
rect 135266 496658 135502 496894
rect 135586 496658 135822 496894
rect 135266 496338 135502 496574
rect 135586 496338 135822 496574
rect 156986 710362 157222 710598
rect 157306 710362 157542 710598
rect 156986 710042 157222 710278
rect 157306 710042 157542 710278
rect 153266 708442 153502 708678
rect 153586 708442 153822 708678
rect 153266 708122 153502 708358
rect 153586 708122 153822 708358
rect 149546 706522 149782 706758
rect 149866 706522 150102 706758
rect 149546 706202 149782 706438
rect 149866 706202 150102 706438
rect 138986 680378 139222 680614
rect 139306 680378 139542 680614
rect 138986 680058 139222 680294
rect 139306 680058 139542 680294
rect 138986 644378 139222 644614
rect 139306 644378 139542 644614
rect 138986 644058 139222 644294
rect 139306 644058 139542 644294
rect 138986 608378 139222 608614
rect 139306 608378 139542 608614
rect 138986 608058 139222 608294
rect 139306 608058 139542 608294
rect 138986 572378 139222 572614
rect 139306 572378 139542 572614
rect 138986 572058 139222 572294
rect 139306 572058 139542 572294
rect 138986 536378 139222 536614
rect 139306 536378 139542 536614
rect 138986 536058 139222 536294
rect 139306 536058 139542 536294
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 138986 500378 139222 500614
rect 139306 500378 139542 500614
rect 138986 500058 139222 500294
rect 139306 500058 139542 500294
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 149546 654938 149782 655174
rect 149866 654938 150102 655174
rect 149546 654618 149782 654854
rect 149866 654618 150102 654854
rect 149546 618938 149782 619174
rect 149866 618938 150102 619174
rect 149546 618618 149782 618854
rect 149866 618618 150102 618854
rect 149546 582938 149782 583174
rect 149866 582938 150102 583174
rect 149546 582618 149782 582854
rect 149866 582618 150102 582854
rect 149546 546938 149782 547174
rect 149866 546938 150102 547174
rect 149546 546618 149782 546854
rect 149866 546618 150102 546854
rect 149546 510938 149782 511174
rect 149866 510938 150102 511174
rect 149546 510618 149782 510854
rect 149866 510618 150102 510854
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 153266 658658 153502 658894
rect 153586 658658 153822 658894
rect 153266 658338 153502 658574
rect 153586 658338 153822 658574
rect 153266 622658 153502 622894
rect 153586 622658 153822 622894
rect 153266 622338 153502 622574
rect 153586 622338 153822 622574
rect 153266 586658 153502 586894
rect 153586 586658 153822 586894
rect 153266 586338 153502 586574
rect 153586 586338 153822 586574
rect 153266 550658 153502 550894
rect 153586 550658 153822 550894
rect 153266 550338 153502 550574
rect 153586 550338 153822 550574
rect 153266 514658 153502 514894
rect 153586 514658 153822 514894
rect 153266 514338 153502 514574
rect 153586 514338 153822 514574
rect 174986 711322 175222 711558
rect 175306 711322 175542 711558
rect 174986 711002 175222 711238
rect 175306 711002 175542 711238
rect 171266 709402 171502 709638
rect 171586 709402 171822 709638
rect 171266 709082 171502 709318
rect 171586 709082 171822 709318
rect 167546 707482 167782 707718
rect 167866 707482 168102 707718
rect 167546 707162 167782 707398
rect 167866 707162 168102 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 156986 662378 157222 662614
rect 157306 662378 157542 662614
rect 156986 662058 157222 662294
rect 157306 662058 157542 662294
rect 156986 626378 157222 626614
rect 157306 626378 157542 626614
rect 156986 626058 157222 626294
rect 157306 626058 157542 626294
rect 156986 590378 157222 590614
rect 157306 590378 157542 590614
rect 156986 590058 157222 590294
rect 157306 590058 157542 590294
rect 156986 554378 157222 554614
rect 157306 554378 157542 554614
rect 156986 554058 157222 554294
rect 157306 554058 157542 554294
rect 156986 518378 157222 518614
rect 157306 518378 157542 518614
rect 156986 518058 157222 518294
rect 157306 518058 157542 518294
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 167546 672938 167782 673174
rect 167866 672938 168102 673174
rect 167546 672618 167782 672854
rect 167866 672618 168102 672854
rect 167546 636938 167782 637174
rect 167866 636938 168102 637174
rect 167546 636618 167782 636854
rect 167866 636618 168102 636854
rect 167546 600938 167782 601174
rect 167866 600938 168102 601174
rect 167546 600618 167782 600854
rect 167866 600618 168102 600854
rect 167546 564938 167782 565174
rect 167866 564938 168102 565174
rect 167546 564618 167782 564854
rect 167866 564618 168102 564854
rect 167546 528938 167782 529174
rect 167866 528938 168102 529174
rect 167546 528618 167782 528854
rect 167866 528618 168102 528854
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 167546 492938 167782 493174
rect 167866 492938 168102 493174
rect 167546 492618 167782 492854
rect 167866 492618 168102 492854
rect 171266 676658 171502 676894
rect 171586 676658 171822 676894
rect 171266 676338 171502 676574
rect 171586 676338 171822 676574
rect 171266 640658 171502 640894
rect 171586 640658 171822 640894
rect 171266 640338 171502 640574
rect 171586 640338 171822 640574
rect 171266 604658 171502 604894
rect 171586 604658 171822 604894
rect 171266 604338 171502 604574
rect 171586 604338 171822 604574
rect 171266 568658 171502 568894
rect 171586 568658 171822 568894
rect 171266 568338 171502 568574
rect 171586 568338 171822 568574
rect 171266 532658 171502 532894
rect 171586 532658 171822 532894
rect 171266 532338 171502 532574
rect 171586 532338 171822 532574
rect 171266 496658 171502 496894
rect 171586 496658 171822 496894
rect 171266 496338 171502 496574
rect 171586 496338 171822 496574
rect 192986 710362 193222 710598
rect 193306 710362 193542 710598
rect 192986 710042 193222 710278
rect 193306 710042 193542 710278
rect 189266 708442 189502 708678
rect 189586 708442 189822 708678
rect 189266 708122 189502 708358
rect 189586 708122 189822 708358
rect 185546 706522 185782 706758
rect 185866 706522 186102 706758
rect 185546 706202 185782 706438
rect 185866 706202 186102 706438
rect 174986 680378 175222 680614
rect 175306 680378 175542 680614
rect 174986 680058 175222 680294
rect 175306 680058 175542 680294
rect 174986 644378 175222 644614
rect 175306 644378 175542 644614
rect 174986 644058 175222 644294
rect 175306 644058 175542 644294
rect 174986 608378 175222 608614
rect 175306 608378 175542 608614
rect 174986 608058 175222 608294
rect 175306 608058 175542 608294
rect 174986 572378 175222 572614
rect 175306 572378 175542 572614
rect 174986 572058 175222 572294
rect 175306 572058 175542 572294
rect 174986 536378 175222 536614
rect 175306 536378 175542 536614
rect 174986 536058 175222 536294
rect 175306 536058 175542 536294
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 174986 500378 175222 500614
rect 175306 500378 175542 500614
rect 174986 500058 175222 500294
rect 175306 500058 175542 500294
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 185546 654938 185782 655174
rect 185866 654938 186102 655174
rect 185546 654618 185782 654854
rect 185866 654618 186102 654854
rect 185546 618938 185782 619174
rect 185866 618938 186102 619174
rect 185546 618618 185782 618854
rect 185866 618618 186102 618854
rect 185546 582938 185782 583174
rect 185866 582938 186102 583174
rect 185546 582618 185782 582854
rect 185866 582618 186102 582854
rect 185546 546938 185782 547174
rect 185866 546938 186102 547174
rect 185546 546618 185782 546854
rect 185866 546618 186102 546854
rect 185546 510938 185782 511174
rect 185866 510938 186102 511174
rect 185546 510618 185782 510854
rect 185866 510618 186102 510854
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 189266 658658 189502 658894
rect 189586 658658 189822 658894
rect 189266 658338 189502 658574
rect 189586 658338 189822 658574
rect 189266 622658 189502 622894
rect 189586 622658 189822 622894
rect 189266 622338 189502 622574
rect 189586 622338 189822 622574
rect 189266 586658 189502 586894
rect 189586 586658 189822 586894
rect 189266 586338 189502 586574
rect 189586 586338 189822 586574
rect 189266 550658 189502 550894
rect 189586 550658 189822 550894
rect 189266 550338 189502 550574
rect 189586 550338 189822 550574
rect 189266 514658 189502 514894
rect 189586 514658 189822 514894
rect 189266 514338 189502 514574
rect 189586 514338 189822 514574
rect 210986 711322 211222 711558
rect 211306 711322 211542 711558
rect 210986 711002 211222 711238
rect 211306 711002 211542 711238
rect 207266 709402 207502 709638
rect 207586 709402 207822 709638
rect 207266 709082 207502 709318
rect 207586 709082 207822 709318
rect 203546 707482 203782 707718
rect 203866 707482 204102 707718
rect 203546 707162 203782 707398
rect 203866 707162 204102 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 192986 662378 193222 662614
rect 193306 662378 193542 662614
rect 192986 662058 193222 662294
rect 193306 662058 193542 662294
rect 192986 626378 193222 626614
rect 193306 626378 193542 626614
rect 192986 626058 193222 626294
rect 193306 626058 193542 626294
rect 192986 590378 193222 590614
rect 193306 590378 193542 590614
rect 192986 590058 193222 590294
rect 193306 590058 193542 590294
rect 192986 554378 193222 554614
rect 193306 554378 193542 554614
rect 192986 554058 193222 554294
rect 193306 554058 193542 554294
rect 192986 518378 193222 518614
rect 193306 518378 193542 518614
rect 192986 518058 193222 518294
rect 193306 518058 193542 518294
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 61008 471218 61244 471454
rect 61008 470898 61244 471134
rect 195376 471218 195612 471454
rect 195376 470898 195612 471134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 60328 453218 60564 453454
rect 60328 452898 60564 453134
rect 196056 453218 196292 453454
rect 196056 452898 196292 453134
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 61008 435218 61244 435454
rect 61008 434898 61244 435134
rect 195376 435218 195612 435454
rect 195376 434898 195612 435134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 60328 417218 60564 417454
rect 60328 416898 60564 417134
rect 196056 417218 196292 417454
rect 196056 416898 196292 417134
rect 199826 417218 200062 417454
rect 200146 417218 200382 417454
rect 199826 416898 200062 417134
rect 200146 416898 200382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 59546 384938 59782 385174
rect 59866 384938 60102 385174
rect 59546 384618 59782 384854
rect 59866 384618 60102 384854
rect 59546 348938 59782 349174
rect 59866 348938 60102 349174
rect 59546 348618 59782 348854
rect 59866 348618 60102 348854
rect 59546 312938 59782 313174
rect 59866 312938 60102 313174
rect 59546 312618 59782 312854
rect 59866 312618 60102 312854
rect 59546 276938 59782 277174
rect 59866 276938 60102 277174
rect 59546 276618 59782 276854
rect 59866 276618 60102 276854
rect 59546 240938 59782 241174
rect 59866 240938 60102 241174
rect 59546 240618 59782 240854
rect 59866 240618 60102 240854
rect 63266 388658 63502 388894
rect 63586 388658 63822 388894
rect 63266 388338 63502 388574
rect 63586 388338 63822 388574
rect 63266 352658 63502 352894
rect 63586 352658 63822 352894
rect 63266 352338 63502 352574
rect 63586 352338 63822 352574
rect 63266 316658 63502 316894
rect 63586 316658 63822 316894
rect 63266 316338 63502 316574
rect 63586 316338 63822 316574
rect 63266 280658 63502 280894
rect 63586 280658 63822 280894
rect 63266 280338 63502 280574
rect 63586 280338 63822 280574
rect 63266 244658 63502 244894
rect 63586 244658 63822 244894
rect 63266 244338 63502 244574
rect 63586 244338 63822 244574
rect 66986 392378 67222 392614
rect 67306 392378 67542 392614
rect 66986 392058 67222 392294
rect 67306 392058 67542 392294
rect 66986 356378 67222 356614
rect 67306 356378 67542 356614
rect 66986 356058 67222 356294
rect 67306 356058 67542 356294
rect 66986 320378 67222 320614
rect 67306 320378 67542 320614
rect 66986 320058 67222 320294
rect 67306 320058 67542 320294
rect 66986 284378 67222 284614
rect 67306 284378 67542 284614
rect 66986 284058 67222 284294
rect 67306 284058 67542 284294
rect 66986 248378 67222 248614
rect 67306 248378 67542 248614
rect 66986 248058 67222 248294
rect 67306 248058 67542 248294
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 73826 291218 74062 291454
rect 74146 291218 74382 291454
rect 73826 290898 74062 291134
rect 74146 290898 74382 291134
rect 73826 255218 74062 255454
rect 74146 255218 74382 255454
rect 73826 254898 74062 255134
rect 74146 254898 74382 255134
rect 77546 366938 77782 367174
rect 77866 366938 78102 367174
rect 77546 366618 77782 366854
rect 77866 366618 78102 366854
rect 77546 330938 77782 331174
rect 77866 330938 78102 331174
rect 77546 330618 77782 330854
rect 77866 330618 78102 330854
rect 77546 294938 77782 295174
rect 77866 294938 78102 295174
rect 77546 294618 77782 294854
rect 77866 294618 78102 294854
rect 77546 258938 77782 259174
rect 77866 258938 78102 259174
rect 77546 258618 77782 258854
rect 77866 258618 78102 258854
rect 81266 370658 81502 370894
rect 81586 370658 81822 370894
rect 81266 370338 81502 370574
rect 81586 370338 81822 370574
rect 81266 334658 81502 334894
rect 81586 334658 81822 334894
rect 81266 334338 81502 334574
rect 81586 334338 81822 334574
rect 81266 298658 81502 298894
rect 81586 298658 81822 298894
rect 81266 298338 81502 298574
rect 81586 298338 81822 298574
rect 81266 262658 81502 262894
rect 81586 262658 81822 262894
rect 81266 262338 81502 262574
rect 81586 262338 81822 262574
rect 84986 374378 85222 374614
rect 85306 374378 85542 374614
rect 84986 374058 85222 374294
rect 85306 374058 85542 374294
rect 84986 338378 85222 338614
rect 85306 338378 85542 338614
rect 84986 338058 85222 338294
rect 85306 338058 85542 338294
rect 84986 302378 85222 302614
rect 85306 302378 85542 302614
rect 84986 302058 85222 302294
rect 85306 302058 85542 302294
rect 84986 266378 85222 266614
rect 85306 266378 85542 266614
rect 84986 266058 85222 266294
rect 85306 266058 85542 266294
rect 84986 230378 85222 230614
rect 85306 230378 85542 230614
rect 84986 230058 85222 230294
rect 85306 230058 85542 230294
rect 91826 381218 92062 381454
rect 92146 381218 92382 381454
rect 91826 380898 92062 381134
rect 92146 380898 92382 381134
rect 91826 345218 92062 345454
rect 92146 345218 92382 345454
rect 91826 344898 92062 345134
rect 92146 344898 92382 345134
rect 91826 309218 92062 309454
rect 92146 309218 92382 309454
rect 91826 308898 92062 309134
rect 92146 308898 92382 309134
rect 91826 273218 92062 273454
rect 92146 273218 92382 273454
rect 91826 272898 92062 273134
rect 92146 272898 92382 273134
rect 91826 237218 92062 237454
rect 92146 237218 92382 237454
rect 91826 236898 92062 237134
rect 92146 236898 92382 237134
rect 95546 384938 95782 385174
rect 95866 384938 96102 385174
rect 95546 384618 95782 384854
rect 95866 384618 96102 384854
rect 95546 348938 95782 349174
rect 95866 348938 96102 349174
rect 95546 348618 95782 348854
rect 95866 348618 96102 348854
rect 95546 312938 95782 313174
rect 95866 312938 96102 313174
rect 95546 312618 95782 312854
rect 95866 312618 96102 312854
rect 95546 276938 95782 277174
rect 95866 276938 96102 277174
rect 95546 276618 95782 276854
rect 95866 276618 96102 276854
rect 95546 240938 95782 241174
rect 95866 240938 96102 241174
rect 95546 240618 95782 240854
rect 95866 240618 96102 240854
rect 99266 388658 99502 388894
rect 99586 388658 99822 388894
rect 99266 388338 99502 388574
rect 99586 388338 99822 388574
rect 99266 352658 99502 352894
rect 99586 352658 99822 352894
rect 99266 352338 99502 352574
rect 99586 352338 99822 352574
rect 99266 316658 99502 316894
rect 99586 316658 99822 316894
rect 99266 316338 99502 316574
rect 99586 316338 99822 316574
rect 99266 280658 99502 280894
rect 99586 280658 99822 280894
rect 99266 280338 99502 280574
rect 99586 280338 99822 280574
rect 99266 244658 99502 244894
rect 99586 244658 99822 244894
rect 99266 244338 99502 244574
rect 99586 244338 99822 244574
rect 102986 392378 103222 392614
rect 103306 392378 103542 392614
rect 102986 392058 103222 392294
rect 103306 392058 103542 392294
rect 102986 356378 103222 356614
rect 103306 356378 103542 356614
rect 102986 356058 103222 356294
rect 103306 356058 103542 356294
rect 102986 320378 103222 320614
rect 103306 320378 103542 320614
rect 102986 320058 103222 320294
rect 103306 320058 103542 320294
rect 102986 284378 103222 284614
rect 103306 284378 103542 284614
rect 102986 284058 103222 284294
rect 103306 284058 103542 284294
rect 102986 248378 103222 248614
rect 103306 248378 103542 248614
rect 102986 248058 103222 248294
rect 103306 248058 103542 248294
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 109826 291218 110062 291454
rect 110146 291218 110382 291454
rect 109826 290898 110062 291134
rect 110146 290898 110382 291134
rect 109826 255218 110062 255454
rect 110146 255218 110382 255454
rect 109826 254898 110062 255134
rect 110146 254898 110382 255134
rect 113546 366938 113782 367174
rect 113866 366938 114102 367174
rect 113546 366618 113782 366854
rect 113866 366618 114102 366854
rect 113546 330938 113782 331174
rect 113866 330938 114102 331174
rect 113546 330618 113782 330854
rect 113866 330618 114102 330854
rect 113546 294938 113782 295174
rect 113866 294938 114102 295174
rect 113546 294618 113782 294854
rect 113866 294618 114102 294854
rect 113546 258938 113782 259174
rect 113866 258938 114102 259174
rect 113546 258618 113782 258854
rect 113866 258618 114102 258854
rect 117266 370658 117502 370894
rect 117586 370658 117822 370894
rect 117266 370338 117502 370574
rect 117586 370338 117822 370574
rect 117266 334658 117502 334894
rect 117586 334658 117822 334894
rect 117266 334338 117502 334574
rect 117586 334338 117822 334574
rect 117266 298658 117502 298894
rect 117586 298658 117822 298894
rect 117266 298338 117502 298574
rect 117586 298338 117822 298574
rect 117266 262658 117502 262894
rect 117586 262658 117822 262894
rect 117266 262338 117502 262574
rect 117586 262338 117822 262574
rect 120986 374378 121222 374614
rect 121306 374378 121542 374614
rect 120986 374058 121222 374294
rect 121306 374058 121542 374294
rect 120986 338378 121222 338614
rect 121306 338378 121542 338614
rect 120986 338058 121222 338294
rect 121306 338058 121542 338294
rect 120986 302378 121222 302614
rect 121306 302378 121542 302614
rect 120986 302058 121222 302294
rect 121306 302058 121542 302294
rect 120986 266378 121222 266614
rect 121306 266378 121542 266614
rect 120986 266058 121222 266294
rect 121306 266058 121542 266294
rect 120986 230378 121222 230614
rect 121306 230378 121542 230614
rect 120986 230058 121222 230294
rect 121306 230058 121542 230294
rect 127826 381218 128062 381454
rect 128146 381218 128382 381454
rect 127826 380898 128062 381134
rect 128146 380898 128382 381134
rect 127826 345218 128062 345454
rect 128146 345218 128382 345454
rect 127826 344898 128062 345134
rect 128146 344898 128382 345134
rect 127826 309218 128062 309454
rect 128146 309218 128382 309454
rect 127826 308898 128062 309134
rect 128146 308898 128382 309134
rect 127826 273218 128062 273454
rect 128146 273218 128382 273454
rect 127826 272898 128062 273134
rect 128146 272898 128382 273134
rect 127826 237218 128062 237454
rect 128146 237218 128382 237454
rect 127826 236898 128062 237134
rect 128146 236898 128382 237134
rect 131546 384938 131782 385174
rect 131866 384938 132102 385174
rect 131546 384618 131782 384854
rect 131866 384618 132102 384854
rect 131546 348938 131782 349174
rect 131866 348938 132102 349174
rect 131546 348618 131782 348854
rect 131866 348618 132102 348854
rect 131546 312938 131782 313174
rect 131866 312938 132102 313174
rect 131546 312618 131782 312854
rect 131866 312618 132102 312854
rect 131546 276938 131782 277174
rect 131866 276938 132102 277174
rect 131546 276618 131782 276854
rect 131866 276618 132102 276854
rect 131546 240938 131782 241174
rect 131866 240938 132102 241174
rect 131546 240618 131782 240854
rect 131866 240618 132102 240854
rect 135266 388658 135502 388894
rect 135586 388658 135822 388894
rect 135266 388338 135502 388574
rect 135586 388338 135822 388574
rect 135266 352658 135502 352894
rect 135586 352658 135822 352894
rect 135266 352338 135502 352574
rect 135586 352338 135822 352574
rect 135266 316658 135502 316894
rect 135586 316658 135822 316894
rect 135266 316338 135502 316574
rect 135586 316338 135822 316574
rect 135266 280658 135502 280894
rect 135586 280658 135822 280894
rect 135266 280338 135502 280574
rect 135586 280338 135822 280574
rect 135266 244658 135502 244894
rect 135586 244658 135822 244894
rect 135266 244338 135502 244574
rect 135586 244338 135822 244574
rect 138986 392378 139222 392614
rect 139306 392378 139542 392614
rect 138986 392058 139222 392294
rect 139306 392058 139542 392294
rect 138986 356378 139222 356614
rect 139306 356378 139542 356614
rect 138986 356058 139222 356294
rect 139306 356058 139542 356294
rect 138986 320378 139222 320614
rect 139306 320378 139542 320614
rect 138986 320058 139222 320294
rect 139306 320058 139542 320294
rect 138986 284378 139222 284614
rect 139306 284378 139542 284614
rect 138986 284058 139222 284294
rect 139306 284058 139542 284294
rect 138986 248378 139222 248614
rect 139306 248378 139542 248614
rect 138986 248058 139222 248294
rect 139306 248058 139542 248294
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 149546 366938 149782 367174
rect 149866 366938 150102 367174
rect 149546 366618 149782 366854
rect 149866 366618 150102 366854
rect 149546 330938 149782 331174
rect 149866 330938 150102 331174
rect 149546 330618 149782 330854
rect 149866 330618 150102 330854
rect 149546 294938 149782 295174
rect 149866 294938 150102 295174
rect 149546 294618 149782 294854
rect 149866 294618 150102 294854
rect 149546 258938 149782 259174
rect 149866 258938 150102 259174
rect 149546 258618 149782 258854
rect 149866 258618 150102 258854
rect 153266 370658 153502 370894
rect 153586 370658 153822 370894
rect 153266 370338 153502 370574
rect 153586 370338 153822 370574
rect 153266 334658 153502 334894
rect 153586 334658 153822 334894
rect 153266 334338 153502 334574
rect 153586 334338 153822 334574
rect 153266 298658 153502 298894
rect 153586 298658 153822 298894
rect 153266 298338 153502 298574
rect 153586 298338 153822 298574
rect 153266 262658 153502 262894
rect 153586 262658 153822 262894
rect 153266 262338 153502 262574
rect 153586 262338 153822 262574
rect 156986 374378 157222 374614
rect 157306 374378 157542 374614
rect 156986 374058 157222 374294
rect 157306 374058 157542 374294
rect 156986 338378 157222 338614
rect 157306 338378 157542 338614
rect 156986 338058 157222 338294
rect 157306 338058 157542 338294
rect 156986 302378 157222 302614
rect 157306 302378 157542 302614
rect 156986 302058 157222 302294
rect 157306 302058 157542 302294
rect 156986 266378 157222 266614
rect 157306 266378 157542 266614
rect 156986 266058 157222 266294
rect 157306 266058 157542 266294
rect 156986 230378 157222 230614
rect 157306 230378 157542 230614
rect 156986 230058 157222 230294
rect 157306 230058 157542 230294
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 163826 345218 164062 345454
rect 164146 345218 164382 345454
rect 163826 344898 164062 345134
rect 164146 344898 164382 345134
rect 163826 309218 164062 309454
rect 164146 309218 164382 309454
rect 163826 308898 164062 309134
rect 164146 308898 164382 309134
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 163826 237218 164062 237454
rect 164146 237218 164382 237454
rect 163826 236898 164062 237134
rect 164146 236898 164382 237134
rect 167546 384938 167782 385174
rect 167866 384938 168102 385174
rect 167546 384618 167782 384854
rect 167866 384618 168102 384854
rect 167546 348938 167782 349174
rect 167866 348938 168102 349174
rect 167546 348618 167782 348854
rect 167866 348618 168102 348854
rect 167546 312938 167782 313174
rect 167866 312938 168102 313174
rect 167546 312618 167782 312854
rect 167866 312618 168102 312854
rect 167546 276938 167782 277174
rect 167866 276938 168102 277174
rect 167546 276618 167782 276854
rect 167866 276618 168102 276854
rect 167546 240938 167782 241174
rect 167866 240938 168102 241174
rect 167546 240618 167782 240854
rect 167866 240618 168102 240854
rect 171266 388658 171502 388894
rect 171586 388658 171822 388894
rect 171266 388338 171502 388574
rect 171586 388338 171822 388574
rect 171266 352658 171502 352894
rect 171586 352658 171822 352894
rect 171266 352338 171502 352574
rect 171586 352338 171822 352574
rect 171266 316658 171502 316894
rect 171586 316658 171822 316894
rect 171266 316338 171502 316574
rect 171586 316338 171822 316574
rect 171266 280658 171502 280894
rect 171586 280658 171822 280894
rect 171266 280338 171502 280574
rect 171586 280338 171822 280574
rect 171266 244658 171502 244894
rect 171586 244658 171822 244894
rect 171266 244338 171502 244574
rect 171586 244338 171822 244574
rect 174986 392378 175222 392614
rect 175306 392378 175542 392614
rect 174986 392058 175222 392294
rect 175306 392058 175542 392294
rect 174986 356378 175222 356614
rect 175306 356378 175542 356614
rect 174986 356058 175222 356294
rect 175306 356058 175542 356294
rect 174986 320378 175222 320614
rect 175306 320378 175542 320614
rect 174986 320058 175222 320294
rect 175306 320058 175542 320294
rect 174986 284378 175222 284614
rect 175306 284378 175542 284614
rect 174986 284058 175222 284294
rect 175306 284058 175542 284294
rect 174986 248378 175222 248614
rect 175306 248378 175542 248614
rect 174986 248058 175222 248294
rect 175306 248058 175542 248294
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 185546 366938 185782 367174
rect 185866 366938 186102 367174
rect 185546 366618 185782 366854
rect 185866 366618 186102 366854
rect 185546 330938 185782 331174
rect 185866 330938 186102 331174
rect 185546 330618 185782 330854
rect 185866 330618 186102 330854
rect 185546 294938 185782 295174
rect 185866 294938 186102 295174
rect 185546 294618 185782 294854
rect 185866 294618 186102 294854
rect 185546 258938 185782 259174
rect 185866 258938 186102 259174
rect 185546 258618 185782 258854
rect 185866 258618 186102 258854
rect 189266 370658 189502 370894
rect 189586 370658 189822 370894
rect 189266 370338 189502 370574
rect 189586 370338 189822 370574
rect 189266 334658 189502 334894
rect 189586 334658 189822 334894
rect 189266 334338 189502 334574
rect 189586 334338 189822 334574
rect 189266 298658 189502 298894
rect 189586 298658 189822 298894
rect 189266 298338 189502 298574
rect 189586 298338 189822 298574
rect 189266 262658 189502 262894
rect 189586 262658 189822 262894
rect 189266 262338 189502 262574
rect 189586 262338 189822 262574
rect 192986 374378 193222 374614
rect 193306 374378 193542 374614
rect 192986 374058 193222 374294
rect 193306 374058 193542 374294
rect 192986 338378 193222 338614
rect 193306 338378 193542 338614
rect 192986 338058 193222 338294
rect 193306 338058 193542 338294
rect 192986 302378 193222 302614
rect 193306 302378 193542 302614
rect 192986 302058 193222 302294
rect 193306 302058 193542 302294
rect 192986 266378 193222 266614
rect 193306 266378 193542 266614
rect 192986 266058 193222 266294
rect 193306 266058 193542 266294
rect 192986 230378 193222 230614
rect 193306 230378 193542 230614
rect 192986 230058 193222 230294
rect 193306 230058 193542 230294
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 199826 345218 200062 345454
rect 200146 345218 200382 345454
rect 199826 344898 200062 345134
rect 200146 344898 200382 345134
rect 199826 309218 200062 309454
rect 200146 309218 200382 309454
rect 199826 308898 200062 309134
rect 200146 308898 200382 309134
rect 199826 273218 200062 273454
rect 200146 273218 200382 273454
rect 199826 272898 200062 273134
rect 200146 272898 200382 273134
rect 199826 237218 200062 237454
rect 200146 237218 200382 237454
rect 199826 236898 200062 237134
rect 200146 236898 200382 237134
rect 203546 672938 203782 673174
rect 203866 672938 204102 673174
rect 203546 672618 203782 672854
rect 203866 672618 204102 672854
rect 203546 636938 203782 637174
rect 203866 636938 204102 637174
rect 203546 636618 203782 636854
rect 203866 636618 204102 636854
rect 203546 600938 203782 601174
rect 203866 600938 204102 601174
rect 203546 600618 203782 600854
rect 203866 600618 204102 600854
rect 203546 564938 203782 565174
rect 203866 564938 204102 565174
rect 203546 564618 203782 564854
rect 203866 564618 204102 564854
rect 203546 528938 203782 529174
rect 203866 528938 204102 529174
rect 203546 528618 203782 528854
rect 203866 528618 204102 528854
rect 203546 492938 203782 493174
rect 203866 492938 204102 493174
rect 203546 492618 203782 492854
rect 203866 492618 204102 492854
rect 203546 456938 203782 457174
rect 203866 456938 204102 457174
rect 203546 456618 203782 456854
rect 203866 456618 204102 456854
rect 203546 420938 203782 421174
rect 203866 420938 204102 421174
rect 203546 420618 203782 420854
rect 203866 420618 204102 420854
rect 203546 384938 203782 385174
rect 203866 384938 204102 385174
rect 203546 384618 203782 384854
rect 203866 384618 204102 384854
rect 203546 348938 203782 349174
rect 203866 348938 204102 349174
rect 203546 348618 203782 348854
rect 203866 348618 204102 348854
rect 203546 312938 203782 313174
rect 203866 312938 204102 313174
rect 203546 312618 203782 312854
rect 203866 312618 204102 312854
rect 203546 276938 203782 277174
rect 203866 276938 204102 277174
rect 203546 276618 203782 276854
rect 203866 276618 204102 276854
rect 203546 240938 203782 241174
rect 203866 240938 204102 241174
rect 203546 240618 203782 240854
rect 203866 240618 204102 240854
rect 207266 676658 207502 676894
rect 207586 676658 207822 676894
rect 207266 676338 207502 676574
rect 207586 676338 207822 676574
rect 207266 640658 207502 640894
rect 207586 640658 207822 640894
rect 207266 640338 207502 640574
rect 207586 640338 207822 640574
rect 207266 604658 207502 604894
rect 207586 604658 207822 604894
rect 207266 604338 207502 604574
rect 207586 604338 207822 604574
rect 207266 568658 207502 568894
rect 207586 568658 207822 568894
rect 207266 568338 207502 568574
rect 207586 568338 207822 568574
rect 207266 532658 207502 532894
rect 207586 532658 207822 532894
rect 207266 532338 207502 532574
rect 207586 532338 207822 532574
rect 207266 496658 207502 496894
rect 207586 496658 207822 496894
rect 207266 496338 207502 496574
rect 207586 496338 207822 496574
rect 207266 460658 207502 460894
rect 207586 460658 207822 460894
rect 207266 460338 207502 460574
rect 207586 460338 207822 460574
rect 207266 424658 207502 424894
rect 207586 424658 207822 424894
rect 207266 424338 207502 424574
rect 207586 424338 207822 424574
rect 207266 388658 207502 388894
rect 207586 388658 207822 388894
rect 207266 388338 207502 388574
rect 207586 388338 207822 388574
rect 207266 352658 207502 352894
rect 207586 352658 207822 352894
rect 207266 352338 207502 352574
rect 207586 352338 207822 352574
rect 207266 316658 207502 316894
rect 207586 316658 207822 316894
rect 207266 316338 207502 316574
rect 207586 316338 207822 316574
rect 207266 280658 207502 280894
rect 207586 280658 207822 280894
rect 207266 280338 207502 280574
rect 207586 280338 207822 280574
rect 207266 244658 207502 244894
rect 207586 244658 207822 244894
rect 207266 244338 207502 244574
rect 207586 244338 207822 244574
rect 228986 710362 229222 710598
rect 229306 710362 229542 710598
rect 228986 710042 229222 710278
rect 229306 710042 229542 710278
rect 225266 708442 225502 708678
rect 225586 708442 225822 708678
rect 225266 708122 225502 708358
rect 225586 708122 225822 708358
rect 221546 706522 221782 706758
rect 221866 706522 222102 706758
rect 221546 706202 221782 706438
rect 221866 706202 222102 706438
rect 210986 680378 211222 680614
rect 211306 680378 211542 680614
rect 210986 680058 211222 680294
rect 211306 680058 211542 680294
rect 210986 644378 211222 644614
rect 211306 644378 211542 644614
rect 210986 644058 211222 644294
rect 211306 644058 211542 644294
rect 210986 608378 211222 608614
rect 211306 608378 211542 608614
rect 210986 608058 211222 608294
rect 211306 608058 211542 608294
rect 210986 572378 211222 572614
rect 211306 572378 211542 572614
rect 210986 572058 211222 572294
rect 211306 572058 211542 572294
rect 210986 536378 211222 536614
rect 211306 536378 211542 536614
rect 210986 536058 211222 536294
rect 211306 536058 211542 536294
rect 210986 500378 211222 500614
rect 211306 500378 211542 500614
rect 210986 500058 211222 500294
rect 211306 500058 211542 500294
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 221546 654938 221782 655174
rect 221866 654938 222102 655174
rect 221546 654618 221782 654854
rect 221866 654618 222102 654854
rect 221546 618938 221782 619174
rect 221866 618938 222102 619174
rect 221546 618618 221782 618854
rect 221866 618618 222102 618854
rect 221546 582938 221782 583174
rect 221866 582938 222102 583174
rect 221546 582618 221782 582854
rect 221866 582618 222102 582854
rect 221546 546938 221782 547174
rect 221866 546938 222102 547174
rect 221546 546618 221782 546854
rect 221866 546618 222102 546854
rect 221546 510938 221782 511174
rect 221866 510938 222102 511174
rect 221546 510618 221782 510854
rect 221866 510618 222102 510854
rect 210986 464378 211222 464614
rect 211306 464378 211542 464614
rect 210986 464058 211222 464294
rect 211306 464058 211542 464294
rect 210986 428378 211222 428614
rect 211306 428378 211542 428614
rect 210986 428058 211222 428294
rect 211306 428058 211542 428294
rect 210986 392378 211222 392614
rect 211306 392378 211542 392614
rect 210986 392058 211222 392294
rect 211306 392058 211542 392294
rect 210986 356378 211222 356614
rect 211306 356378 211542 356614
rect 210986 356058 211222 356294
rect 211306 356058 211542 356294
rect 210986 320378 211222 320614
rect 211306 320378 211542 320614
rect 210986 320058 211222 320294
rect 211306 320058 211542 320294
rect 210986 284378 211222 284614
rect 211306 284378 211542 284614
rect 210986 284058 211222 284294
rect 211306 284058 211542 284294
rect 210986 248378 211222 248614
rect 211306 248378 211542 248614
rect 210986 248058 211222 248294
rect 211306 248058 211542 248294
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 217826 291218 218062 291454
rect 218146 291218 218382 291454
rect 217826 290898 218062 291134
rect 218146 290898 218382 291134
rect 217826 255218 218062 255454
rect 218146 255218 218382 255454
rect 217826 254898 218062 255134
rect 218146 254898 218382 255134
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 225266 658658 225502 658894
rect 225586 658658 225822 658894
rect 225266 658338 225502 658574
rect 225586 658338 225822 658574
rect 225266 622658 225502 622894
rect 225586 622658 225822 622894
rect 225266 622338 225502 622574
rect 225586 622338 225822 622574
rect 225266 586658 225502 586894
rect 225586 586658 225822 586894
rect 225266 586338 225502 586574
rect 225586 586338 225822 586574
rect 225266 550658 225502 550894
rect 225586 550658 225822 550894
rect 225266 550338 225502 550574
rect 225586 550338 225822 550574
rect 225266 514658 225502 514894
rect 225586 514658 225822 514894
rect 225266 514338 225502 514574
rect 225586 514338 225822 514574
rect 246986 711322 247222 711558
rect 247306 711322 247542 711558
rect 246986 711002 247222 711238
rect 247306 711002 247542 711238
rect 243266 709402 243502 709638
rect 243586 709402 243822 709638
rect 243266 709082 243502 709318
rect 243586 709082 243822 709318
rect 239546 707482 239782 707718
rect 239866 707482 240102 707718
rect 239546 707162 239782 707398
rect 239866 707162 240102 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 228986 662378 229222 662614
rect 229306 662378 229542 662614
rect 228986 662058 229222 662294
rect 229306 662058 229542 662294
rect 228986 626378 229222 626614
rect 229306 626378 229542 626614
rect 228986 626058 229222 626294
rect 229306 626058 229542 626294
rect 228986 590378 229222 590614
rect 229306 590378 229542 590614
rect 228986 590058 229222 590294
rect 229306 590058 229542 590294
rect 228986 554378 229222 554614
rect 229306 554378 229542 554614
rect 228986 554058 229222 554294
rect 229306 554058 229542 554294
rect 228986 518378 229222 518614
rect 229306 518378 229542 518614
rect 228986 518058 229222 518294
rect 229306 518058 229542 518294
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 235826 525218 236062 525454
rect 236146 525218 236382 525454
rect 235826 524898 236062 525134
rect 236146 524898 236382 525134
rect 235826 489218 236062 489454
rect 236146 489218 236382 489454
rect 235826 488898 236062 489134
rect 236146 488898 236382 489134
rect 239546 672938 239782 673174
rect 239866 672938 240102 673174
rect 239546 672618 239782 672854
rect 239866 672618 240102 672854
rect 239546 636938 239782 637174
rect 239866 636938 240102 637174
rect 239546 636618 239782 636854
rect 239866 636618 240102 636854
rect 239546 600938 239782 601174
rect 239866 600938 240102 601174
rect 239546 600618 239782 600854
rect 239866 600618 240102 600854
rect 239546 564938 239782 565174
rect 239866 564938 240102 565174
rect 239546 564618 239782 564854
rect 239866 564618 240102 564854
rect 239546 528938 239782 529174
rect 239866 528938 240102 529174
rect 239546 528618 239782 528854
rect 239866 528618 240102 528854
rect 239546 492938 239782 493174
rect 239866 492938 240102 493174
rect 239546 492618 239782 492854
rect 239866 492618 240102 492854
rect 243266 676658 243502 676894
rect 243586 676658 243822 676894
rect 243266 676338 243502 676574
rect 243586 676338 243822 676574
rect 243266 640658 243502 640894
rect 243586 640658 243822 640894
rect 243266 640338 243502 640574
rect 243586 640338 243822 640574
rect 243266 604658 243502 604894
rect 243586 604658 243822 604894
rect 243266 604338 243502 604574
rect 243586 604338 243822 604574
rect 243266 568658 243502 568894
rect 243586 568658 243822 568894
rect 243266 568338 243502 568574
rect 243586 568338 243822 568574
rect 243266 532658 243502 532894
rect 243586 532658 243822 532894
rect 243266 532338 243502 532574
rect 243586 532338 243822 532574
rect 243266 496658 243502 496894
rect 243586 496658 243822 496894
rect 243266 496338 243502 496574
rect 243586 496338 243822 496574
rect 264986 710362 265222 710598
rect 265306 710362 265542 710598
rect 264986 710042 265222 710278
rect 265306 710042 265542 710278
rect 261266 708442 261502 708678
rect 261586 708442 261822 708678
rect 261266 708122 261502 708358
rect 261586 708122 261822 708358
rect 257546 706522 257782 706758
rect 257866 706522 258102 706758
rect 257546 706202 257782 706438
rect 257866 706202 258102 706438
rect 246986 680378 247222 680614
rect 247306 680378 247542 680614
rect 246986 680058 247222 680294
rect 247306 680058 247542 680294
rect 246986 644378 247222 644614
rect 247306 644378 247542 644614
rect 246986 644058 247222 644294
rect 247306 644058 247542 644294
rect 246986 608378 247222 608614
rect 247306 608378 247542 608614
rect 246986 608058 247222 608294
rect 247306 608058 247542 608294
rect 246986 572378 247222 572614
rect 247306 572378 247542 572614
rect 246986 572058 247222 572294
rect 247306 572058 247542 572294
rect 246986 536378 247222 536614
rect 247306 536378 247542 536614
rect 246986 536058 247222 536294
rect 247306 536058 247542 536294
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 246986 500378 247222 500614
rect 247306 500378 247542 500614
rect 246986 500058 247222 500294
rect 247306 500058 247542 500294
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 257546 654938 257782 655174
rect 257866 654938 258102 655174
rect 257546 654618 257782 654854
rect 257866 654618 258102 654854
rect 257546 618938 257782 619174
rect 257866 618938 258102 619174
rect 257546 618618 257782 618854
rect 257866 618618 258102 618854
rect 257546 582938 257782 583174
rect 257866 582938 258102 583174
rect 257546 582618 257782 582854
rect 257866 582618 258102 582854
rect 257546 546938 257782 547174
rect 257866 546938 258102 547174
rect 257546 546618 257782 546854
rect 257866 546618 258102 546854
rect 257546 510938 257782 511174
rect 257866 510938 258102 511174
rect 257546 510618 257782 510854
rect 257866 510618 258102 510854
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 261266 658658 261502 658894
rect 261586 658658 261822 658894
rect 261266 658338 261502 658574
rect 261586 658338 261822 658574
rect 261266 622658 261502 622894
rect 261586 622658 261822 622894
rect 261266 622338 261502 622574
rect 261586 622338 261822 622574
rect 261266 586658 261502 586894
rect 261586 586658 261822 586894
rect 261266 586338 261502 586574
rect 261586 586338 261822 586574
rect 261266 550658 261502 550894
rect 261586 550658 261822 550894
rect 261266 550338 261502 550574
rect 261586 550338 261822 550574
rect 261266 514658 261502 514894
rect 261586 514658 261822 514894
rect 261266 514338 261502 514574
rect 261586 514338 261822 514574
rect 282986 711322 283222 711558
rect 283306 711322 283542 711558
rect 282986 711002 283222 711238
rect 283306 711002 283542 711238
rect 279266 709402 279502 709638
rect 279586 709402 279822 709638
rect 279266 709082 279502 709318
rect 279586 709082 279822 709318
rect 275546 707482 275782 707718
rect 275866 707482 276102 707718
rect 275546 707162 275782 707398
rect 275866 707162 276102 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 264986 662378 265222 662614
rect 265306 662378 265542 662614
rect 264986 662058 265222 662294
rect 265306 662058 265542 662294
rect 264986 626378 265222 626614
rect 265306 626378 265542 626614
rect 264986 626058 265222 626294
rect 265306 626058 265542 626294
rect 264986 590378 265222 590614
rect 265306 590378 265542 590614
rect 264986 590058 265222 590294
rect 265306 590058 265542 590294
rect 264986 554378 265222 554614
rect 265306 554378 265542 554614
rect 264986 554058 265222 554294
rect 265306 554058 265542 554294
rect 264986 518378 265222 518614
rect 265306 518378 265542 518614
rect 264986 518058 265222 518294
rect 265306 518058 265542 518294
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 271826 525218 272062 525454
rect 272146 525218 272382 525454
rect 271826 524898 272062 525134
rect 272146 524898 272382 525134
rect 275546 672938 275782 673174
rect 275866 672938 276102 673174
rect 275546 672618 275782 672854
rect 275866 672618 276102 672854
rect 275546 636938 275782 637174
rect 275866 636938 276102 637174
rect 275546 636618 275782 636854
rect 275866 636618 276102 636854
rect 275546 600938 275782 601174
rect 275866 600938 276102 601174
rect 275546 600618 275782 600854
rect 275866 600618 276102 600854
rect 275546 564938 275782 565174
rect 275866 564938 276102 565174
rect 275546 564618 275782 564854
rect 275866 564618 276102 564854
rect 275546 528938 275782 529174
rect 275866 528938 276102 529174
rect 275546 528618 275782 528854
rect 275866 528618 276102 528854
rect 271826 489218 272062 489454
rect 272146 489218 272382 489454
rect 271826 488898 272062 489134
rect 272146 488898 272382 489134
rect 279266 676658 279502 676894
rect 279586 676658 279822 676894
rect 279266 676338 279502 676574
rect 279586 676338 279822 676574
rect 279266 640658 279502 640894
rect 279586 640658 279822 640894
rect 279266 640338 279502 640574
rect 279586 640338 279822 640574
rect 279266 604658 279502 604894
rect 279586 604658 279822 604894
rect 279266 604338 279502 604574
rect 279586 604338 279822 604574
rect 279266 568658 279502 568894
rect 279586 568658 279822 568894
rect 279266 568338 279502 568574
rect 279586 568338 279822 568574
rect 279266 532658 279502 532894
rect 279586 532658 279822 532894
rect 279266 532338 279502 532574
rect 279586 532338 279822 532574
rect 275546 492938 275782 493174
rect 275866 492938 276102 493174
rect 275546 492618 275782 492854
rect 275866 492618 276102 492854
rect 300986 710362 301222 710598
rect 301306 710362 301542 710598
rect 300986 710042 301222 710278
rect 301306 710042 301542 710278
rect 297266 708442 297502 708678
rect 297586 708442 297822 708678
rect 297266 708122 297502 708358
rect 297586 708122 297822 708358
rect 293546 706522 293782 706758
rect 293866 706522 294102 706758
rect 293546 706202 293782 706438
rect 293866 706202 294102 706438
rect 282986 680378 283222 680614
rect 283306 680378 283542 680614
rect 282986 680058 283222 680294
rect 283306 680058 283542 680294
rect 282986 644378 283222 644614
rect 283306 644378 283542 644614
rect 282986 644058 283222 644294
rect 283306 644058 283542 644294
rect 282986 608378 283222 608614
rect 283306 608378 283542 608614
rect 282986 608058 283222 608294
rect 283306 608058 283542 608294
rect 282986 572378 283222 572614
rect 283306 572378 283542 572614
rect 282986 572058 283222 572294
rect 283306 572058 283542 572294
rect 282986 536378 283222 536614
rect 283306 536378 283542 536614
rect 282986 536058 283222 536294
rect 283306 536058 283542 536294
rect 279266 496658 279502 496894
rect 279586 496658 279822 496894
rect 279266 496338 279502 496574
rect 279586 496338 279822 496574
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 282986 500378 283222 500614
rect 283306 500378 283542 500614
rect 282986 500058 283222 500294
rect 283306 500058 283542 500294
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 293546 654938 293782 655174
rect 293866 654938 294102 655174
rect 293546 654618 293782 654854
rect 293866 654618 294102 654854
rect 293546 618938 293782 619174
rect 293866 618938 294102 619174
rect 293546 618618 293782 618854
rect 293866 618618 294102 618854
rect 293546 582938 293782 583174
rect 293866 582938 294102 583174
rect 293546 582618 293782 582854
rect 293866 582618 294102 582854
rect 293546 546938 293782 547174
rect 293866 546938 294102 547174
rect 293546 546618 293782 546854
rect 293866 546618 294102 546854
rect 293546 510938 293782 511174
rect 293866 510938 294102 511174
rect 293546 510618 293782 510854
rect 293866 510618 294102 510854
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 297266 658658 297502 658894
rect 297586 658658 297822 658894
rect 297266 658338 297502 658574
rect 297586 658338 297822 658574
rect 297266 622658 297502 622894
rect 297586 622658 297822 622894
rect 297266 622338 297502 622574
rect 297586 622338 297822 622574
rect 297266 586658 297502 586894
rect 297586 586658 297822 586894
rect 297266 586338 297502 586574
rect 297586 586338 297822 586574
rect 297266 550658 297502 550894
rect 297586 550658 297822 550894
rect 297266 550338 297502 550574
rect 297586 550338 297822 550574
rect 297266 514658 297502 514894
rect 297586 514658 297822 514894
rect 297266 514338 297502 514574
rect 297586 514338 297822 514574
rect 318986 711322 319222 711558
rect 319306 711322 319542 711558
rect 318986 711002 319222 711238
rect 319306 711002 319542 711238
rect 315266 709402 315502 709638
rect 315586 709402 315822 709638
rect 315266 709082 315502 709318
rect 315586 709082 315822 709318
rect 311546 707482 311782 707718
rect 311866 707482 312102 707718
rect 311546 707162 311782 707398
rect 311866 707162 312102 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 300986 662378 301222 662614
rect 301306 662378 301542 662614
rect 300986 662058 301222 662294
rect 301306 662058 301542 662294
rect 300986 626378 301222 626614
rect 301306 626378 301542 626614
rect 300986 626058 301222 626294
rect 301306 626058 301542 626294
rect 300986 590378 301222 590614
rect 301306 590378 301542 590614
rect 300986 590058 301222 590294
rect 301306 590058 301542 590294
rect 300986 554378 301222 554614
rect 301306 554378 301542 554614
rect 300986 554058 301222 554294
rect 301306 554058 301542 554294
rect 300986 518378 301222 518614
rect 301306 518378 301542 518614
rect 300986 518058 301222 518294
rect 301306 518058 301542 518294
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 311546 672938 311782 673174
rect 311866 672938 312102 673174
rect 311546 672618 311782 672854
rect 311866 672618 312102 672854
rect 311546 636938 311782 637174
rect 311866 636938 312102 637174
rect 311546 636618 311782 636854
rect 311866 636618 312102 636854
rect 311546 600938 311782 601174
rect 311866 600938 312102 601174
rect 311546 600618 311782 600854
rect 311866 600618 312102 600854
rect 311546 564938 311782 565174
rect 311866 564938 312102 565174
rect 311546 564618 311782 564854
rect 311866 564618 312102 564854
rect 311546 528938 311782 529174
rect 311866 528938 312102 529174
rect 311546 528618 311782 528854
rect 311866 528618 312102 528854
rect 311546 492938 311782 493174
rect 311866 492938 312102 493174
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 311546 492618 311782 492854
rect 311866 492618 312102 492854
rect 315266 676658 315502 676894
rect 315586 676658 315822 676894
rect 315266 676338 315502 676574
rect 315586 676338 315822 676574
rect 315266 640658 315502 640894
rect 315586 640658 315822 640894
rect 315266 640338 315502 640574
rect 315586 640338 315822 640574
rect 315266 604658 315502 604894
rect 315586 604658 315822 604894
rect 315266 604338 315502 604574
rect 315586 604338 315822 604574
rect 315266 568658 315502 568894
rect 315586 568658 315822 568894
rect 315266 568338 315502 568574
rect 315586 568338 315822 568574
rect 315266 532658 315502 532894
rect 315586 532658 315822 532894
rect 315266 532338 315502 532574
rect 315586 532338 315822 532574
rect 315266 496658 315502 496894
rect 315586 496658 315822 496894
rect 315266 496338 315502 496574
rect 315586 496338 315822 496574
rect 336986 710362 337222 710598
rect 337306 710362 337542 710598
rect 336986 710042 337222 710278
rect 337306 710042 337542 710278
rect 333266 708442 333502 708678
rect 333586 708442 333822 708678
rect 333266 708122 333502 708358
rect 333586 708122 333822 708358
rect 329546 706522 329782 706758
rect 329866 706522 330102 706758
rect 329546 706202 329782 706438
rect 329866 706202 330102 706438
rect 318986 680378 319222 680614
rect 319306 680378 319542 680614
rect 318986 680058 319222 680294
rect 319306 680058 319542 680294
rect 318986 644378 319222 644614
rect 319306 644378 319542 644614
rect 318986 644058 319222 644294
rect 319306 644058 319542 644294
rect 318986 608378 319222 608614
rect 319306 608378 319542 608614
rect 318986 608058 319222 608294
rect 319306 608058 319542 608294
rect 318986 572378 319222 572614
rect 319306 572378 319542 572614
rect 318986 572058 319222 572294
rect 319306 572058 319542 572294
rect 318986 536378 319222 536614
rect 319306 536378 319542 536614
rect 318986 536058 319222 536294
rect 319306 536058 319542 536294
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 318986 500378 319222 500614
rect 319306 500378 319542 500614
rect 318986 500058 319222 500294
rect 319306 500058 319542 500294
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 329546 654938 329782 655174
rect 329866 654938 330102 655174
rect 329546 654618 329782 654854
rect 329866 654618 330102 654854
rect 329546 618938 329782 619174
rect 329866 618938 330102 619174
rect 329546 618618 329782 618854
rect 329866 618618 330102 618854
rect 329546 582938 329782 583174
rect 329866 582938 330102 583174
rect 329546 582618 329782 582854
rect 329866 582618 330102 582854
rect 329546 546938 329782 547174
rect 329866 546938 330102 547174
rect 329546 546618 329782 546854
rect 329866 546618 330102 546854
rect 329546 510938 329782 511174
rect 329866 510938 330102 511174
rect 329546 510618 329782 510854
rect 329866 510618 330102 510854
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 333266 658658 333502 658894
rect 333586 658658 333822 658894
rect 333266 658338 333502 658574
rect 333586 658338 333822 658574
rect 333266 622658 333502 622894
rect 333586 622658 333822 622894
rect 333266 622338 333502 622574
rect 333586 622338 333822 622574
rect 333266 586658 333502 586894
rect 333586 586658 333822 586894
rect 333266 586338 333502 586574
rect 333586 586338 333822 586574
rect 333266 550658 333502 550894
rect 333586 550658 333822 550894
rect 333266 550338 333502 550574
rect 333586 550338 333822 550574
rect 333266 514658 333502 514894
rect 333586 514658 333822 514894
rect 333266 514338 333502 514574
rect 333586 514338 333822 514574
rect 354986 711322 355222 711558
rect 355306 711322 355542 711558
rect 354986 711002 355222 711238
rect 355306 711002 355542 711238
rect 351266 709402 351502 709638
rect 351586 709402 351822 709638
rect 351266 709082 351502 709318
rect 351586 709082 351822 709318
rect 347546 707482 347782 707718
rect 347866 707482 348102 707718
rect 347546 707162 347782 707398
rect 347866 707162 348102 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 336986 662378 337222 662614
rect 337306 662378 337542 662614
rect 336986 662058 337222 662294
rect 337306 662058 337542 662294
rect 336986 626378 337222 626614
rect 337306 626378 337542 626614
rect 336986 626058 337222 626294
rect 337306 626058 337542 626294
rect 336986 590378 337222 590614
rect 337306 590378 337542 590614
rect 336986 590058 337222 590294
rect 337306 590058 337542 590294
rect 336986 554378 337222 554614
rect 337306 554378 337542 554614
rect 336986 554058 337222 554294
rect 337306 554058 337542 554294
rect 336986 518378 337222 518614
rect 337306 518378 337542 518614
rect 336986 518058 337222 518294
rect 337306 518058 337542 518294
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 347546 672938 347782 673174
rect 347866 672938 348102 673174
rect 347546 672618 347782 672854
rect 347866 672618 348102 672854
rect 347546 636938 347782 637174
rect 347866 636938 348102 637174
rect 347546 636618 347782 636854
rect 347866 636618 348102 636854
rect 347546 600938 347782 601174
rect 347866 600938 348102 601174
rect 347546 600618 347782 600854
rect 347866 600618 348102 600854
rect 347546 564938 347782 565174
rect 347866 564938 348102 565174
rect 347546 564618 347782 564854
rect 347866 564618 348102 564854
rect 347546 528938 347782 529174
rect 347866 528938 348102 529174
rect 347546 528618 347782 528854
rect 347866 528618 348102 528854
rect 347546 492938 347782 493174
rect 347866 492938 348102 493174
rect 347546 492618 347782 492854
rect 347866 492618 348102 492854
rect 351266 676658 351502 676894
rect 351586 676658 351822 676894
rect 351266 676338 351502 676574
rect 351586 676338 351822 676574
rect 351266 640658 351502 640894
rect 351586 640658 351822 640894
rect 351266 640338 351502 640574
rect 351586 640338 351822 640574
rect 351266 604658 351502 604894
rect 351586 604658 351822 604894
rect 351266 604338 351502 604574
rect 351586 604338 351822 604574
rect 351266 568658 351502 568894
rect 351586 568658 351822 568894
rect 351266 568338 351502 568574
rect 351586 568338 351822 568574
rect 351266 532658 351502 532894
rect 351586 532658 351822 532894
rect 351266 532338 351502 532574
rect 351586 532338 351822 532574
rect 351266 496658 351502 496894
rect 351586 496658 351822 496894
rect 351266 496338 351502 496574
rect 351586 496338 351822 496574
rect 372986 710362 373222 710598
rect 373306 710362 373542 710598
rect 372986 710042 373222 710278
rect 373306 710042 373542 710278
rect 369266 708442 369502 708678
rect 369586 708442 369822 708678
rect 369266 708122 369502 708358
rect 369586 708122 369822 708358
rect 365546 706522 365782 706758
rect 365866 706522 366102 706758
rect 365546 706202 365782 706438
rect 365866 706202 366102 706438
rect 354986 680378 355222 680614
rect 355306 680378 355542 680614
rect 354986 680058 355222 680294
rect 355306 680058 355542 680294
rect 354986 644378 355222 644614
rect 355306 644378 355542 644614
rect 354986 644058 355222 644294
rect 355306 644058 355542 644294
rect 354986 608378 355222 608614
rect 355306 608378 355542 608614
rect 354986 608058 355222 608294
rect 355306 608058 355542 608294
rect 354986 572378 355222 572614
rect 355306 572378 355542 572614
rect 354986 572058 355222 572294
rect 355306 572058 355542 572294
rect 354986 536378 355222 536614
rect 355306 536378 355542 536614
rect 354986 536058 355222 536294
rect 355306 536058 355542 536294
rect 354986 500378 355222 500614
rect 355306 500378 355542 500614
rect 354986 500058 355222 500294
rect 355306 500058 355542 500294
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 221008 471218 221244 471454
rect 221008 470898 221244 471134
rect 355376 471218 355612 471454
rect 355376 470898 355612 471134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 220328 453218 220564 453454
rect 220328 452898 220564 453134
rect 356056 453218 356292 453454
rect 356056 452898 356292 453134
rect 221008 435218 221244 435454
rect 221008 434898 221244 435134
rect 355376 435218 355612 435454
rect 355376 434898 355612 435134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 220328 417218 220564 417454
rect 220328 416898 220564 417134
rect 356056 417218 356292 417454
rect 356056 416898 356292 417134
rect 221546 366938 221782 367174
rect 221866 366938 222102 367174
rect 221546 366618 221782 366854
rect 221866 366618 222102 366854
rect 221546 330938 221782 331174
rect 221866 330938 222102 331174
rect 221546 330618 221782 330854
rect 221866 330618 222102 330854
rect 221546 294938 221782 295174
rect 221866 294938 222102 295174
rect 221546 294618 221782 294854
rect 221866 294618 222102 294854
rect 221546 258938 221782 259174
rect 221866 258938 222102 259174
rect 221546 258618 221782 258854
rect 221866 258618 222102 258854
rect 225266 370658 225502 370894
rect 225586 370658 225822 370894
rect 225266 370338 225502 370574
rect 225586 370338 225822 370574
rect 225266 334658 225502 334894
rect 225586 334658 225822 334894
rect 225266 334338 225502 334574
rect 225586 334338 225822 334574
rect 225266 298658 225502 298894
rect 225586 298658 225822 298894
rect 225266 298338 225502 298574
rect 225586 298338 225822 298574
rect 225266 262658 225502 262894
rect 225586 262658 225822 262894
rect 225266 262338 225502 262574
rect 225586 262338 225822 262574
rect 64250 219218 64486 219454
rect 64250 218898 64486 219134
rect 94970 219218 95206 219454
rect 94970 218898 95206 219134
rect 125690 219218 125926 219454
rect 125690 218898 125926 219134
rect 156410 219218 156646 219454
rect 156410 218898 156646 219134
rect 187130 219218 187366 219454
rect 187130 218898 187366 219134
rect 217850 219218 218086 219454
rect 217850 218898 218086 219134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 79610 201218 79846 201454
rect 79610 200898 79846 201134
rect 110330 201218 110566 201454
rect 110330 200898 110566 201134
rect 141050 201218 141286 201454
rect 141050 200898 141286 201134
rect 171770 201218 172006 201454
rect 171770 200898 172006 201134
rect 202490 201218 202726 201454
rect 202490 200898 202726 201134
rect 64250 183218 64486 183454
rect 64250 182898 64486 183134
rect 94970 183218 95206 183454
rect 94970 182898 95206 183134
rect 125690 183218 125926 183454
rect 125690 182898 125926 183134
rect 156410 183218 156646 183454
rect 156410 182898 156646 183134
rect 187130 183218 187366 183454
rect 187130 182898 187366 183134
rect 217850 183218 218086 183454
rect 217850 182898 218086 183134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 79610 165218 79846 165454
rect 79610 164898 79846 165134
rect 110330 165218 110566 165454
rect 110330 164898 110566 165134
rect 141050 165218 141286 165454
rect 141050 164898 141286 165134
rect 171770 165218 172006 165454
rect 171770 164898 172006 165134
rect 202490 165218 202726 165454
rect 202490 164898 202726 165134
rect 64250 147218 64486 147454
rect 64250 146898 64486 147134
rect 94970 147218 95206 147454
rect 94970 146898 95206 147134
rect 125690 147218 125926 147454
rect 125690 146898 125926 147134
rect 156410 147218 156646 147454
rect 156410 146898 156646 147134
rect 187130 147218 187366 147454
rect 187130 146898 187366 147134
rect 217850 147218 218086 147454
rect 217850 146898 218086 147134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 79610 129218 79846 129454
rect 79610 128898 79846 129134
rect 110330 129218 110566 129454
rect 110330 128898 110566 129134
rect 141050 129218 141286 129454
rect 141050 128898 141286 129134
rect 171770 129218 172006 129454
rect 171770 128898 172006 129134
rect 202490 129218 202726 129454
rect 202490 128898 202726 129134
rect 64250 111218 64486 111454
rect 64250 110898 64486 111134
rect 94970 111218 95206 111454
rect 94970 110898 95206 111134
rect 125690 111218 125926 111454
rect 125690 110898 125926 111134
rect 156410 111218 156646 111454
rect 156410 110898 156646 111134
rect 187130 111218 187366 111454
rect 187130 110898 187366 111134
rect 217850 111218 218086 111454
rect 217850 110898 218086 111134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 79610 93218 79846 93454
rect 79610 92898 79846 93134
rect 110330 93218 110566 93454
rect 110330 92898 110566 93134
rect 141050 93218 141286 93454
rect 141050 92898 141286 93134
rect 171770 93218 172006 93454
rect 171770 92898 172006 93134
rect 202490 93218 202726 93454
rect 202490 92898 202726 93134
rect 64250 75218 64486 75454
rect 64250 74898 64486 75134
rect 94970 75218 95206 75454
rect 94970 74898 95206 75134
rect 125690 75218 125926 75454
rect 125690 74898 125926 75134
rect 156410 75218 156646 75454
rect 156410 74898 156646 75134
rect 187130 75218 187366 75454
rect 187130 74898 187366 75134
rect 217850 75218 218086 75454
rect 217850 74898 218086 75134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -1542 56062 -1306
rect 56146 -1542 56382 -1306
rect 55826 -1862 56062 -1626
rect 56146 -1862 56382 -1626
rect 59546 24938 59782 25174
rect 59866 24938 60102 25174
rect 59546 24618 59782 24854
rect 59866 24618 60102 24854
rect 59546 -3462 59782 -3226
rect 59866 -3462 60102 -3226
rect 59546 -3782 59782 -3546
rect 59866 -3782 60102 -3546
rect 63266 28658 63502 28894
rect 63586 28658 63822 28894
rect 63266 28338 63502 28574
rect 63586 28338 63822 28574
rect 63266 -5382 63502 -5146
rect 63586 -5382 63822 -5146
rect 63266 -5702 63502 -5466
rect 63586 -5702 63822 -5466
rect 66986 32378 67222 32614
rect 67306 32378 67542 32614
rect 66986 32058 67222 32294
rect 67306 32058 67542 32294
rect 48986 -6342 49222 -6106
rect 49306 -6342 49542 -6106
rect 48986 -6662 49222 -6426
rect 49306 -6662 49542 -6426
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 42938 77782 43174
rect 77866 42938 78102 43174
rect 77546 42618 77782 42854
rect 77866 42618 78102 42854
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -2502 77782 -2266
rect 77866 -2502 78102 -2266
rect 77546 -2822 77782 -2586
rect 77866 -2822 78102 -2586
rect 81266 46658 81502 46894
rect 81586 46658 81822 46894
rect 81266 46338 81502 46574
rect 81586 46338 81822 46574
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -4422 81502 -4186
rect 81586 -4422 81822 -4186
rect 81266 -4742 81502 -4506
rect 81586 -4742 81822 -4506
rect 84986 50378 85222 50614
rect 85306 50378 85542 50614
rect 84986 50058 85222 50294
rect 85306 50058 85542 50294
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 66986 -7302 67222 -7066
rect 67306 -7302 67542 -7066
rect 66986 -7622 67222 -7386
rect 67306 -7622 67542 -7386
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -1542 92062 -1306
rect 92146 -1542 92382 -1306
rect 91826 -1862 92062 -1626
rect 92146 -1862 92382 -1626
rect 95546 24938 95782 25174
rect 95866 24938 96102 25174
rect 95546 24618 95782 24854
rect 95866 24618 96102 24854
rect 95546 -3462 95782 -3226
rect 95866 -3462 96102 -3226
rect 95546 -3782 95782 -3546
rect 95866 -3782 96102 -3546
rect 99266 28658 99502 28894
rect 99586 28658 99822 28894
rect 99266 28338 99502 28574
rect 99586 28338 99822 28574
rect 99266 -5382 99502 -5146
rect 99586 -5382 99822 -5146
rect 99266 -5702 99502 -5466
rect 99586 -5702 99822 -5466
rect 102986 32378 103222 32614
rect 103306 32378 103542 32614
rect 102986 32058 103222 32294
rect 103306 32058 103542 32294
rect 84986 -6342 85222 -6106
rect 85306 -6342 85542 -6106
rect 84986 -6662 85222 -6426
rect 85306 -6662 85542 -6426
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 42938 113782 43174
rect 113866 42938 114102 43174
rect 113546 42618 113782 42854
rect 113866 42618 114102 42854
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -2502 113782 -2266
rect 113866 -2502 114102 -2266
rect 113546 -2822 113782 -2586
rect 113866 -2822 114102 -2586
rect 117266 46658 117502 46894
rect 117586 46658 117822 46894
rect 117266 46338 117502 46574
rect 117586 46338 117822 46574
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -4422 117502 -4186
rect 117586 -4422 117822 -4186
rect 117266 -4742 117502 -4506
rect 117586 -4742 117822 -4506
rect 120986 50378 121222 50614
rect 121306 50378 121542 50614
rect 120986 50058 121222 50294
rect 121306 50058 121542 50294
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 102986 -7302 103222 -7066
rect 103306 -7302 103542 -7066
rect 102986 -7622 103222 -7386
rect 103306 -7622 103542 -7386
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -1542 128062 -1306
rect 128146 -1542 128382 -1306
rect 127826 -1862 128062 -1626
rect 128146 -1862 128382 -1626
rect 131546 24938 131782 25174
rect 131866 24938 132102 25174
rect 131546 24618 131782 24854
rect 131866 24618 132102 24854
rect 131546 -3462 131782 -3226
rect 131866 -3462 132102 -3226
rect 131546 -3782 131782 -3546
rect 131866 -3782 132102 -3546
rect 135266 28658 135502 28894
rect 135586 28658 135822 28894
rect 135266 28338 135502 28574
rect 135586 28338 135822 28574
rect 135266 -5382 135502 -5146
rect 135586 -5382 135822 -5146
rect 135266 -5702 135502 -5466
rect 135586 -5702 135822 -5466
rect 138986 32378 139222 32614
rect 139306 32378 139542 32614
rect 138986 32058 139222 32294
rect 139306 32058 139542 32294
rect 120986 -6342 121222 -6106
rect 121306 -6342 121542 -6106
rect 120986 -6662 121222 -6426
rect 121306 -6662 121542 -6426
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 42938 149782 43174
rect 149866 42938 150102 43174
rect 149546 42618 149782 42854
rect 149866 42618 150102 42854
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -2502 149782 -2266
rect 149866 -2502 150102 -2266
rect 149546 -2822 149782 -2586
rect 149866 -2822 150102 -2586
rect 153266 46658 153502 46894
rect 153586 46658 153822 46894
rect 153266 46338 153502 46574
rect 153586 46338 153822 46574
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -4422 153502 -4186
rect 153586 -4422 153822 -4186
rect 153266 -4742 153502 -4506
rect 153586 -4742 153822 -4506
rect 156986 50378 157222 50614
rect 157306 50378 157542 50614
rect 156986 50058 157222 50294
rect 157306 50058 157542 50294
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 138986 -7302 139222 -7066
rect 139306 -7302 139542 -7066
rect 138986 -7622 139222 -7386
rect 139306 -7622 139542 -7386
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -1542 164062 -1306
rect 164146 -1542 164382 -1306
rect 163826 -1862 164062 -1626
rect 164146 -1862 164382 -1626
rect 167546 24938 167782 25174
rect 167866 24938 168102 25174
rect 167546 24618 167782 24854
rect 167866 24618 168102 24854
rect 167546 -3462 167782 -3226
rect 167866 -3462 168102 -3226
rect 167546 -3782 167782 -3546
rect 167866 -3782 168102 -3546
rect 171266 28658 171502 28894
rect 171586 28658 171822 28894
rect 171266 28338 171502 28574
rect 171586 28338 171822 28574
rect 171266 -5382 171502 -5146
rect 171586 -5382 171822 -5146
rect 171266 -5702 171502 -5466
rect 171586 -5702 171822 -5466
rect 174986 32378 175222 32614
rect 175306 32378 175542 32614
rect 174986 32058 175222 32294
rect 175306 32058 175542 32294
rect 156986 -6342 157222 -6106
rect 157306 -6342 157542 -6106
rect 156986 -6662 157222 -6426
rect 157306 -6662 157542 -6426
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 42938 185782 43174
rect 185866 42938 186102 43174
rect 185546 42618 185782 42854
rect 185866 42618 186102 42854
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -2502 185782 -2266
rect 185866 -2502 186102 -2266
rect 185546 -2822 185782 -2586
rect 185866 -2822 186102 -2586
rect 189266 46658 189502 46894
rect 189586 46658 189822 46894
rect 189266 46338 189502 46574
rect 189586 46338 189822 46574
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -4422 189502 -4186
rect 189586 -4422 189822 -4186
rect 189266 -4742 189502 -4506
rect 189586 -4742 189822 -4506
rect 192986 50378 193222 50614
rect 193306 50378 193542 50614
rect 192986 50058 193222 50294
rect 193306 50058 193542 50294
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 174986 -7302 175222 -7066
rect 175306 -7302 175542 -7066
rect 174986 -7622 175222 -7386
rect 175306 -7622 175542 -7386
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -1542 200062 -1306
rect 200146 -1542 200382 -1306
rect 199826 -1862 200062 -1626
rect 200146 -1862 200382 -1626
rect 203546 24938 203782 25174
rect 203866 24938 204102 25174
rect 203546 24618 203782 24854
rect 203866 24618 204102 24854
rect 203546 -3462 203782 -3226
rect 203866 -3462 204102 -3226
rect 203546 -3782 203782 -3546
rect 203866 -3782 204102 -3546
rect 207266 28658 207502 28894
rect 207586 28658 207822 28894
rect 207266 28338 207502 28574
rect 207586 28338 207822 28574
rect 207266 -5382 207502 -5146
rect 207586 -5382 207822 -5146
rect 207266 -5702 207502 -5466
rect 207586 -5702 207822 -5466
rect 210986 32378 211222 32614
rect 211306 32378 211542 32614
rect 210986 32058 211222 32294
rect 211306 32058 211542 32294
rect 192986 -6342 193222 -6106
rect 193306 -6342 193542 -6106
rect 192986 -6662 193222 -6426
rect 193306 -6662 193542 -6426
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 42938 221782 43174
rect 221866 42938 222102 43174
rect 221546 42618 221782 42854
rect 221866 42618 222102 42854
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -2502 221782 -2266
rect 221866 -2502 222102 -2266
rect 221546 -2822 221782 -2586
rect 221866 -2822 222102 -2586
rect 228986 374378 229222 374614
rect 229306 374378 229542 374614
rect 228986 374058 229222 374294
rect 229306 374058 229542 374294
rect 228986 338378 229222 338614
rect 229306 338378 229542 338614
rect 228986 338058 229222 338294
rect 229306 338058 229542 338294
rect 228986 302378 229222 302614
rect 229306 302378 229542 302614
rect 228986 302058 229222 302294
rect 229306 302058 229542 302294
rect 228986 266378 229222 266614
rect 229306 266378 229542 266614
rect 228986 266058 229222 266294
rect 229306 266058 229542 266294
rect 228986 230378 229222 230614
rect 229306 230378 229542 230614
rect 228986 230058 229222 230294
rect 229306 230058 229542 230294
rect 228986 194378 229222 194614
rect 229306 194378 229542 194614
rect 228986 194058 229222 194294
rect 229306 194058 229542 194294
rect 228986 158378 229222 158614
rect 229306 158378 229542 158614
rect 228986 158058 229222 158294
rect 229306 158058 229542 158294
rect 228986 122378 229222 122614
rect 229306 122378 229542 122614
rect 228986 122058 229222 122294
rect 229306 122058 229542 122294
rect 228986 86378 229222 86614
rect 229306 86378 229542 86614
rect 228986 86058 229222 86294
rect 229306 86058 229542 86294
rect 225266 46658 225502 46894
rect 225586 46658 225822 46894
rect 225266 46338 225502 46574
rect 225586 46338 225822 46574
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -4422 225502 -4186
rect 225586 -4422 225822 -4186
rect 225266 -4742 225502 -4506
rect 225586 -4742 225822 -4506
rect 228986 50378 229222 50614
rect 229306 50378 229542 50614
rect 228986 50058 229222 50294
rect 229306 50058 229542 50294
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 210986 -7302 211222 -7066
rect 211306 -7302 211542 -7066
rect 210986 -7622 211222 -7386
rect 211306 -7622 211542 -7386
rect 235826 381218 236062 381454
rect 236146 381218 236382 381454
rect 235826 380898 236062 381134
rect 236146 380898 236382 381134
rect 235826 345218 236062 345454
rect 236146 345218 236382 345454
rect 235826 344898 236062 345134
rect 236146 344898 236382 345134
rect 235826 309218 236062 309454
rect 236146 309218 236382 309454
rect 235826 308898 236062 309134
rect 236146 308898 236382 309134
rect 235826 273218 236062 273454
rect 236146 273218 236382 273454
rect 235826 272898 236062 273134
rect 236146 272898 236382 273134
rect 235826 237218 236062 237454
rect 236146 237218 236382 237454
rect 235826 236898 236062 237134
rect 236146 236898 236382 237134
rect 235826 201218 236062 201454
rect 236146 201218 236382 201454
rect 235826 200898 236062 201134
rect 236146 200898 236382 201134
rect 235826 165218 236062 165454
rect 236146 165218 236382 165454
rect 235826 164898 236062 165134
rect 236146 164898 236382 165134
rect 235826 129218 236062 129454
rect 236146 129218 236382 129454
rect 235826 128898 236062 129134
rect 236146 128898 236382 129134
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -1542 236062 -1306
rect 236146 -1542 236382 -1306
rect 235826 -1862 236062 -1626
rect 236146 -1862 236382 -1626
rect 239546 384938 239782 385174
rect 239866 384938 240102 385174
rect 239546 384618 239782 384854
rect 239866 384618 240102 384854
rect 239546 348938 239782 349174
rect 239866 348938 240102 349174
rect 239546 348618 239782 348854
rect 239866 348618 240102 348854
rect 239546 312938 239782 313174
rect 239866 312938 240102 313174
rect 239546 312618 239782 312854
rect 239866 312618 240102 312854
rect 239546 276938 239782 277174
rect 239866 276938 240102 277174
rect 239546 276618 239782 276854
rect 239866 276618 240102 276854
rect 239546 240938 239782 241174
rect 239866 240938 240102 241174
rect 239546 240618 239782 240854
rect 239866 240618 240102 240854
rect 239546 204938 239782 205174
rect 239866 204938 240102 205174
rect 239546 204618 239782 204854
rect 239866 204618 240102 204854
rect 239546 168938 239782 169174
rect 239866 168938 240102 169174
rect 239546 168618 239782 168854
rect 239866 168618 240102 168854
rect 239546 132938 239782 133174
rect 239866 132938 240102 133174
rect 239546 132618 239782 132854
rect 239866 132618 240102 132854
rect 239546 96938 239782 97174
rect 239866 96938 240102 97174
rect 239546 96618 239782 96854
rect 239866 96618 240102 96854
rect 239546 60938 239782 61174
rect 239866 60938 240102 61174
rect 239546 60618 239782 60854
rect 239866 60618 240102 60854
rect 239546 24938 239782 25174
rect 239866 24938 240102 25174
rect 239546 24618 239782 24854
rect 239866 24618 240102 24854
rect 239546 -3462 239782 -3226
rect 239866 -3462 240102 -3226
rect 239546 -3782 239782 -3546
rect 239866 -3782 240102 -3546
rect 243266 388658 243502 388894
rect 243586 388658 243822 388894
rect 243266 388338 243502 388574
rect 243586 388338 243822 388574
rect 243266 352658 243502 352894
rect 243586 352658 243822 352894
rect 243266 352338 243502 352574
rect 243586 352338 243822 352574
rect 243266 316658 243502 316894
rect 243586 316658 243822 316894
rect 243266 316338 243502 316574
rect 243586 316338 243822 316574
rect 243266 280658 243502 280894
rect 243586 280658 243822 280894
rect 243266 280338 243502 280574
rect 243586 280338 243822 280574
rect 243266 244658 243502 244894
rect 243586 244658 243822 244894
rect 243266 244338 243502 244574
rect 243586 244338 243822 244574
rect 243266 208658 243502 208894
rect 243586 208658 243822 208894
rect 243266 208338 243502 208574
rect 243586 208338 243822 208574
rect 243266 172658 243502 172894
rect 243586 172658 243822 172894
rect 243266 172338 243502 172574
rect 243586 172338 243822 172574
rect 243266 136658 243502 136894
rect 243586 136658 243822 136894
rect 243266 136338 243502 136574
rect 243586 136338 243822 136574
rect 243266 100658 243502 100894
rect 243586 100658 243822 100894
rect 243266 100338 243502 100574
rect 243586 100338 243822 100574
rect 243266 64658 243502 64894
rect 243586 64658 243822 64894
rect 243266 64338 243502 64574
rect 243586 64338 243822 64574
rect 243266 28658 243502 28894
rect 243586 28658 243822 28894
rect 243266 28338 243502 28574
rect 243586 28338 243822 28574
rect 243266 -5382 243502 -5146
rect 243586 -5382 243822 -5146
rect 243266 -5702 243502 -5466
rect 243586 -5702 243822 -5466
rect 246986 392378 247222 392614
rect 247306 392378 247542 392614
rect 246986 392058 247222 392294
rect 247306 392058 247542 392294
rect 246986 356378 247222 356614
rect 247306 356378 247542 356614
rect 246986 356058 247222 356294
rect 247306 356058 247542 356294
rect 246986 320378 247222 320614
rect 247306 320378 247542 320614
rect 246986 320058 247222 320294
rect 247306 320058 247542 320294
rect 246986 284378 247222 284614
rect 247306 284378 247542 284614
rect 246986 284058 247222 284294
rect 247306 284058 247542 284294
rect 246986 248378 247222 248614
rect 247306 248378 247542 248614
rect 246986 248058 247222 248294
rect 247306 248058 247542 248294
rect 246986 212378 247222 212614
rect 247306 212378 247542 212614
rect 246986 212058 247222 212294
rect 247306 212058 247542 212294
rect 246986 176378 247222 176614
rect 247306 176378 247542 176614
rect 246986 176058 247222 176294
rect 247306 176058 247542 176294
rect 246986 140378 247222 140614
rect 247306 140378 247542 140614
rect 246986 140058 247222 140294
rect 247306 140058 247542 140294
rect 246986 104378 247222 104614
rect 247306 104378 247542 104614
rect 246986 104058 247222 104294
rect 247306 104058 247542 104294
rect 246986 68378 247222 68614
rect 247306 68378 247542 68614
rect 246986 68058 247222 68294
rect 247306 68058 247542 68294
rect 246986 32378 247222 32614
rect 247306 32378 247542 32614
rect 246986 32058 247222 32294
rect 247306 32058 247542 32294
rect 228986 -6342 229222 -6106
rect 229306 -6342 229542 -6106
rect 228986 -6662 229222 -6426
rect 229306 -6662 229542 -6426
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 253826 327218 254062 327454
rect 254146 327218 254382 327454
rect 253826 326898 254062 327134
rect 254146 326898 254382 327134
rect 253826 291218 254062 291454
rect 254146 291218 254382 291454
rect 253826 290898 254062 291134
rect 254146 290898 254382 291134
rect 253826 255218 254062 255454
rect 254146 255218 254382 255454
rect 253826 254898 254062 255134
rect 254146 254898 254382 255134
rect 253826 219218 254062 219454
rect 254146 219218 254382 219454
rect 253826 218898 254062 219134
rect 254146 218898 254382 219134
rect 253826 183218 254062 183454
rect 254146 183218 254382 183454
rect 253826 182898 254062 183134
rect 254146 182898 254382 183134
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 366938 257782 367174
rect 257866 366938 258102 367174
rect 257546 366618 257782 366854
rect 257866 366618 258102 366854
rect 257546 330938 257782 331174
rect 257866 330938 258102 331174
rect 257546 330618 257782 330854
rect 257866 330618 258102 330854
rect 257546 294938 257782 295174
rect 257866 294938 258102 295174
rect 257546 294618 257782 294854
rect 257866 294618 258102 294854
rect 257546 258938 257782 259174
rect 257866 258938 258102 259174
rect 257546 258618 257782 258854
rect 257866 258618 258102 258854
rect 257546 222938 257782 223174
rect 257866 222938 258102 223174
rect 257546 222618 257782 222854
rect 257866 222618 258102 222854
rect 257546 186938 257782 187174
rect 257866 186938 258102 187174
rect 257546 186618 257782 186854
rect 257866 186618 258102 186854
rect 257546 150938 257782 151174
rect 257866 150938 258102 151174
rect 257546 150618 257782 150854
rect 257866 150618 258102 150854
rect 257546 114938 257782 115174
rect 257866 114938 258102 115174
rect 257546 114618 257782 114854
rect 257866 114618 258102 114854
rect 257546 78938 257782 79174
rect 257866 78938 258102 79174
rect 257546 78618 257782 78854
rect 257866 78618 258102 78854
rect 257546 42938 257782 43174
rect 257866 42938 258102 43174
rect 257546 42618 257782 42854
rect 257866 42618 258102 42854
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -2502 257782 -2266
rect 257866 -2502 258102 -2266
rect 257546 -2822 257782 -2586
rect 257866 -2822 258102 -2586
rect 261266 370658 261502 370894
rect 261586 370658 261822 370894
rect 261266 370338 261502 370574
rect 261586 370338 261822 370574
rect 261266 334658 261502 334894
rect 261586 334658 261822 334894
rect 261266 334338 261502 334574
rect 261586 334338 261822 334574
rect 261266 298658 261502 298894
rect 261586 298658 261822 298894
rect 261266 298338 261502 298574
rect 261586 298338 261822 298574
rect 261266 262658 261502 262894
rect 261586 262658 261822 262894
rect 261266 262338 261502 262574
rect 261586 262338 261822 262574
rect 261266 226658 261502 226894
rect 261586 226658 261822 226894
rect 261266 226338 261502 226574
rect 261586 226338 261822 226574
rect 261266 190658 261502 190894
rect 261586 190658 261822 190894
rect 261266 190338 261502 190574
rect 261586 190338 261822 190574
rect 261266 154658 261502 154894
rect 261586 154658 261822 154894
rect 261266 154338 261502 154574
rect 261586 154338 261822 154574
rect 261266 118658 261502 118894
rect 261586 118658 261822 118894
rect 261266 118338 261502 118574
rect 261586 118338 261822 118574
rect 261266 82658 261502 82894
rect 261586 82658 261822 82894
rect 261266 82338 261502 82574
rect 261586 82338 261822 82574
rect 261266 46658 261502 46894
rect 261586 46658 261822 46894
rect 261266 46338 261502 46574
rect 261586 46338 261822 46574
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -4422 261502 -4186
rect 261586 -4422 261822 -4186
rect 261266 -4742 261502 -4506
rect 261586 -4742 261822 -4506
rect 264986 374378 265222 374614
rect 265306 374378 265542 374614
rect 264986 374058 265222 374294
rect 265306 374058 265542 374294
rect 264986 338378 265222 338614
rect 265306 338378 265542 338614
rect 264986 338058 265222 338294
rect 265306 338058 265542 338294
rect 264986 302378 265222 302614
rect 265306 302378 265542 302614
rect 264986 302058 265222 302294
rect 265306 302058 265542 302294
rect 264986 266378 265222 266614
rect 265306 266378 265542 266614
rect 264986 266058 265222 266294
rect 265306 266058 265542 266294
rect 264986 230378 265222 230614
rect 265306 230378 265542 230614
rect 264986 230058 265222 230294
rect 265306 230058 265542 230294
rect 264986 194378 265222 194614
rect 265306 194378 265542 194614
rect 264986 194058 265222 194294
rect 265306 194058 265542 194294
rect 264986 158378 265222 158614
rect 265306 158378 265542 158614
rect 264986 158058 265222 158294
rect 265306 158058 265542 158294
rect 264986 122378 265222 122614
rect 265306 122378 265542 122614
rect 264986 122058 265222 122294
rect 265306 122058 265542 122294
rect 264986 86378 265222 86614
rect 265306 86378 265542 86614
rect 264986 86058 265222 86294
rect 265306 86058 265542 86294
rect 264986 50378 265222 50614
rect 265306 50378 265542 50614
rect 264986 50058 265222 50294
rect 265306 50058 265542 50294
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 246986 -7302 247222 -7066
rect 247306 -7302 247542 -7066
rect 246986 -7622 247222 -7386
rect 247306 -7622 247542 -7386
rect 271826 381218 272062 381454
rect 272146 381218 272382 381454
rect 271826 380898 272062 381134
rect 272146 380898 272382 381134
rect 271826 345218 272062 345454
rect 272146 345218 272382 345454
rect 271826 344898 272062 345134
rect 272146 344898 272382 345134
rect 271826 309218 272062 309454
rect 272146 309218 272382 309454
rect 271826 308898 272062 309134
rect 272146 308898 272382 309134
rect 271826 273218 272062 273454
rect 272146 273218 272382 273454
rect 271826 272898 272062 273134
rect 272146 272898 272382 273134
rect 271826 237218 272062 237454
rect 272146 237218 272382 237454
rect 271826 236898 272062 237134
rect 272146 236898 272382 237134
rect 271826 201218 272062 201454
rect 272146 201218 272382 201454
rect 271826 200898 272062 201134
rect 272146 200898 272382 201134
rect 271826 165218 272062 165454
rect 272146 165218 272382 165454
rect 271826 164898 272062 165134
rect 272146 164898 272382 165134
rect 271826 129218 272062 129454
rect 272146 129218 272382 129454
rect 271826 128898 272062 129134
rect 272146 128898 272382 129134
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -1542 272062 -1306
rect 272146 -1542 272382 -1306
rect 271826 -1862 272062 -1626
rect 272146 -1862 272382 -1626
rect 275546 384938 275782 385174
rect 275866 384938 276102 385174
rect 275546 384618 275782 384854
rect 275866 384618 276102 384854
rect 275546 348938 275782 349174
rect 275866 348938 276102 349174
rect 275546 348618 275782 348854
rect 275866 348618 276102 348854
rect 275546 312938 275782 313174
rect 275866 312938 276102 313174
rect 275546 312618 275782 312854
rect 275866 312618 276102 312854
rect 275546 276938 275782 277174
rect 275866 276938 276102 277174
rect 275546 276618 275782 276854
rect 275866 276618 276102 276854
rect 275546 240938 275782 241174
rect 275866 240938 276102 241174
rect 275546 240618 275782 240854
rect 275866 240618 276102 240854
rect 275546 204938 275782 205174
rect 275866 204938 276102 205174
rect 275546 204618 275782 204854
rect 275866 204618 276102 204854
rect 275546 168938 275782 169174
rect 275866 168938 276102 169174
rect 275546 168618 275782 168854
rect 275866 168618 276102 168854
rect 275546 132938 275782 133174
rect 275866 132938 276102 133174
rect 275546 132618 275782 132854
rect 275866 132618 276102 132854
rect 275546 96938 275782 97174
rect 275866 96938 276102 97174
rect 275546 96618 275782 96854
rect 275866 96618 276102 96854
rect 275546 60938 275782 61174
rect 275866 60938 276102 61174
rect 275546 60618 275782 60854
rect 275866 60618 276102 60854
rect 275546 24938 275782 25174
rect 275866 24938 276102 25174
rect 275546 24618 275782 24854
rect 275866 24618 276102 24854
rect 275546 -3462 275782 -3226
rect 275866 -3462 276102 -3226
rect 275546 -3782 275782 -3546
rect 275866 -3782 276102 -3546
rect 279266 388658 279502 388894
rect 279586 388658 279822 388894
rect 279266 388338 279502 388574
rect 279586 388338 279822 388574
rect 279266 352658 279502 352894
rect 279586 352658 279822 352894
rect 279266 352338 279502 352574
rect 279586 352338 279822 352574
rect 279266 316658 279502 316894
rect 279586 316658 279822 316894
rect 279266 316338 279502 316574
rect 279586 316338 279822 316574
rect 279266 280658 279502 280894
rect 279586 280658 279822 280894
rect 279266 280338 279502 280574
rect 279586 280338 279822 280574
rect 279266 244658 279502 244894
rect 279586 244658 279822 244894
rect 279266 244338 279502 244574
rect 279586 244338 279822 244574
rect 279266 208658 279502 208894
rect 279586 208658 279822 208894
rect 279266 208338 279502 208574
rect 279586 208338 279822 208574
rect 279266 172658 279502 172894
rect 279586 172658 279822 172894
rect 279266 172338 279502 172574
rect 279586 172338 279822 172574
rect 279266 136658 279502 136894
rect 279586 136658 279822 136894
rect 279266 136338 279502 136574
rect 279586 136338 279822 136574
rect 279266 100658 279502 100894
rect 279586 100658 279822 100894
rect 279266 100338 279502 100574
rect 279586 100338 279822 100574
rect 279266 64658 279502 64894
rect 279586 64658 279822 64894
rect 279266 64338 279502 64574
rect 279586 64338 279822 64574
rect 279266 28658 279502 28894
rect 279586 28658 279822 28894
rect 279266 28338 279502 28574
rect 279586 28338 279822 28574
rect 279266 -5382 279502 -5146
rect 279586 -5382 279822 -5146
rect 279266 -5702 279502 -5466
rect 279586 -5702 279822 -5466
rect 282986 392378 283222 392614
rect 283306 392378 283542 392614
rect 282986 392058 283222 392294
rect 283306 392058 283542 392294
rect 282986 356378 283222 356614
rect 283306 356378 283542 356614
rect 282986 356058 283222 356294
rect 283306 356058 283542 356294
rect 282986 320378 283222 320614
rect 283306 320378 283542 320614
rect 282986 320058 283222 320294
rect 283306 320058 283542 320294
rect 282986 284378 283222 284614
rect 283306 284378 283542 284614
rect 282986 284058 283222 284294
rect 283306 284058 283542 284294
rect 282986 248378 283222 248614
rect 283306 248378 283542 248614
rect 282986 248058 283222 248294
rect 283306 248058 283542 248294
rect 282986 212378 283222 212614
rect 283306 212378 283542 212614
rect 282986 212058 283222 212294
rect 283306 212058 283542 212294
rect 282986 176378 283222 176614
rect 283306 176378 283542 176614
rect 282986 176058 283222 176294
rect 283306 176058 283542 176294
rect 282986 140378 283222 140614
rect 283306 140378 283542 140614
rect 282986 140058 283222 140294
rect 283306 140058 283542 140294
rect 282986 104378 283222 104614
rect 283306 104378 283542 104614
rect 282986 104058 283222 104294
rect 283306 104058 283542 104294
rect 282986 68378 283222 68614
rect 283306 68378 283542 68614
rect 282986 68058 283222 68294
rect 283306 68058 283542 68294
rect 282986 32378 283222 32614
rect 283306 32378 283542 32614
rect 282986 32058 283222 32294
rect 283306 32058 283542 32294
rect 264986 -6342 265222 -6106
rect 265306 -6342 265542 -6106
rect 264986 -6662 265222 -6426
rect 265306 -6662 265542 -6426
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 289826 327218 290062 327454
rect 290146 327218 290382 327454
rect 289826 326898 290062 327134
rect 290146 326898 290382 327134
rect 289826 291218 290062 291454
rect 290146 291218 290382 291454
rect 289826 290898 290062 291134
rect 290146 290898 290382 291134
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 289826 219218 290062 219454
rect 290146 219218 290382 219454
rect 289826 218898 290062 219134
rect 290146 218898 290382 219134
rect 289826 183218 290062 183454
rect 290146 183218 290382 183454
rect 289826 182898 290062 183134
rect 290146 182898 290382 183134
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 366938 293782 367174
rect 293866 366938 294102 367174
rect 293546 366618 293782 366854
rect 293866 366618 294102 366854
rect 293546 330938 293782 331174
rect 293866 330938 294102 331174
rect 293546 330618 293782 330854
rect 293866 330618 294102 330854
rect 293546 294938 293782 295174
rect 293866 294938 294102 295174
rect 293546 294618 293782 294854
rect 293866 294618 294102 294854
rect 293546 258938 293782 259174
rect 293866 258938 294102 259174
rect 293546 258618 293782 258854
rect 293866 258618 294102 258854
rect 293546 222938 293782 223174
rect 293866 222938 294102 223174
rect 293546 222618 293782 222854
rect 293866 222618 294102 222854
rect 293546 186938 293782 187174
rect 293866 186938 294102 187174
rect 293546 186618 293782 186854
rect 293866 186618 294102 186854
rect 293546 150938 293782 151174
rect 293866 150938 294102 151174
rect 293546 150618 293782 150854
rect 293866 150618 294102 150854
rect 293546 114938 293782 115174
rect 293866 114938 294102 115174
rect 293546 114618 293782 114854
rect 293866 114618 294102 114854
rect 293546 78938 293782 79174
rect 293866 78938 294102 79174
rect 293546 78618 293782 78854
rect 293866 78618 294102 78854
rect 293546 42938 293782 43174
rect 293866 42938 294102 43174
rect 293546 42618 293782 42854
rect 293866 42618 294102 42854
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -2502 293782 -2266
rect 293866 -2502 294102 -2266
rect 293546 -2822 293782 -2586
rect 293866 -2822 294102 -2586
rect 297266 370658 297502 370894
rect 297586 370658 297822 370894
rect 297266 370338 297502 370574
rect 297586 370338 297822 370574
rect 297266 334658 297502 334894
rect 297586 334658 297822 334894
rect 297266 334338 297502 334574
rect 297586 334338 297822 334574
rect 297266 298658 297502 298894
rect 297586 298658 297822 298894
rect 297266 298338 297502 298574
rect 297586 298338 297822 298574
rect 297266 262658 297502 262894
rect 297586 262658 297822 262894
rect 297266 262338 297502 262574
rect 297586 262338 297822 262574
rect 297266 226658 297502 226894
rect 297586 226658 297822 226894
rect 297266 226338 297502 226574
rect 297586 226338 297822 226574
rect 297266 190658 297502 190894
rect 297586 190658 297822 190894
rect 297266 190338 297502 190574
rect 297586 190338 297822 190574
rect 297266 154658 297502 154894
rect 297586 154658 297822 154894
rect 297266 154338 297502 154574
rect 297586 154338 297822 154574
rect 297266 118658 297502 118894
rect 297586 118658 297822 118894
rect 297266 118338 297502 118574
rect 297586 118338 297822 118574
rect 297266 82658 297502 82894
rect 297586 82658 297822 82894
rect 297266 82338 297502 82574
rect 297586 82338 297822 82574
rect 297266 46658 297502 46894
rect 297586 46658 297822 46894
rect 297266 46338 297502 46574
rect 297586 46338 297822 46574
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -4422 297502 -4186
rect 297586 -4422 297822 -4186
rect 297266 -4742 297502 -4506
rect 297586 -4742 297822 -4506
rect 300986 374378 301222 374614
rect 301306 374378 301542 374614
rect 300986 374058 301222 374294
rect 301306 374058 301542 374294
rect 300986 338378 301222 338614
rect 301306 338378 301542 338614
rect 300986 338058 301222 338294
rect 301306 338058 301542 338294
rect 300986 302378 301222 302614
rect 301306 302378 301542 302614
rect 300986 302058 301222 302294
rect 301306 302058 301542 302294
rect 300986 266378 301222 266614
rect 301306 266378 301542 266614
rect 300986 266058 301222 266294
rect 301306 266058 301542 266294
rect 300986 230378 301222 230614
rect 301306 230378 301542 230614
rect 300986 230058 301222 230294
rect 301306 230058 301542 230294
rect 300986 194378 301222 194614
rect 301306 194378 301542 194614
rect 300986 194058 301222 194294
rect 301306 194058 301542 194294
rect 300986 158378 301222 158614
rect 301306 158378 301542 158614
rect 300986 158058 301222 158294
rect 301306 158058 301542 158294
rect 300986 122378 301222 122614
rect 301306 122378 301542 122614
rect 300986 122058 301222 122294
rect 301306 122058 301542 122294
rect 300986 86378 301222 86614
rect 301306 86378 301542 86614
rect 300986 86058 301222 86294
rect 301306 86058 301542 86294
rect 300986 50378 301222 50614
rect 301306 50378 301542 50614
rect 300986 50058 301222 50294
rect 301306 50058 301542 50294
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 282986 -7302 283222 -7066
rect 283306 -7302 283542 -7066
rect 282986 -7622 283222 -7386
rect 283306 -7622 283542 -7386
rect 307826 381218 308062 381454
rect 308146 381218 308382 381454
rect 307826 380898 308062 381134
rect 308146 380898 308382 381134
rect 307826 345218 308062 345454
rect 308146 345218 308382 345454
rect 307826 344898 308062 345134
rect 308146 344898 308382 345134
rect 307826 309218 308062 309454
rect 308146 309218 308382 309454
rect 307826 308898 308062 309134
rect 308146 308898 308382 309134
rect 307826 273218 308062 273454
rect 308146 273218 308382 273454
rect 307826 272898 308062 273134
rect 308146 272898 308382 273134
rect 307826 237218 308062 237454
rect 308146 237218 308382 237454
rect 307826 236898 308062 237134
rect 308146 236898 308382 237134
rect 307826 201218 308062 201454
rect 308146 201218 308382 201454
rect 307826 200898 308062 201134
rect 308146 200898 308382 201134
rect 307826 165218 308062 165454
rect 308146 165218 308382 165454
rect 307826 164898 308062 165134
rect 308146 164898 308382 165134
rect 307826 129218 308062 129454
rect 308146 129218 308382 129454
rect 307826 128898 308062 129134
rect 308146 128898 308382 129134
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -1542 308062 -1306
rect 308146 -1542 308382 -1306
rect 307826 -1862 308062 -1626
rect 308146 -1862 308382 -1626
rect 311546 384938 311782 385174
rect 311866 384938 312102 385174
rect 311546 384618 311782 384854
rect 311866 384618 312102 384854
rect 311546 348938 311782 349174
rect 311866 348938 312102 349174
rect 311546 348618 311782 348854
rect 311866 348618 312102 348854
rect 311546 312938 311782 313174
rect 311866 312938 312102 313174
rect 311546 312618 311782 312854
rect 311866 312618 312102 312854
rect 311546 276938 311782 277174
rect 311866 276938 312102 277174
rect 311546 276618 311782 276854
rect 311866 276618 312102 276854
rect 311546 240938 311782 241174
rect 311866 240938 312102 241174
rect 311546 240618 311782 240854
rect 311866 240618 312102 240854
rect 311546 204938 311782 205174
rect 311866 204938 312102 205174
rect 311546 204618 311782 204854
rect 311866 204618 312102 204854
rect 311546 168938 311782 169174
rect 311866 168938 312102 169174
rect 311546 168618 311782 168854
rect 311866 168618 312102 168854
rect 311546 132938 311782 133174
rect 311866 132938 312102 133174
rect 311546 132618 311782 132854
rect 311866 132618 312102 132854
rect 311546 96938 311782 97174
rect 311866 96938 312102 97174
rect 311546 96618 311782 96854
rect 311866 96618 312102 96854
rect 311546 60938 311782 61174
rect 311866 60938 312102 61174
rect 311546 60618 311782 60854
rect 311866 60618 312102 60854
rect 311546 24938 311782 25174
rect 311866 24938 312102 25174
rect 311546 24618 311782 24854
rect 311866 24618 312102 24854
rect 311546 -3462 311782 -3226
rect 311866 -3462 312102 -3226
rect 311546 -3782 311782 -3546
rect 311866 -3782 312102 -3546
rect 315266 388658 315502 388894
rect 315586 388658 315822 388894
rect 315266 388338 315502 388574
rect 315586 388338 315822 388574
rect 315266 352658 315502 352894
rect 315586 352658 315822 352894
rect 315266 352338 315502 352574
rect 315586 352338 315822 352574
rect 315266 316658 315502 316894
rect 315586 316658 315822 316894
rect 315266 316338 315502 316574
rect 315586 316338 315822 316574
rect 315266 280658 315502 280894
rect 315586 280658 315822 280894
rect 315266 280338 315502 280574
rect 315586 280338 315822 280574
rect 315266 244658 315502 244894
rect 315586 244658 315822 244894
rect 315266 244338 315502 244574
rect 315586 244338 315822 244574
rect 315266 208658 315502 208894
rect 315586 208658 315822 208894
rect 315266 208338 315502 208574
rect 315586 208338 315822 208574
rect 315266 172658 315502 172894
rect 315586 172658 315822 172894
rect 315266 172338 315502 172574
rect 315586 172338 315822 172574
rect 315266 136658 315502 136894
rect 315586 136658 315822 136894
rect 315266 136338 315502 136574
rect 315586 136338 315822 136574
rect 315266 100658 315502 100894
rect 315586 100658 315822 100894
rect 315266 100338 315502 100574
rect 315586 100338 315822 100574
rect 315266 64658 315502 64894
rect 315586 64658 315822 64894
rect 315266 64338 315502 64574
rect 315586 64338 315822 64574
rect 315266 28658 315502 28894
rect 315586 28658 315822 28894
rect 315266 28338 315502 28574
rect 315586 28338 315822 28574
rect 315266 -5382 315502 -5146
rect 315586 -5382 315822 -5146
rect 315266 -5702 315502 -5466
rect 315586 -5702 315822 -5466
rect 318986 392378 319222 392614
rect 319306 392378 319542 392614
rect 318986 392058 319222 392294
rect 319306 392058 319542 392294
rect 318986 356378 319222 356614
rect 319306 356378 319542 356614
rect 318986 356058 319222 356294
rect 319306 356058 319542 356294
rect 318986 320378 319222 320614
rect 319306 320378 319542 320614
rect 318986 320058 319222 320294
rect 319306 320058 319542 320294
rect 318986 284378 319222 284614
rect 319306 284378 319542 284614
rect 318986 284058 319222 284294
rect 319306 284058 319542 284294
rect 318986 248378 319222 248614
rect 319306 248378 319542 248614
rect 318986 248058 319222 248294
rect 319306 248058 319542 248294
rect 318986 212378 319222 212614
rect 319306 212378 319542 212614
rect 318986 212058 319222 212294
rect 319306 212058 319542 212294
rect 318986 176378 319222 176614
rect 319306 176378 319542 176614
rect 318986 176058 319222 176294
rect 319306 176058 319542 176294
rect 318986 140378 319222 140614
rect 319306 140378 319542 140614
rect 318986 140058 319222 140294
rect 319306 140058 319542 140294
rect 318986 104378 319222 104614
rect 319306 104378 319542 104614
rect 318986 104058 319222 104294
rect 319306 104058 319542 104294
rect 318986 68378 319222 68614
rect 319306 68378 319542 68614
rect 318986 68058 319222 68294
rect 319306 68058 319542 68294
rect 318986 32378 319222 32614
rect 319306 32378 319542 32614
rect 318986 32058 319222 32294
rect 319306 32058 319542 32294
rect 300986 -6342 301222 -6106
rect 301306 -6342 301542 -6106
rect 300986 -6662 301222 -6426
rect 301306 -6662 301542 -6426
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 325826 327218 326062 327454
rect 326146 327218 326382 327454
rect 325826 326898 326062 327134
rect 326146 326898 326382 327134
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 325826 219218 326062 219454
rect 326146 219218 326382 219454
rect 325826 218898 326062 219134
rect 326146 218898 326382 219134
rect 325826 183218 326062 183454
rect 326146 183218 326382 183454
rect 325826 182898 326062 183134
rect 326146 182898 326382 183134
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 366938 329782 367174
rect 329866 366938 330102 367174
rect 329546 366618 329782 366854
rect 329866 366618 330102 366854
rect 329546 330938 329782 331174
rect 329866 330938 330102 331174
rect 329546 330618 329782 330854
rect 329866 330618 330102 330854
rect 329546 294938 329782 295174
rect 329866 294938 330102 295174
rect 329546 294618 329782 294854
rect 329866 294618 330102 294854
rect 329546 258938 329782 259174
rect 329866 258938 330102 259174
rect 329546 258618 329782 258854
rect 329866 258618 330102 258854
rect 329546 222938 329782 223174
rect 329866 222938 330102 223174
rect 329546 222618 329782 222854
rect 329866 222618 330102 222854
rect 329546 186938 329782 187174
rect 329866 186938 330102 187174
rect 329546 186618 329782 186854
rect 329866 186618 330102 186854
rect 329546 150938 329782 151174
rect 329866 150938 330102 151174
rect 329546 150618 329782 150854
rect 329866 150618 330102 150854
rect 329546 114938 329782 115174
rect 329866 114938 330102 115174
rect 329546 114618 329782 114854
rect 329866 114618 330102 114854
rect 329546 78938 329782 79174
rect 329866 78938 330102 79174
rect 329546 78618 329782 78854
rect 329866 78618 330102 78854
rect 329546 42938 329782 43174
rect 329866 42938 330102 43174
rect 329546 42618 329782 42854
rect 329866 42618 330102 42854
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -2502 329782 -2266
rect 329866 -2502 330102 -2266
rect 329546 -2822 329782 -2586
rect 329866 -2822 330102 -2586
rect 333266 370658 333502 370894
rect 333586 370658 333822 370894
rect 333266 370338 333502 370574
rect 333586 370338 333822 370574
rect 333266 334658 333502 334894
rect 333586 334658 333822 334894
rect 333266 334338 333502 334574
rect 333586 334338 333822 334574
rect 333266 298658 333502 298894
rect 333586 298658 333822 298894
rect 333266 298338 333502 298574
rect 333586 298338 333822 298574
rect 333266 262658 333502 262894
rect 333586 262658 333822 262894
rect 333266 262338 333502 262574
rect 333586 262338 333822 262574
rect 333266 226658 333502 226894
rect 333586 226658 333822 226894
rect 333266 226338 333502 226574
rect 333586 226338 333822 226574
rect 333266 190658 333502 190894
rect 333586 190658 333822 190894
rect 333266 190338 333502 190574
rect 333586 190338 333822 190574
rect 333266 154658 333502 154894
rect 333586 154658 333822 154894
rect 333266 154338 333502 154574
rect 333586 154338 333822 154574
rect 333266 118658 333502 118894
rect 333586 118658 333822 118894
rect 333266 118338 333502 118574
rect 333586 118338 333822 118574
rect 333266 82658 333502 82894
rect 333586 82658 333822 82894
rect 333266 82338 333502 82574
rect 333586 82338 333822 82574
rect 333266 46658 333502 46894
rect 333586 46658 333822 46894
rect 333266 46338 333502 46574
rect 333586 46338 333822 46574
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -4422 333502 -4186
rect 333586 -4422 333822 -4186
rect 333266 -4742 333502 -4506
rect 333586 -4742 333822 -4506
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 336986 374378 337222 374614
rect 337306 374378 337542 374614
rect 336986 374058 337222 374294
rect 337306 374058 337542 374294
rect 336986 338378 337222 338614
rect 337306 338378 337542 338614
rect 336986 338058 337222 338294
rect 337306 338058 337542 338294
rect 336986 302378 337222 302614
rect 337306 302378 337542 302614
rect 336986 302058 337222 302294
rect 337306 302058 337542 302294
rect 336986 266378 337222 266614
rect 337306 266378 337542 266614
rect 336986 266058 337222 266294
rect 337306 266058 337542 266294
rect 336986 230378 337222 230614
rect 337306 230378 337542 230614
rect 336986 230058 337222 230294
rect 337306 230058 337542 230294
rect 336986 194378 337222 194614
rect 337306 194378 337542 194614
rect 336986 194058 337222 194294
rect 337306 194058 337542 194294
rect 336986 158378 337222 158614
rect 337306 158378 337542 158614
rect 336986 158058 337222 158294
rect 337306 158058 337542 158294
rect 336986 122378 337222 122614
rect 337306 122378 337542 122614
rect 336986 122058 337222 122294
rect 337306 122058 337542 122294
rect 336986 86378 337222 86614
rect 337306 86378 337542 86614
rect 336986 86058 337222 86294
rect 337306 86058 337542 86294
rect 336986 50378 337222 50614
rect 337306 50378 337542 50614
rect 336986 50058 337222 50294
rect 337306 50058 337542 50294
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 318986 -7302 319222 -7066
rect 319306 -7302 319542 -7066
rect 318986 -7622 319222 -7386
rect 319306 -7622 319542 -7386
rect 343826 381218 344062 381454
rect 344146 381218 344382 381454
rect 343826 380898 344062 381134
rect 344146 380898 344382 381134
rect 343826 345218 344062 345454
rect 344146 345218 344382 345454
rect 343826 344898 344062 345134
rect 344146 344898 344382 345134
rect 343826 309218 344062 309454
rect 344146 309218 344382 309454
rect 343826 308898 344062 309134
rect 344146 308898 344382 309134
rect 343826 273218 344062 273454
rect 344146 273218 344382 273454
rect 343826 272898 344062 273134
rect 344146 272898 344382 273134
rect 343826 237218 344062 237454
rect 344146 237218 344382 237454
rect 343826 236898 344062 237134
rect 344146 236898 344382 237134
rect 343826 201218 344062 201454
rect 344146 201218 344382 201454
rect 343826 200898 344062 201134
rect 344146 200898 344382 201134
rect 343826 165218 344062 165454
rect 344146 165218 344382 165454
rect 343826 164898 344062 165134
rect 344146 164898 344382 165134
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -1542 344062 -1306
rect 344146 -1542 344382 -1306
rect 343826 -1862 344062 -1626
rect 344146 -1862 344382 -1626
rect 347546 384938 347782 385174
rect 347866 384938 348102 385174
rect 347546 384618 347782 384854
rect 347866 384618 348102 384854
rect 347546 348938 347782 349174
rect 347866 348938 348102 349174
rect 347546 348618 347782 348854
rect 347866 348618 348102 348854
rect 347546 312938 347782 313174
rect 347866 312938 348102 313174
rect 347546 312618 347782 312854
rect 347866 312618 348102 312854
rect 347546 276938 347782 277174
rect 347866 276938 348102 277174
rect 347546 276618 347782 276854
rect 347866 276618 348102 276854
rect 347546 240938 347782 241174
rect 347866 240938 348102 241174
rect 347546 240618 347782 240854
rect 347866 240618 348102 240854
rect 347546 204938 347782 205174
rect 347866 204938 348102 205174
rect 347546 204618 347782 204854
rect 347866 204618 348102 204854
rect 347546 168938 347782 169174
rect 347866 168938 348102 169174
rect 347546 168618 347782 168854
rect 347866 168618 348102 168854
rect 347546 132938 347782 133174
rect 347866 132938 348102 133174
rect 347546 132618 347782 132854
rect 347866 132618 348102 132854
rect 347546 96938 347782 97174
rect 347866 96938 348102 97174
rect 347546 96618 347782 96854
rect 347866 96618 348102 96854
rect 347546 60938 347782 61174
rect 347866 60938 348102 61174
rect 347546 60618 347782 60854
rect 347866 60618 348102 60854
rect 347546 24938 347782 25174
rect 347866 24938 348102 25174
rect 347546 24618 347782 24854
rect 347866 24618 348102 24854
rect 347546 -3462 347782 -3226
rect 347866 -3462 348102 -3226
rect 347546 -3782 347782 -3546
rect 347866 -3782 348102 -3546
rect 351266 388658 351502 388894
rect 351586 388658 351822 388894
rect 351266 388338 351502 388574
rect 351586 388338 351822 388574
rect 351266 352658 351502 352894
rect 351586 352658 351822 352894
rect 351266 352338 351502 352574
rect 351586 352338 351822 352574
rect 351266 316658 351502 316894
rect 351586 316658 351822 316894
rect 351266 316338 351502 316574
rect 351586 316338 351822 316574
rect 351266 280658 351502 280894
rect 351586 280658 351822 280894
rect 351266 280338 351502 280574
rect 351586 280338 351822 280574
rect 351266 244658 351502 244894
rect 351586 244658 351822 244894
rect 351266 244338 351502 244574
rect 351586 244338 351822 244574
rect 351266 208658 351502 208894
rect 351586 208658 351822 208894
rect 351266 208338 351502 208574
rect 351586 208338 351822 208574
rect 351266 172658 351502 172894
rect 351586 172658 351822 172894
rect 351266 172338 351502 172574
rect 351586 172338 351822 172574
rect 351266 136658 351502 136894
rect 351586 136658 351822 136894
rect 351266 136338 351502 136574
rect 351586 136338 351822 136574
rect 351266 100658 351502 100894
rect 351586 100658 351822 100894
rect 351266 100338 351502 100574
rect 351586 100338 351822 100574
rect 351266 64658 351502 64894
rect 351586 64658 351822 64894
rect 351266 64338 351502 64574
rect 351586 64338 351822 64574
rect 351266 28658 351502 28894
rect 351586 28658 351822 28894
rect 351266 28338 351502 28574
rect 351586 28338 351822 28574
rect 351266 -5382 351502 -5146
rect 351586 -5382 351822 -5146
rect 351266 -5702 351502 -5466
rect 351586 -5702 351822 -5466
rect 354986 392378 355222 392614
rect 355306 392378 355542 392614
rect 354986 392058 355222 392294
rect 355306 392058 355542 392294
rect 354986 356378 355222 356614
rect 355306 356378 355542 356614
rect 354986 356058 355222 356294
rect 355306 356058 355542 356294
rect 354986 320378 355222 320614
rect 355306 320378 355542 320614
rect 354986 320058 355222 320294
rect 355306 320058 355542 320294
rect 354986 284378 355222 284614
rect 355306 284378 355542 284614
rect 354986 284058 355222 284294
rect 355306 284058 355542 284294
rect 354986 248378 355222 248614
rect 355306 248378 355542 248614
rect 354986 248058 355222 248294
rect 355306 248058 355542 248294
rect 354986 212378 355222 212614
rect 355306 212378 355542 212614
rect 354986 212058 355222 212294
rect 355306 212058 355542 212294
rect 354986 176378 355222 176614
rect 355306 176378 355542 176614
rect 354986 176058 355222 176294
rect 355306 176058 355542 176294
rect 354986 140378 355222 140614
rect 355306 140378 355542 140614
rect 354986 140058 355222 140294
rect 355306 140058 355542 140294
rect 354986 104378 355222 104614
rect 355306 104378 355542 104614
rect 354986 104058 355222 104294
rect 355306 104058 355542 104294
rect 354986 68378 355222 68614
rect 355306 68378 355542 68614
rect 354986 68058 355222 68294
rect 355306 68058 355542 68294
rect 354986 32378 355222 32614
rect 355306 32378 355542 32614
rect 354986 32058 355222 32294
rect 355306 32058 355542 32294
rect 336986 -6342 337222 -6106
rect 337306 -6342 337542 -6106
rect 336986 -6662 337222 -6426
rect 337306 -6662 337542 -6426
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 365546 618938 365782 619174
rect 365866 618938 366102 619174
rect 365546 618618 365782 618854
rect 365866 618618 366102 618854
rect 365546 582938 365782 583174
rect 365866 582938 366102 583174
rect 365546 582618 365782 582854
rect 365866 582618 366102 582854
rect 365546 546938 365782 547174
rect 365866 546938 366102 547174
rect 365546 546618 365782 546854
rect 365866 546618 366102 546854
rect 365546 510938 365782 511174
rect 365866 510938 366102 511174
rect 365546 510618 365782 510854
rect 365866 510618 366102 510854
rect 365546 474938 365782 475174
rect 365866 474938 366102 475174
rect 365546 474618 365782 474854
rect 365866 474618 366102 474854
rect 365546 438938 365782 439174
rect 365866 438938 366102 439174
rect 365546 438618 365782 438854
rect 365866 438618 366102 438854
rect 365546 402938 365782 403174
rect 365866 402938 366102 403174
rect 365546 402618 365782 402854
rect 365866 402618 366102 402854
rect 365546 366938 365782 367174
rect 365866 366938 366102 367174
rect 365546 366618 365782 366854
rect 365866 366618 366102 366854
rect 365546 330938 365782 331174
rect 365866 330938 366102 331174
rect 365546 330618 365782 330854
rect 365866 330618 366102 330854
rect 365546 294938 365782 295174
rect 365866 294938 366102 295174
rect 365546 294618 365782 294854
rect 365866 294618 366102 294854
rect 365546 258938 365782 259174
rect 365866 258938 366102 259174
rect 365546 258618 365782 258854
rect 365866 258618 366102 258854
rect 365546 222938 365782 223174
rect 365866 222938 366102 223174
rect 365546 222618 365782 222854
rect 365866 222618 366102 222854
rect 365546 186938 365782 187174
rect 365866 186938 366102 187174
rect 365546 186618 365782 186854
rect 365866 186618 366102 186854
rect 365546 150938 365782 151174
rect 365866 150938 366102 151174
rect 365546 150618 365782 150854
rect 365866 150618 366102 150854
rect 365546 114938 365782 115174
rect 365866 114938 366102 115174
rect 365546 114618 365782 114854
rect 365866 114618 366102 114854
rect 365546 78938 365782 79174
rect 365866 78938 366102 79174
rect 365546 78618 365782 78854
rect 365866 78618 366102 78854
rect 365546 42938 365782 43174
rect 365866 42938 366102 43174
rect 365546 42618 365782 42854
rect 365866 42618 366102 42854
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -2502 365782 -2266
rect 365866 -2502 366102 -2266
rect 365546 -2822 365782 -2586
rect 365866 -2822 366102 -2586
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 369266 622658 369502 622894
rect 369586 622658 369822 622894
rect 369266 622338 369502 622574
rect 369586 622338 369822 622574
rect 369266 586658 369502 586894
rect 369586 586658 369822 586894
rect 369266 586338 369502 586574
rect 369586 586338 369822 586574
rect 369266 550658 369502 550894
rect 369586 550658 369822 550894
rect 369266 550338 369502 550574
rect 369586 550338 369822 550574
rect 369266 514658 369502 514894
rect 369586 514658 369822 514894
rect 369266 514338 369502 514574
rect 369586 514338 369822 514574
rect 369266 478658 369502 478894
rect 369586 478658 369822 478894
rect 369266 478338 369502 478574
rect 369586 478338 369822 478574
rect 369266 442658 369502 442894
rect 369586 442658 369822 442894
rect 369266 442338 369502 442574
rect 369586 442338 369822 442574
rect 369266 406658 369502 406894
rect 369586 406658 369822 406894
rect 369266 406338 369502 406574
rect 369586 406338 369822 406574
rect 369266 370658 369502 370894
rect 369586 370658 369822 370894
rect 369266 370338 369502 370574
rect 369586 370338 369822 370574
rect 369266 334658 369502 334894
rect 369586 334658 369822 334894
rect 369266 334338 369502 334574
rect 369586 334338 369822 334574
rect 369266 298658 369502 298894
rect 369586 298658 369822 298894
rect 369266 298338 369502 298574
rect 369586 298338 369822 298574
rect 369266 262658 369502 262894
rect 369586 262658 369822 262894
rect 369266 262338 369502 262574
rect 369586 262338 369822 262574
rect 369266 226658 369502 226894
rect 369586 226658 369822 226894
rect 369266 226338 369502 226574
rect 369586 226338 369822 226574
rect 369266 190658 369502 190894
rect 369586 190658 369822 190894
rect 369266 190338 369502 190574
rect 369586 190338 369822 190574
rect 369266 154658 369502 154894
rect 369586 154658 369822 154894
rect 369266 154338 369502 154574
rect 369586 154338 369822 154574
rect 369266 118658 369502 118894
rect 369586 118658 369822 118894
rect 369266 118338 369502 118574
rect 369586 118338 369822 118574
rect 369266 82658 369502 82894
rect 369586 82658 369822 82894
rect 369266 82338 369502 82574
rect 369586 82338 369822 82574
rect 369266 46658 369502 46894
rect 369586 46658 369822 46894
rect 369266 46338 369502 46574
rect 369586 46338 369822 46574
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -4422 369502 -4186
rect 369586 -4422 369822 -4186
rect 369266 -4742 369502 -4506
rect 369586 -4742 369822 -4506
rect 390986 711322 391222 711558
rect 391306 711322 391542 711558
rect 390986 711002 391222 711238
rect 391306 711002 391542 711238
rect 387266 709402 387502 709638
rect 387586 709402 387822 709638
rect 387266 709082 387502 709318
rect 387586 709082 387822 709318
rect 383546 707482 383782 707718
rect 383866 707482 384102 707718
rect 383546 707162 383782 707398
rect 383866 707162 384102 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 372986 626378 373222 626614
rect 373306 626378 373542 626614
rect 372986 626058 373222 626294
rect 373306 626058 373542 626294
rect 372986 590378 373222 590614
rect 373306 590378 373542 590614
rect 372986 590058 373222 590294
rect 373306 590058 373542 590294
rect 372986 554378 373222 554614
rect 373306 554378 373542 554614
rect 372986 554058 373222 554294
rect 373306 554058 373542 554294
rect 372986 518378 373222 518614
rect 373306 518378 373542 518614
rect 372986 518058 373222 518294
rect 373306 518058 373542 518294
rect 372986 482378 373222 482614
rect 373306 482378 373542 482614
rect 372986 482058 373222 482294
rect 373306 482058 373542 482294
rect 372986 446378 373222 446614
rect 373306 446378 373542 446614
rect 372986 446058 373222 446294
rect 373306 446058 373542 446294
rect 372986 410378 373222 410614
rect 373306 410378 373542 410614
rect 372986 410058 373222 410294
rect 373306 410058 373542 410294
rect 372986 374378 373222 374614
rect 373306 374378 373542 374614
rect 372986 374058 373222 374294
rect 373306 374058 373542 374294
rect 372986 338378 373222 338614
rect 373306 338378 373542 338614
rect 372986 338058 373222 338294
rect 373306 338058 373542 338294
rect 372986 302378 373222 302614
rect 373306 302378 373542 302614
rect 372986 302058 373222 302294
rect 373306 302058 373542 302294
rect 372986 266378 373222 266614
rect 373306 266378 373542 266614
rect 372986 266058 373222 266294
rect 373306 266058 373542 266294
rect 372986 230378 373222 230614
rect 373306 230378 373542 230614
rect 372986 230058 373222 230294
rect 373306 230058 373542 230294
rect 372986 194378 373222 194614
rect 373306 194378 373542 194614
rect 372986 194058 373222 194294
rect 373306 194058 373542 194294
rect 372986 158378 373222 158614
rect 373306 158378 373542 158614
rect 372986 158058 373222 158294
rect 373306 158058 373542 158294
rect 372986 122378 373222 122614
rect 373306 122378 373542 122614
rect 372986 122058 373222 122294
rect 373306 122058 373542 122294
rect 372986 86378 373222 86614
rect 373306 86378 373542 86614
rect 372986 86058 373222 86294
rect 373306 86058 373542 86294
rect 372986 50378 373222 50614
rect 373306 50378 373542 50614
rect 372986 50058 373222 50294
rect 373306 50058 373542 50294
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 354986 -7302 355222 -7066
rect 355306 -7302 355542 -7066
rect 354986 -7622 355222 -7386
rect 355306 -7622 355542 -7386
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 379826 345218 380062 345454
rect 380146 345218 380382 345454
rect 379826 344898 380062 345134
rect 380146 344898 380382 345134
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 379826 237218 380062 237454
rect 380146 237218 380382 237454
rect 379826 236898 380062 237134
rect 380146 236898 380382 237134
rect 379826 201218 380062 201454
rect 380146 201218 380382 201454
rect 379826 200898 380062 201134
rect 380146 200898 380382 201134
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -1542 380062 -1306
rect 380146 -1542 380382 -1306
rect 379826 -1862 380062 -1626
rect 380146 -1862 380382 -1626
rect 383546 672938 383782 673174
rect 383866 672938 384102 673174
rect 383546 672618 383782 672854
rect 383866 672618 384102 672854
rect 383546 636938 383782 637174
rect 383866 636938 384102 637174
rect 383546 636618 383782 636854
rect 383866 636618 384102 636854
rect 383546 600938 383782 601174
rect 383866 600938 384102 601174
rect 383546 600618 383782 600854
rect 383866 600618 384102 600854
rect 383546 564938 383782 565174
rect 383866 564938 384102 565174
rect 383546 564618 383782 564854
rect 383866 564618 384102 564854
rect 383546 528938 383782 529174
rect 383866 528938 384102 529174
rect 383546 528618 383782 528854
rect 383866 528618 384102 528854
rect 383546 492938 383782 493174
rect 383866 492938 384102 493174
rect 383546 492618 383782 492854
rect 383866 492618 384102 492854
rect 383546 456938 383782 457174
rect 383866 456938 384102 457174
rect 383546 456618 383782 456854
rect 383866 456618 384102 456854
rect 383546 420938 383782 421174
rect 383866 420938 384102 421174
rect 383546 420618 383782 420854
rect 383866 420618 384102 420854
rect 383546 384938 383782 385174
rect 383866 384938 384102 385174
rect 383546 384618 383782 384854
rect 383866 384618 384102 384854
rect 383546 348938 383782 349174
rect 383866 348938 384102 349174
rect 383546 348618 383782 348854
rect 383866 348618 384102 348854
rect 383546 312938 383782 313174
rect 383866 312938 384102 313174
rect 383546 312618 383782 312854
rect 383866 312618 384102 312854
rect 383546 276938 383782 277174
rect 383866 276938 384102 277174
rect 383546 276618 383782 276854
rect 383866 276618 384102 276854
rect 383546 240938 383782 241174
rect 383866 240938 384102 241174
rect 383546 240618 383782 240854
rect 383866 240618 384102 240854
rect 383546 204938 383782 205174
rect 383866 204938 384102 205174
rect 383546 204618 383782 204854
rect 383866 204618 384102 204854
rect 383546 168938 383782 169174
rect 383866 168938 384102 169174
rect 383546 168618 383782 168854
rect 383866 168618 384102 168854
rect 383546 132938 383782 133174
rect 383866 132938 384102 133174
rect 383546 132618 383782 132854
rect 383866 132618 384102 132854
rect 383546 96938 383782 97174
rect 383866 96938 384102 97174
rect 383546 96618 383782 96854
rect 383866 96618 384102 96854
rect 383546 60938 383782 61174
rect 383866 60938 384102 61174
rect 383546 60618 383782 60854
rect 383866 60618 384102 60854
rect 383546 24938 383782 25174
rect 383866 24938 384102 25174
rect 383546 24618 383782 24854
rect 383866 24618 384102 24854
rect 383546 -3462 383782 -3226
rect 383866 -3462 384102 -3226
rect 383546 -3782 383782 -3546
rect 383866 -3782 384102 -3546
rect 387266 676658 387502 676894
rect 387586 676658 387822 676894
rect 387266 676338 387502 676574
rect 387586 676338 387822 676574
rect 387266 640658 387502 640894
rect 387586 640658 387822 640894
rect 387266 640338 387502 640574
rect 387586 640338 387822 640574
rect 387266 604658 387502 604894
rect 387586 604658 387822 604894
rect 387266 604338 387502 604574
rect 387586 604338 387822 604574
rect 387266 568658 387502 568894
rect 387586 568658 387822 568894
rect 387266 568338 387502 568574
rect 387586 568338 387822 568574
rect 387266 532658 387502 532894
rect 387586 532658 387822 532894
rect 387266 532338 387502 532574
rect 387586 532338 387822 532574
rect 387266 496658 387502 496894
rect 387586 496658 387822 496894
rect 387266 496338 387502 496574
rect 387586 496338 387822 496574
rect 387266 460658 387502 460894
rect 387586 460658 387822 460894
rect 387266 460338 387502 460574
rect 387586 460338 387822 460574
rect 387266 424658 387502 424894
rect 387586 424658 387822 424894
rect 387266 424338 387502 424574
rect 387586 424338 387822 424574
rect 387266 388658 387502 388894
rect 387586 388658 387822 388894
rect 387266 388338 387502 388574
rect 387586 388338 387822 388574
rect 387266 352658 387502 352894
rect 387586 352658 387822 352894
rect 387266 352338 387502 352574
rect 387586 352338 387822 352574
rect 387266 316658 387502 316894
rect 387586 316658 387822 316894
rect 387266 316338 387502 316574
rect 387586 316338 387822 316574
rect 387266 280658 387502 280894
rect 387586 280658 387822 280894
rect 387266 280338 387502 280574
rect 387586 280338 387822 280574
rect 387266 244658 387502 244894
rect 387586 244658 387822 244894
rect 387266 244338 387502 244574
rect 387586 244338 387822 244574
rect 387266 208658 387502 208894
rect 387586 208658 387822 208894
rect 387266 208338 387502 208574
rect 387586 208338 387822 208574
rect 387266 172658 387502 172894
rect 387586 172658 387822 172894
rect 387266 172338 387502 172574
rect 387586 172338 387822 172574
rect 387266 136658 387502 136894
rect 387586 136658 387822 136894
rect 387266 136338 387502 136574
rect 387586 136338 387822 136574
rect 387266 100658 387502 100894
rect 387586 100658 387822 100894
rect 387266 100338 387502 100574
rect 387586 100338 387822 100574
rect 387266 64658 387502 64894
rect 387586 64658 387822 64894
rect 387266 64338 387502 64574
rect 387586 64338 387822 64574
rect 387266 28658 387502 28894
rect 387586 28658 387822 28894
rect 387266 28338 387502 28574
rect 387586 28338 387822 28574
rect 387266 -5382 387502 -5146
rect 387586 -5382 387822 -5146
rect 387266 -5702 387502 -5466
rect 387586 -5702 387822 -5466
rect 408986 710362 409222 710598
rect 409306 710362 409542 710598
rect 408986 710042 409222 710278
rect 409306 710042 409542 710278
rect 405266 708442 405502 708678
rect 405586 708442 405822 708678
rect 405266 708122 405502 708358
rect 405586 708122 405822 708358
rect 401546 706522 401782 706758
rect 401866 706522 402102 706758
rect 401546 706202 401782 706438
rect 401866 706202 402102 706438
rect 390986 680378 391222 680614
rect 391306 680378 391542 680614
rect 390986 680058 391222 680294
rect 391306 680058 391542 680294
rect 390986 644378 391222 644614
rect 391306 644378 391542 644614
rect 390986 644058 391222 644294
rect 391306 644058 391542 644294
rect 390986 608378 391222 608614
rect 391306 608378 391542 608614
rect 390986 608058 391222 608294
rect 391306 608058 391542 608294
rect 390986 572378 391222 572614
rect 391306 572378 391542 572614
rect 390986 572058 391222 572294
rect 391306 572058 391542 572294
rect 390986 536378 391222 536614
rect 391306 536378 391542 536614
rect 390986 536058 391222 536294
rect 391306 536058 391542 536294
rect 390986 500378 391222 500614
rect 391306 500378 391542 500614
rect 390986 500058 391222 500294
rect 391306 500058 391542 500294
rect 390986 464378 391222 464614
rect 391306 464378 391542 464614
rect 390986 464058 391222 464294
rect 391306 464058 391542 464294
rect 390986 428378 391222 428614
rect 391306 428378 391542 428614
rect 390986 428058 391222 428294
rect 391306 428058 391542 428294
rect 390986 392378 391222 392614
rect 391306 392378 391542 392614
rect 390986 392058 391222 392294
rect 391306 392058 391542 392294
rect 390986 356378 391222 356614
rect 391306 356378 391542 356614
rect 390986 356058 391222 356294
rect 391306 356058 391542 356294
rect 390986 320378 391222 320614
rect 391306 320378 391542 320614
rect 390986 320058 391222 320294
rect 391306 320058 391542 320294
rect 390986 284378 391222 284614
rect 391306 284378 391542 284614
rect 390986 284058 391222 284294
rect 391306 284058 391542 284294
rect 390986 248378 391222 248614
rect 391306 248378 391542 248614
rect 390986 248058 391222 248294
rect 391306 248058 391542 248294
rect 390986 212378 391222 212614
rect 391306 212378 391542 212614
rect 390986 212058 391222 212294
rect 391306 212058 391542 212294
rect 390986 176378 391222 176614
rect 391306 176378 391542 176614
rect 390986 176058 391222 176294
rect 391306 176058 391542 176294
rect 390986 140378 391222 140614
rect 391306 140378 391542 140614
rect 390986 140058 391222 140294
rect 391306 140058 391542 140294
rect 390986 104378 391222 104614
rect 391306 104378 391542 104614
rect 390986 104058 391222 104294
rect 391306 104058 391542 104294
rect 390986 68378 391222 68614
rect 391306 68378 391542 68614
rect 390986 68058 391222 68294
rect 391306 68058 391542 68294
rect 390986 32378 391222 32614
rect 391306 32378 391542 32614
rect 390986 32058 391222 32294
rect 391306 32058 391542 32294
rect 372986 -6342 373222 -6106
rect 373306 -6342 373542 -6106
rect 372986 -6662 373222 -6426
rect 373306 -6662 373542 -6426
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 401546 618938 401782 619174
rect 401866 618938 402102 619174
rect 401546 618618 401782 618854
rect 401866 618618 402102 618854
rect 401546 582938 401782 583174
rect 401866 582938 402102 583174
rect 401546 582618 401782 582854
rect 401866 582618 402102 582854
rect 401546 546938 401782 547174
rect 401866 546938 402102 547174
rect 401546 546618 401782 546854
rect 401866 546618 402102 546854
rect 401546 510938 401782 511174
rect 401866 510938 402102 511174
rect 401546 510618 401782 510854
rect 401866 510618 402102 510854
rect 401546 474938 401782 475174
rect 401866 474938 402102 475174
rect 401546 474618 401782 474854
rect 401866 474618 402102 474854
rect 401546 438938 401782 439174
rect 401866 438938 402102 439174
rect 401546 438618 401782 438854
rect 401866 438618 402102 438854
rect 401546 402938 401782 403174
rect 401866 402938 402102 403174
rect 401546 402618 401782 402854
rect 401866 402618 402102 402854
rect 401546 366938 401782 367174
rect 401866 366938 402102 367174
rect 401546 366618 401782 366854
rect 401866 366618 402102 366854
rect 401546 330938 401782 331174
rect 401866 330938 402102 331174
rect 401546 330618 401782 330854
rect 401866 330618 402102 330854
rect 401546 294938 401782 295174
rect 401866 294938 402102 295174
rect 401546 294618 401782 294854
rect 401866 294618 402102 294854
rect 401546 258938 401782 259174
rect 401866 258938 402102 259174
rect 401546 258618 401782 258854
rect 401866 258618 402102 258854
rect 401546 222938 401782 223174
rect 401866 222938 402102 223174
rect 401546 222618 401782 222854
rect 401866 222618 402102 222854
rect 401546 186938 401782 187174
rect 401866 186938 402102 187174
rect 401546 186618 401782 186854
rect 401866 186618 402102 186854
rect 401546 150938 401782 151174
rect 401866 150938 402102 151174
rect 401546 150618 401782 150854
rect 401866 150618 402102 150854
rect 401546 114938 401782 115174
rect 401866 114938 402102 115174
rect 401546 114618 401782 114854
rect 401866 114618 402102 114854
rect 401546 78938 401782 79174
rect 401866 78938 402102 79174
rect 401546 78618 401782 78854
rect 401866 78618 402102 78854
rect 401546 42938 401782 43174
rect 401866 42938 402102 43174
rect 401546 42618 401782 42854
rect 401866 42618 402102 42854
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -2502 401782 -2266
rect 401866 -2502 402102 -2266
rect 401546 -2822 401782 -2586
rect 401866 -2822 402102 -2586
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 405266 658658 405502 658894
rect 405586 658658 405822 658894
rect 405266 658338 405502 658574
rect 405586 658338 405822 658574
rect 405266 622658 405502 622894
rect 405586 622658 405822 622894
rect 405266 622338 405502 622574
rect 405586 622338 405822 622574
rect 405266 586658 405502 586894
rect 405586 586658 405822 586894
rect 405266 586338 405502 586574
rect 405586 586338 405822 586574
rect 405266 550658 405502 550894
rect 405586 550658 405822 550894
rect 405266 550338 405502 550574
rect 405586 550338 405822 550574
rect 405266 514658 405502 514894
rect 405586 514658 405822 514894
rect 405266 514338 405502 514574
rect 405586 514338 405822 514574
rect 405266 478658 405502 478894
rect 405586 478658 405822 478894
rect 405266 478338 405502 478574
rect 405586 478338 405822 478574
rect 405266 442658 405502 442894
rect 405586 442658 405822 442894
rect 405266 442338 405502 442574
rect 405586 442338 405822 442574
rect 405266 406658 405502 406894
rect 405586 406658 405822 406894
rect 405266 406338 405502 406574
rect 405586 406338 405822 406574
rect 405266 370658 405502 370894
rect 405586 370658 405822 370894
rect 405266 370338 405502 370574
rect 405586 370338 405822 370574
rect 405266 334658 405502 334894
rect 405586 334658 405822 334894
rect 405266 334338 405502 334574
rect 405586 334338 405822 334574
rect 405266 298658 405502 298894
rect 405586 298658 405822 298894
rect 405266 298338 405502 298574
rect 405586 298338 405822 298574
rect 405266 262658 405502 262894
rect 405586 262658 405822 262894
rect 405266 262338 405502 262574
rect 405586 262338 405822 262574
rect 405266 226658 405502 226894
rect 405586 226658 405822 226894
rect 405266 226338 405502 226574
rect 405586 226338 405822 226574
rect 405266 190658 405502 190894
rect 405586 190658 405822 190894
rect 405266 190338 405502 190574
rect 405586 190338 405822 190574
rect 405266 154658 405502 154894
rect 405586 154658 405822 154894
rect 405266 154338 405502 154574
rect 405586 154338 405822 154574
rect 405266 118658 405502 118894
rect 405586 118658 405822 118894
rect 405266 118338 405502 118574
rect 405586 118338 405822 118574
rect 405266 82658 405502 82894
rect 405586 82658 405822 82894
rect 405266 82338 405502 82574
rect 405586 82338 405822 82574
rect 405266 46658 405502 46894
rect 405586 46658 405822 46894
rect 405266 46338 405502 46574
rect 405586 46338 405822 46574
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -4422 405502 -4186
rect 405586 -4422 405822 -4186
rect 405266 -4742 405502 -4506
rect 405586 -4742 405822 -4506
rect 426986 711322 427222 711558
rect 427306 711322 427542 711558
rect 426986 711002 427222 711238
rect 427306 711002 427542 711238
rect 423266 709402 423502 709638
rect 423586 709402 423822 709638
rect 423266 709082 423502 709318
rect 423586 709082 423822 709318
rect 419546 707482 419782 707718
rect 419866 707482 420102 707718
rect 419546 707162 419782 707398
rect 419866 707162 420102 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 408986 626378 409222 626614
rect 409306 626378 409542 626614
rect 408986 626058 409222 626294
rect 409306 626058 409542 626294
rect 408986 590378 409222 590614
rect 409306 590378 409542 590614
rect 408986 590058 409222 590294
rect 409306 590058 409542 590294
rect 408986 554378 409222 554614
rect 409306 554378 409542 554614
rect 408986 554058 409222 554294
rect 409306 554058 409542 554294
rect 408986 518378 409222 518614
rect 409306 518378 409542 518614
rect 408986 518058 409222 518294
rect 409306 518058 409542 518294
rect 408986 482378 409222 482614
rect 409306 482378 409542 482614
rect 408986 482058 409222 482294
rect 409306 482058 409542 482294
rect 408986 446378 409222 446614
rect 409306 446378 409542 446614
rect 408986 446058 409222 446294
rect 409306 446058 409542 446294
rect 408986 410378 409222 410614
rect 409306 410378 409542 410614
rect 408986 410058 409222 410294
rect 409306 410058 409542 410294
rect 408986 374378 409222 374614
rect 409306 374378 409542 374614
rect 408986 374058 409222 374294
rect 409306 374058 409542 374294
rect 408986 338378 409222 338614
rect 409306 338378 409542 338614
rect 408986 338058 409222 338294
rect 409306 338058 409542 338294
rect 408986 302378 409222 302614
rect 409306 302378 409542 302614
rect 408986 302058 409222 302294
rect 409306 302058 409542 302294
rect 408986 266378 409222 266614
rect 409306 266378 409542 266614
rect 408986 266058 409222 266294
rect 409306 266058 409542 266294
rect 408986 230378 409222 230614
rect 409306 230378 409542 230614
rect 408986 230058 409222 230294
rect 409306 230058 409542 230294
rect 408986 194378 409222 194614
rect 409306 194378 409542 194614
rect 408986 194058 409222 194294
rect 409306 194058 409542 194294
rect 408986 158378 409222 158614
rect 409306 158378 409542 158614
rect 408986 158058 409222 158294
rect 409306 158058 409542 158294
rect 408986 122378 409222 122614
rect 409306 122378 409542 122614
rect 408986 122058 409222 122294
rect 409306 122058 409542 122294
rect 408986 86378 409222 86614
rect 409306 86378 409542 86614
rect 408986 86058 409222 86294
rect 409306 86058 409542 86294
rect 408986 50378 409222 50614
rect 409306 50378 409542 50614
rect 408986 50058 409222 50294
rect 409306 50058 409542 50294
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 390986 -7302 391222 -7066
rect 391306 -7302 391542 -7066
rect 390986 -7622 391222 -7386
rect 391306 -7622 391542 -7386
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -1542 416062 -1306
rect 416146 -1542 416382 -1306
rect 415826 -1862 416062 -1626
rect 416146 -1862 416382 -1626
rect 419546 672938 419782 673174
rect 419866 672938 420102 673174
rect 419546 672618 419782 672854
rect 419866 672618 420102 672854
rect 419546 636938 419782 637174
rect 419866 636938 420102 637174
rect 419546 636618 419782 636854
rect 419866 636618 420102 636854
rect 419546 600938 419782 601174
rect 419866 600938 420102 601174
rect 419546 600618 419782 600854
rect 419866 600618 420102 600854
rect 419546 564938 419782 565174
rect 419866 564938 420102 565174
rect 419546 564618 419782 564854
rect 419866 564618 420102 564854
rect 419546 528938 419782 529174
rect 419866 528938 420102 529174
rect 419546 528618 419782 528854
rect 419866 528618 420102 528854
rect 419546 492938 419782 493174
rect 419866 492938 420102 493174
rect 419546 492618 419782 492854
rect 419866 492618 420102 492854
rect 419546 456938 419782 457174
rect 419866 456938 420102 457174
rect 419546 456618 419782 456854
rect 419866 456618 420102 456854
rect 419546 420938 419782 421174
rect 419866 420938 420102 421174
rect 419546 420618 419782 420854
rect 419866 420618 420102 420854
rect 419546 384938 419782 385174
rect 419866 384938 420102 385174
rect 419546 384618 419782 384854
rect 419866 384618 420102 384854
rect 419546 348938 419782 349174
rect 419866 348938 420102 349174
rect 419546 348618 419782 348854
rect 419866 348618 420102 348854
rect 419546 312938 419782 313174
rect 419866 312938 420102 313174
rect 419546 312618 419782 312854
rect 419866 312618 420102 312854
rect 419546 276938 419782 277174
rect 419866 276938 420102 277174
rect 419546 276618 419782 276854
rect 419866 276618 420102 276854
rect 419546 240938 419782 241174
rect 419866 240938 420102 241174
rect 419546 240618 419782 240854
rect 419866 240618 420102 240854
rect 419546 204938 419782 205174
rect 419866 204938 420102 205174
rect 419546 204618 419782 204854
rect 419866 204618 420102 204854
rect 419546 168938 419782 169174
rect 419866 168938 420102 169174
rect 419546 168618 419782 168854
rect 419866 168618 420102 168854
rect 419546 132938 419782 133174
rect 419866 132938 420102 133174
rect 419546 132618 419782 132854
rect 419866 132618 420102 132854
rect 419546 96938 419782 97174
rect 419866 96938 420102 97174
rect 419546 96618 419782 96854
rect 419866 96618 420102 96854
rect 419546 60938 419782 61174
rect 419866 60938 420102 61174
rect 419546 60618 419782 60854
rect 419866 60618 420102 60854
rect 419546 24938 419782 25174
rect 419866 24938 420102 25174
rect 419546 24618 419782 24854
rect 419866 24618 420102 24854
rect 419546 -3462 419782 -3226
rect 419866 -3462 420102 -3226
rect 419546 -3782 419782 -3546
rect 419866 -3782 420102 -3546
rect 423266 676658 423502 676894
rect 423586 676658 423822 676894
rect 423266 676338 423502 676574
rect 423586 676338 423822 676574
rect 423266 640658 423502 640894
rect 423586 640658 423822 640894
rect 423266 640338 423502 640574
rect 423586 640338 423822 640574
rect 423266 604658 423502 604894
rect 423586 604658 423822 604894
rect 423266 604338 423502 604574
rect 423586 604338 423822 604574
rect 423266 568658 423502 568894
rect 423586 568658 423822 568894
rect 423266 568338 423502 568574
rect 423586 568338 423822 568574
rect 423266 532658 423502 532894
rect 423586 532658 423822 532894
rect 423266 532338 423502 532574
rect 423586 532338 423822 532574
rect 423266 496658 423502 496894
rect 423586 496658 423822 496894
rect 423266 496338 423502 496574
rect 423586 496338 423822 496574
rect 423266 460658 423502 460894
rect 423586 460658 423822 460894
rect 423266 460338 423502 460574
rect 423586 460338 423822 460574
rect 423266 424658 423502 424894
rect 423586 424658 423822 424894
rect 423266 424338 423502 424574
rect 423586 424338 423822 424574
rect 423266 388658 423502 388894
rect 423586 388658 423822 388894
rect 423266 388338 423502 388574
rect 423586 388338 423822 388574
rect 423266 352658 423502 352894
rect 423586 352658 423822 352894
rect 423266 352338 423502 352574
rect 423586 352338 423822 352574
rect 423266 316658 423502 316894
rect 423586 316658 423822 316894
rect 423266 316338 423502 316574
rect 423586 316338 423822 316574
rect 423266 280658 423502 280894
rect 423586 280658 423822 280894
rect 423266 280338 423502 280574
rect 423586 280338 423822 280574
rect 423266 244658 423502 244894
rect 423586 244658 423822 244894
rect 423266 244338 423502 244574
rect 423586 244338 423822 244574
rect 423266 208658 423502 208894
rect 423586 208658 423822 208894
rect 423266 208338 423502 208574
rect 423586 208338 423822 208574
rect 423266 172658 423502 172894
rect 423586 172658 423822 172894
rect 423266 172338 423502 172574
rect 423586 172338 423822 172574
rect 423266 136658 423502 136894
rect 423586 136658 423822 136894
rect 423266 136338 423502 136574
rect 423586 136338 423822 136574
rect 423266 100658 423502 100894
rect 423586 100658 423822 100894
rect 423266 100338 423502 100574
rect 423586 100338 423822 100574
rect 423266 64658 423502 64894
rect 423586 64658 423822 64894
rect 423266 64338 423502 64574
rect 423586 64338 423822 64574
rect 423266 28658 423502 28894
rect 423586 28658 423822 28894
rect 423266 28338 423502 28574
rect 423586 28338 423822 28574
rect 423266 -5382 423502 -5146
rect 423586 -5382 423822 -5146
rect 423266 -5702 423502 -5466
rect 423586 -5702 423822 -5466
rect 444986 710362 445222 710598
rect 445306 710362 445542 710598
rect 444986 710042 445222 710278
rect 445306 710042 445542 710278
rect 441266 708442 441502 708678
rect 441586 708442 441822 708678
rect 441266 708122 441502 708358
rect 441586 708122 441822 708358
rect 437546 706522 437782 706758
rect 437866 706522 438102 706758
rect 437546 706202 437782 706438
rect 437866 706202 438102 706438
rect 426986 680378 427222 680614
rect 427306 680378 427542 680614
rect 426986 680058 427222 680294
rect 427306 680058 427542 680294
rect 426986 644378 427222 644614
rect 427306 644378 427542 644614
rect 426986 644058 427222 644294
rect 427306 644058 427542 644294
rect 426986 608378 427222 608614
rect 427306 608378 427542 608614
rect 426986 608058 427222 608294
rect 427306 608058 427542 608294
rect 426986 572378 427222 572614
rect 427306 572378 427542 572614
rect 426986 572058 427222 572294
rect 427306 572058 427542 572294
rect 426986 536378 427222 536614
rect 427306 536378 427542 536614
rect 426986 536058 427222 536294
rect 427306 536058 427542 536294
rect 426986 500378 427222 500614
rect 427306 500378 427542 500614
rect 426986 500058 427222 500294
rect 427306 500058 427542 500294
rect 426986 464378 427222 464614
rect 427306 464378 427542 464614
rect 426986 464058 427222 464294
rect 427306 464058 427542 464294
rect 426986 428378 427222 428614
rect 427306 428378 427542 428614
rect 426986 428058 427222 428294
rect 427306 428058 427542 428294
rect 426986 392378 427222 392614
rect 427306 392378 427542 392614
rect 426986 392058 427222 392294
rect 427306 392058 427542 392294
rect 426986 356378 427222 356614
rect 427306 356378 427542 356614
rect 426986 356058 427222 356294
rect 427306 356058 427542 356294
rect 426986 320378 427222 320614
rect 427306 320378 427542 320614
rect 426986 320058 427222 320294
rect 427306 320058 427542 320294
rect 426986 284378 427222 284614
rect 427306 284378 427542 284614
rect 426986 284058 427222 284294
rect 427306 284058 427542 284294
rect 426986 248378 427222 248614
rect 427306 248378 427542 248614
rect 426986 248058 427222 248294
rect 427306 248058 427542 248294
rect 426986 212378 427222 212614
rect 427306 212378 427542 212614
rect 426986 212058 427222 212294
rect 427306 212058 427542 212294
rect 426986 176378 427222 176614
rect 427306 176378 427542 176614
rect 426986 176058 427222 176294
rect 427306 176058 427542 176294
rect 426986 140378 427222 140614
rect 427306 140378 427542 140614
rect 426986 140058 427222 140294
rect 427306 140058 427542 140294
rect 426986 104378 427222 104614
rect 427306 104378 427542 104614
rect 426986 104058 427222 104294
rect 427306 104058 427542 104294
rect 426986 68378 427222 68614
rect 427306 68378 427542 68614
rect 426986 68058 427222 68294
rect 427306 68058 427542 68294
rect 426986 32378 427222 32614
rect 427306 32378 427542 32614
rect 426986 32058 427222 32294
rect 427306 32058 427542 32294
rect 408986 -6342 409222 -6106
rect 409306 -6342 409542 -6106
rect 408986 -6662 409222 -6426
rect 409306 -6662 409542 -6426
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 437546 654938 437782 655174
rect 437866 654938 438102 655174
rect 437546 654618 437782 654854
rect 437866 654618 438102 654854
rect 437546 618938 437782 619174
rect 437866 618938 438102 619174
rect 437546 618618 437782 618854
rect 437866 618618 438102 618854
rect 437546 582938 437782 583174
rect 437866 582938 438102 583174
rect 437546 582618 437782 582854
rect 437866 582618 438102 582854
rect 437546 546938 437782 547174
rect 437866 546938 438102 547174
rect 437546 546618 437782 546854
rect 437866 546618 438102 546854
rect 437546 510938 437782 511174
rect 437866 510938 438102 511174
rect 437546 510618 437782 510854
rect 437866 510618 438102 510854
rect 437546 474938 437782 475174
rect 437866 474938 438102 475174
rect 437546 474618 437782 474854
rect 437866 474618 438102 474854
rect 437546 438938 437782 439174
rect 437866 438938 438102 439174
rect 437546 438618 437782 438854
rect 437866 438618 438102 438854
rect 437546 402938 437782 403174
rect 437866 402938 438102 403174
rect 437546 402618 437782 402854
rect 437866 402618 438102 402854
rect 437546 366938 437782 367174
rect 437866 366938 438102 367174
rect 437546 366618 437782 366854
rect 437866 366618 438102 366854
rect 437546 330938 437782 331174
rect 437866 330938 438102 331174
rect 437546 330618 437782 330854
rect 437866 330618 438102 330854
rect 437546 294938 437782 295174
rect 437866 294938 438102 295174
rect 437546 294618 437782 294854
rect 437866 294618 438102 294854
rect 437546 258938 437782 259174
rect 437866 258938 438102 259174
rect 437546 258618 437782 258854
rect 437866 258618 438102 258854
rect 437546 222938 437782 223174
rect 437866 222938 438102 223174
rect 437546 222618 437782 222854
rect 437866 222618 438102 222854
rect 437546 186938 437782 187174
rect 437866 186938 438102 187174
rect 437546 186618 437782 186854
rect 437866 186618 438102 186854
rect 437546 150938 437782 151174
rect 437866 150938 438102 151174
rect 437546 150618 437782 150854
rect 437866 150618 438102 150854
rect 437546 114938 437782 115174
rect 437866 114938 438102 115174
rect 437546 114618 437782 114854
rect 437866 114618 438102 114854
rect 437546 78938 437782 79174
rect 437866 78938 438102 79174
rect 437546 78618 437782 78854
rect 437866 78618 438102 78854
rect 437546 42938 437782 43174
rect 437866 42938 438102 43174
rect 437546 42618 437782 42854
rect 437866 42618 438102 42854
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -2502 437782 -2266
rect 437866 -2502 438102 -2266
rect 437546 -2822 437782 -2586
rect 437866 -2822 438102 -2586
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 441266 658658 441502 658894
rect 441586 658658 441822 658894
rect 441266 658338 441502 658574
rect 441586 658338 441822 658574
rect 441266 622658 441502 622894
rect 441586 622658 441822 622894
rect 441266 622338 441502 622574
rect 441586 622338 441822 622574
rect 441266 586658 441502 586894
rect 441586 586658 441822 586894
rect 441266 586338 441502 586574
rect 441586 586338 441822 586574
rect 441266 550658 441502 550894
rect 441586 550658 441822 550894
rect 441266 550338 441502 550574
rect 441586 550338 441822 550574
rect 441266 514658 441502 514894
rect 441586 514658 441822 514894
rect 441266 514338 441502 514574
rect 441586 514338 441822 514574
rect 441266 478658 441502 478894
rect 441586 478658 441822 478894
rect 441266 478338 441502 478574
rect 441586 478338 441822 478574
rect 441266 442658 441502 442894
rect 441586 442658 441822 442894
rect 441266 442338 441502 442574
rect 441586 442338 441822 442574
rect 441266 406658 441502 406894
rect 441586 406658 441822 406894
rect 441266 406338 441502 406574
rect 441586 406338 441822 406574
rect 441266 370658 441502 370894
rect 441586 370658 441822 370894
rect 441266 370338 441502 370574
rect 441586 370338 441822 370574
rect 441266 334658 441502 334894
rect 441586 334658 441822 334894
rect 441266 334338 441502 334574
rect 441586 334338 441822 334574
rect 441266 298658 441502 298894
rect 441586 298658 441822 298894
rect 441266 298338 441502 298574
rect 441586 298338 441822 298574
rect 441266 262658 441502 262894
rect 441586 262658 441822 262894
rect 441266 262338 441502 262574
rect 441586 262338 441822 262574
rect 441266 226658 441502 226894
rect 441586 226658 441822 226894
rect 441266 226338 441502 226574
rect 441586 226338 441822 226574
rect 441266 190658 441502 190894
rect 441586 190658 441822 190894
rect 441266 190338 441502 190574
rect 441586 190338 441822 190574
rect 441266 154658 441502 154894
rect 441586 154658 441822 154894
rect 441266 154338 441502 154574
rect 441586 154338 441822 154574
rect 441266 118658 441502 118894
rect 441586 118658 441822 118894
rect 441266 118338 441502 118574
rect 441586 118338 441822 118574
rect 441266 82658 441502 82894
rect 441586 82658 441822 82894
rect 441266 82338 441502 82574
rect 441586 82338 441822 82574
rect 441266 46658 441502 46894
rect 441586 46658 441822 46894
rect 441266 46338 441502 46574
rect 441586 46338 441822 46574
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -4422 441502 -4186
rect 441586 -4422 441822 -4186
rect 441266 -4742 441502 -4506
rect 441586 -4742 441822 -4506
rect 462986 711322 463222 711558
rect 463306 711322 463542 711558
rect 462986 711002 463222 711238
rect 463306 711002 463542 711238
rect 459266 709402 459502 709638
rect 459586 709402 459822 709638
rect 459266 709082 459502 709318
rect 459586 709082 459822 709318
rect 455546 707482 455782 707718
rect 455866 707482 456102 707718
rect 455546 707162 455782 707398
rect 455866 707162 456102 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 444986 662378 445222 662614
rect 445306 662378 445542 662614
rect 444986 662058 445222 662294
rect 445306 662058 445542 662294
rect 444986 626378 445222 626614
rect 445306 626378 445542 626614
rect 444986 626058 445222 626294
rect 445306 626058 445542 626294
rect 444986 590378 445222 590614
rect 445306 590378 445542 590614
rect 444986 590058 445222 590294
rect 445306 590058 445542 590294
rect 444986 554378 445222 554614
rect 445306 554378 445542 554614
rect 444986 554058 445222 554294
rect 445306 554058 445542 554294
rect 444986 518378 445222 518614
rect 445306 518378 445542 518614
rect 444986 518058 445222 518294
rect 445306 518058 445542 518294
rect 444986 482378 445222 482614
rect 445306 482378 445542 482614
rect 444986 482058 445222 482294
rect 445306 482058 445542 482294
rect 444986 446378 445222 446614
rect 445306 446378 445542 446614
rect 444986 446058 445222 446294
rect 445306 446058 445542 446294
rect 444986 410378 445222 410614
rect 445306 410378 445542 410614
rect 444986 410058 445222 410294
rect 445306 410058 445542 410294
rect 444986 374378 445222 374614
rect 445306 374378 445542 374614
rect 444986 374058 445222 374294
rect 445306 374058 445542 374294
rect 444986 338378 445222 338614
rect 445306 338378 445542 338614
rect 444986 338058 445222 338294
rect 445306 338058 445542 338294
rect 444986 302378 445222 302614
rect 445306 302378 445542 302614
rect 444986 302058 445222 302294
rect 445306 302058 445542 302294
rect 444986 266378 445222 266614
rect 445306 266378 445542 266614
rect 444986 266058 445222 266294
rect 445306 266058 445542 266294
rect 444986 230378 445222 230614
rect 445306 230378 445542 230614
rect 444986 230058 445222 230294
rect 445306 230058 445542 230294
rect 444986 194378 445222 194614
rect 445306 194378 445542 194614
rect 444986 194058 445222 194294
rect 445306 194058 445542 194294
rect 444986 158378 445222 158614
rect 445306 158378 445542 158614
rect 444986 158058 445222 158294
rect 445306 158058 445542 158294
rect 444986 122378 445222 122614
rect 445306 122378 445542 122614
rect 444986 122058 445222 122294
rect 445306 122058 445542 122294
rect 444986 86378 445222 86614
rect 445306 86378 445542 86614
rect 444986 86058 445222 86294
rect 445306 86058 445542 86294
rect 444986 50378 445222 50614
rect 445306 50378 445542 50614
rect 444986 50058 445222 50294
rect 445306 50058 445542 50294
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 426986 -7302 427222 -7066
rect 427306 -7302 427542 -7066
rect 426986 -7622 427222 -7386
rect 427306 -7622 427542 -7386
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -1542 452062 -1306
rect 452146 -1542 452382 -1306
rect 451826 -1862 452062 -1626
rect 452146 -1862 452382 -1626
rect 455546 672938 455782 673174
rect 455866 672938 456102 673174
rect 455546 672618 455782 672854
rect 455866 672618 456102 672854
rect 455546 636938 455782 637174
rect 455866 636938 456102 637174
rect 455546 636618 455782 636854
rect 455866 636618 456102 636854
rect 455546 600938 455782 601174
rect 455866 600938 456102 601174
rect 455546 600618 455782 600854
rect 455866 600618 456102 600854
rect 455546 564938 455782 565174
rect 455866 564938 456102 565174
rect 455546 564618 455782 564854
rect 455866 564618 456102 564854
rect 455546 528938 455782 529174
rect 455866 528938 456102 529174
rect 455546 528618 455782 528854
rect 455866 528618 456102 528854
rect 455546 492938 455782 493174
rect 455866 492938 456102 493174
rect 455546 492618 455782 492854
rect 455866 492618 456102 492854
rect 455546 456938 455782 457174
rect 455866 456938 456102 457174
rect 455546 456618 455782 456854
rect 455866 456618 456102 456854
rect 455546 420938 455782 421174
rect 455866 420938 456102 421174
rect 455546 420618 455782 420854
rect 455866 420618 456102 420854
rect 455546 384938 455782 385174
rect 455866 384938 456102 385174
rect 455546 384618 455782 384854
rect 455866 384618 456102 384854
rect 455546 348938 455782 349174
rect 455866 348938 456102 349174
rect 455546 348618 455782 348854
rect 455866 348618 456102 348854
rect 455546 312938 455782 313174
rect 455866 312938 456102 313174
rect 455546 312618 455782 312854
rect 455866 312618 456102 312854
rect 455546 276938 455782 277174
rect 455866 276938 456102 277174
rect 455546 276618 455782 276854
rect 455866 276618 456102 276854
rect 455546 240938 455782 241174
rect 455866 240938 456102 241174
rect 455546 240618 455782 240854
rect 455866 240618 456102 240854
rect 455546 204938 455782 205174
rect 455866 204938 456102 205174
rect 455546 204618 455782 204854
rect 455866 204618 456102 204854
rect 455546 168938 455782 169174
rect 455866 168938 456102 169174
rect 455546 168618 455782 168854
rect 455866 168618 456102 168854
rect 455546 132938 455782 133174
rect 455866 132938 456102 133174
rect 455546 132618 455782 132854
rect 455866 132618 456102 132854
rect 455546 96938 455782 97174
rect 455866 96938 456102 97174
rect 455546 96618 455782 96854
rect 455866 96618 456102 96854
rect 455546 60938 455782 61174
rect 455866 60938 456102 61174
rect 455546 60618 455782 60854
rect 455866 60618 456102 60854
rect 455546 24938 455782 25174
rect 455866 24938 456102 25174
rect 455546 24618 455782 24854
rect 455866 24618 456102 24854
rect 455546 -3462 455782 -3226
rect 455866 -3462 456102 -3226
rect 455546 -3782 455782 -3546
rect 455866 -3782 456102 -3546
rect 459266 676658 459502 676894
rect 459586 676658 459822 676894
rect 459266 676338 459502 676574
rect 459586 676338 459822 676574
rect 459266 640658 459502 640894
rect 459586 640658 459822 640894
rect 459266 640338 459502 640574
rect 459586 640338 459822 640574
rect 459266 604658 459502 604894
rect 459586 604658 459822 604894
rect 459266 604338 459502 604574
rect 459586 604338 459822 604574
rect 459266 568658 459502 568894
rect 459586 568658 459822 568894
rect 459266 568338 459502 568574
rect 459586 568338 459822 568574
rect 459266 532658 459502 532894
rect 459586 532658 459822 532894
rect 459266 532338 459502 532574
rect 459586 532338 459822 532574
rect 459266 496658 459502 496894
rect 459586 496658 459822 496894
rect 459266 496338 459502 496574
rect 459586 496338 459822 496574
rect 459266 460658 459502 460894
rect 459586 460658 459822 460894
rect 459266 460338 459502 460574
rect 459586 460338 459822 460574
rect 459266 424658 459502 424894
rect 459586 424658 459822 424894
rect 459266 424338 459502 424574
rect 459586 424338 459822 424574
rect 459266 388658 459502 388894
rect 459586 388658 459822 388894
rect 459266 388338 459502 388574
rect 459586 388338 459822 388574
rect 459266 352658 459502 352894
rect 459586 352658 459822 352894
rect 459266 352338 459502 352574
rect 459586 352338 459822 352574
rect 459266 316658 459502 316894
rect 459586 316658 459822 316894
rect 459266 316338 459502 316574
rect 459586 316338 459822 316574
rect 459266 280658 459502 280894
rect 459586 280658 459822 280894
rect 459266 280338 459502 280574
rect 459586 280338 459822 280574
rect 459266 244658 459502 244894
rect 459586 244658 459822 244894
rect 459266 244338 459502 244574
rect 459586 244338 459822 244574
rect 459266 208658 459502 208894
rect 459586 208658 459822 208894
rect 459266 208338 459502 208574
rect 459586 208338 459822 208574
rect 459266 172658 459502 172894
rect 459586 172658 459822 172894
rect 459266 172338 459502 172574
rect 459586 172338 459822 172574
rect 459266 136658 459502 136894
rect 459586 136658 459822 136894
rect 459266 136338 459502 136574
rect 459586 136338 459822 136574
rect 459266 100658 459502 100894
rect 459586 100658 459822 100894
rect 459266 100338 459502 100574
rect 459586 100338 459822 100574
rect 459266 64658 459502 64894
rect 459586 64658 459822 64894
rect 459266 64338 459502 64574
rect 459586 64338 459822 64574
rect 459266 28658 459502 28894
rect 459586 28658 459822 28894
rect 459266 28338 459502 28574
rect 459586 28338 459822 28574
rect 459266 -5382 459502 -5146
rect 459586 -5382 459822 -5146
rect 459266 -5702 459502 -5466
rect 459586 -5702 459822 -5466
rect 480986 710362 481222 710598
rect 481306 710362 481542 710598
rect 480986 710042 481222 710278
rect 481306 710042 481542 710278
rect 477266 708442 477502 708678
rect 477586 708442 477822 708678
rect 477266 708122 477502 708358
rect 477586 708122 477822 708358
rect 473546 706522 473782 706758
rect 473866 706522 474102 706758
rect 473546 706202 473782 706438
rect 473866 706202 474102 706438
rect 462986 680378 463222 680614
rect 463306 680378 463542 680614
rect 462986 680058 463222 680294
rect 463306 680058 463542 680294
rect 462986 644378 463222 644614
rect 463306 644378 463542 644614
rect 462986 644058 463222 644294
rect 463306 644058 463542 644294
rect 462986 608378 463222 608614
rect 463306 608378 463542 608614
rect 462986 608058 463222 608294
rect 463306 608058 463542 608294
rect 462986 572378 463222 572614
rect 463306 572378 463542 572614
rect 462986 572058 463222 572294
rect 463306 572058 463542 572294
rect 462986 536378 463222 536614
rect 463306 536378 463542 536614
rect 462986 536058 463222 536294
rect 463306 536058 463542 536294
rect 462986 500378 463222 500614
rect 463306 500378 463542 500614
rect 462986 500058 463222 500294
rect 463306 500058 463542 500294
rect 462986 464378 463222 464614
rect 463306 464378 463542 464614
rect 462986 464058 463222 464294
rect 463306 464058 463542 464294
rect 462986 428378 463222 428614
rect 463306 428378 463542 428614
rect 462986 428058 463222 428294
rect 463306 428058 463542 428294
rect 462986 392378 463222 392614
rect 463306 392378 463542 392614
rect 462986 392058 463222 392294
rect 463306 392058 463542 392294
rect 462986 356378 463222 356614
rect 463306 356378 463542 356614
rect 462986 356058 463222 356294
rect 463306 356058 463542 356294
rect 462986 320378 463222 320614
rect 463306 320378 463542 320614
rect 462986 320058 463222 320294
rect 463306 320058 463542 320294
rect 462986 284378 463222 284614
rect 463306 284378 463542 284614
rect 462986 284058 463222 284294
rect 463306 284058 463542 284294
rect 462986 248378 463222 248614
rect 463306 248378 463542 248614
rect 462986 248058 463222 248294
rect 463306 248058 463542 248294
rect 462986 212378 463222 212614
rect 463306 212378 463542 212614
rect 462986 212058 463222 212294
rect 463306 212058 463542 212294
rect 462986 176378 463222 176614
rect 463306 176378 463542 176614
rect 462986 176058 463222 176294
rect 463306 176058 463542 176294
rect 462986 140378 463222 140614
rect 463306 140378 463542 140614
rect 462986 140058 463222 140294
rect 463306 140058 463542 140294
rect 462986 104378 463222 104614
rect 463306 104378 463542 104614
rect 462986 104058 463222 104294
rect 463306 104058 463542 104294
rect 462986 68378 463222 68614
rect 463306 68378 463542 68614
rect 462986 68058 463222 68294
rect 463306 68058 463542 68294
rect 462986 32378 463222 32614
rect 463306 32378 463542 32614
rect 462986 32058 463222 32294
rect 463306 32058 463542 32294
rect 444986 -6342 445222 -6106
rect 445306 -6342 445542 -6106
rect 444986 -6662 445222 -6426
rect 445306 -6662 445542 -6426
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 473546 654938 473782 655174
rect 473866 654938 474102 655174
rect 473546 654618 473782 654854
rect 473866 654618 474102 654854
rect 473546 618938 473782 619174
rect 473866 618938 474102 619174
rect 473546 618618 473782 618854
rect 473866 618618 474102 618854
rect 473546 582938 473782 583174
rect 473866 582938 474102 583174
rect 473546 582618 473782 582854
rect 473866 582618 474102 582854
rect 473546 546938 473782 547174
rect 473866 546938 474102 547174
rect 473546 546618 473782 546854
rect 473866 546618 474102 546854
rect 473546 510938 473782 511174
rect 473866 510938 474102 511174
rect 473546 510618 473782 510854
rect 473866 510618 474102 510854
rect 473546 474938 473782 475174
rect 473866 474938 474102 475174
rect 473546 474618 473782 474854
rect 473866 474618 474102 474854
rect 473546 438938 473782 439174
rect 473866 438938 474102 439174
rect 473546 438618 473782 438854
rect 473866 438618 474102 438854
rect 473546 402938 473782 403174
rect 473866 402938 474102 403174
rect 473546 402618 473782 402854
rect 473866 402618 474102 402854
rect 473546 366938 473782 367174
rect 473866 366938 474102 367174
rect 473546 366618 473782 366854
rect 473866 366618 474102 366854
rect 473546 330938 473782 331174
rect 473866 330938 474102 331174
rect 473546 330618 473782 330854
rect 473866 330618 474102 330854
rect 473546 294938 473782 295174
rect 473866 294938 474102 295174
rect 473546 294618 473782 294854
rect 473866 294618 474102 294854
rect 473546 258938 473782 259174
rect 473866 258938 474102 259174
rect 473546 258618 473782 258854
rect 473866 258618 474102 258854
rect 473546 222938 473782 223174
rect 473866 222938 474102 223174
rect 473546 222618 473782 222854
rect 473866 222618 474102 222854
rect 473546 186938 473782 187174
rect 473866 186938 474102 187174
rect 473546 186618 473782 186854
rect 473866 186618 474102 186854
rect 473546 150938 473782 151174
rect 473866 150938 474102 151174
rect 473546 150618 473782 150854
rect 473866 150618 474102 150854
rect 473546 114938 473782 115174
rect 473866 114938 474102 115174
rect 473546 114618 473782 114854
rect 473866 114618 474102 114854
rect 473546 78938 473782 79174
rect 473866 78938 474102 79174
rect 473546 78618 473782 78854
rect 473866 78618 474102 78854
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -2502 473782 -2266
rect 473866 -2502 474102 -2266
rect 473546 -2822 473782 -2586
rect 473866 -2822 474102 -2586
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 477266 658658 477502 658894
rect 477586 658658 477822 658894
rect 477266 658338 477502 658574
rect 477586 658338 477822 658574
rect 477266 622658 477502 622894
rect 477586 622658 477822 622894
rect 477266 622338 477502 622574
rect 477586 622338 477822 622574
rect 477266 586658 477502 586894
rect 477586 586658 477822 586894
rect 477266 586338 477502 586574
rect 477586 586338 477822 586574
rect 477266 550658 477502 550894
rect 477586 550658 477822 550894
rect 477266 550338 477502 550574
rect 477586 550338 477822 550574
rect 477266 514658 477502 514894
rect 477586 514658 477822 514894
rect 477266 514338 477502 514574
rect 477586 514338 477822 514574
rect 477266 478658 477502 478894
rect 477586 478658 477822 478894
rect 477266 478338 477502 478574
rect 477586 478338 477822 478574
rect 477266 442658 477502 442894
rect 477586 442658 477822 442894
rect 477266 442338 477502 442574
rect 477586 442338 477822 442574
rect 477266 406658 477502 406894
rect 477586 406658 477822 406894
rect 477266 406338 477502 406574
rect 477586 406338 477822 406574
rect 477266 370658 477502 370894
rect 477586 370658 477822 370894
rect 477266 370338 477502 370574
rect 477586 370338 477822 370574
rect 477266 334658 477502 334894
rect 477586 334658 477822 334894
rect 477266 334338 477502 334574
rect 477586 334338 477822 334574
rect 477266 298658 477502 298894
rect 477586 298658 477822 298894
rect 477266 298338 477502 298574
rect 477586 298338 477822 298574
rect 477266 262658 477502 262894
rect 477586 262658 477822 262894
rect 477266 262338 477502 262574
rect 477586 262338 477822 262574
rect 477266 226658 477502 226894
rect 477586 226658 477822 226894
rect 477266 226338 477502 226574
rect 477586 226338 477822 226574
rect 477266 190658 477502 190894
rect 477586 190658 477822 190894
rect 477266 190338 477502 190574
rect 477586 190338 477822 190574
rect 477266 154658 477502 154894
rect 477586 154658 477822 154894
rect 477266 154338 477502 154574
rect 477586 154338 477822 154574
rect 477266 118658 477502 118894
rect 477586 118658 477822 118894
rect 477266 118338 477502 118574
rect 477586 118338 477822 118574
rect 477266 82658 477502 82894
rect 477586 82658 477822 82894
rect 477266 82338 477502 82574
rect 477586 82338 477822 82574
rect 477266 46658 477502 46894
rect 477586 46658 477822 46894
rect 477266 46338 477502 46574
rect 477586 46338 477822 46574
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -4422 477502 -4186
rect 477586 -4422 477822 -4186
rect 477266 -4742 477502 -4506
rect 477586 -4742 477822 -4506
rect 498986 711322 499222 711558
rect 499306 711322 499542 711558
rect 498986 711002 499222 711238
rect 499306 711002 499542 711238
rect 495266 709402 495502 709638
rect 495586 709402 495822 709638
rect 495266 709082 495502 709318
rect 495586 709082 495822 709318
rect 491546 707482 491782 707718
rect 491866 707482 492102 707718
rect 491546 707162 491782 707398
rect 491866 707162 492102 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 480986 662378 481222 662614
rect 481306 662378 481542 662614
rect 480986 662058 481222 662294
rect 481306 662058 481542 662294
rect 480986 626378 481222 626614
rect 481306 626378 481542 626614
rect 480986 626058 481222 626294
rect 481306 626058 481542 626294
rect 480986 590378 481222 590614
rect 481306 590378 481542 590614
rect 480986 590058 481222 590294
rect 481306 590058 481542 590294
rect 480986 554378 481222 554614
rect 481306 554378 481542 554614
rect 480986 554058 481222 554294
rect 481306 554058 481542 554294
rect 480986 518378 481222 518614
rect 481306 518378 481542 518614
rect 480986 518058 481222 518294
rect 481306 518058 481542 518294
rect 480986 482378 481222 482614
rect 481306 482378 481542 482614
rect 480986 482058 481222 482294
rect 481306 482058 481542 482294
rect 480986 446378 481222 446614
rect 481306 446378 481542 446614
rect 480986 446058 481222 446294
rect 481306 446058 481542 446294
rect 480986 410378 481222 410614
rect 481306 410378 481542 410614
rect 480986 410058 481222 410294
rect 481306 410058 481542 410294
rect 480986 374378 481222 374614
rect 481306 374378 481542 374614
rect 480986 374058 481222 374294
rect 481306 374058 481542 374294
rect 480986 338378 481222 338614
rect 481306 338378 481542 338614
rect 480986 338058 481222 338294
rect 481306 338058 481542 338294
rect 480986 302378 481222 302614
rect 481306 302378 481542 302614
rect 480986 302058 481222 302294
rect 481306 302058 481542 302294
rect 480986 266378 481222 266614
rect 481306 266378 481542 266614
rect 480986 266058 481222 266294
rect 481306 266058 481542 266294
rect 480986 230378 481222 230614
rect 481306 230378 481542 230614
rect 480986 230058 481222 230294
rect 481306 230058 481542 230294
rect 480986 194378 481222 194614
rect 481306 194378 481542 194614
rect 480986 194058 481222 194294
rect 481306 194058 481542 194294
rect 480986 158378 481222 158614
rect 481306 158378 481542 158614
rect 480986 158058 481222 158294
rect 481306 158058 481542 158294
rect 480986 122378 481222 122614
rect 481306 122378 481542 122614
rect 480986 122058 481222 122294
rect 481306 122058 481542 122294
rect 480986 86378 481222 86614
rect 481306 86378 481542 86614
rect 480986 86058 481222 86294
rect 481306 86058 481542 86294
rect 480986 50378 481222 50614
rect 481306 50378 481542 50614
rect 480986 50058 481222 50294
rect 481306 50058 481542 50294
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 462986 -7302 463222 -7066
rect 463306 -7302 463542 -7066
rect 462986 -7622 463222 -7386
rect 463306 -7622 463542 -7386
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -1542 488062 -1306
rect 488146 -1542 488382 -1306
rect 487826 -1862 488062 -1626
rect 488146 -1862 488382 -1626
rect 491546 672938 491782 673174
rect 491866 672938 492102 673174
rect 491546 672618 491782 672854
rect 491866 672618 492102 672854
rect 491546 636938 491782 637174
rect 491866 636938 492102 637174
rect 491546 636618 491782 636854
rect 491866 636618 492102 636854
rect 491546 600938 491782 601174
rect 491866 600938 492102 601174
rect 491546 600618 491782 600854
rect 491866 600618 492102 600854
rect 491546 564938 491782 565174
rect 491866 564938 492102 565174
rect 491546 564618 491782 564854
rect 491866 564618 492102 564854
rect 491546 528938 491782 529174
rect 491866 528938 492102 529174
rect 491546 528618 491782 528854
rect 491866 528618 492102 528854
rect 491546 492938 491782 493174
rect 491866 492938 492102 493174
rect 491546 492618 491782 492854
rect 491866 492618 492102 492854
rect 491546 456938 491782 457174
rect 491866 456938 492102 457174
rect 491546 456618 491782 456854
rect 491866 456618 492102 456854
rect 491546 420938 491782 421174
rect 491866 420938 492102 421174
rect 491546 420618 491782 420854
rect 491866 420618 492102 420854
rect 491546 384938 491782 385174
rect 491866 384938 492102 385174
rect 491546 384618 491782 384854
rect 491866 384618 492102 384854
rect 491546 348938 491782 349174
rect 491866 348938 492102 349174
rect 491546 348618 491782 348854
rect 491866 348618 492102 348854
rect 491546 312938 491782 313174
rect 491866 312938 492102 313174
rect 491546 312618 491782 312854
rect 491866 312618 492102 312854
rect 491546 276938 491782 277174
rect 491866 276938 492102 277174
rect 491546 276618 491782 276854
rect 491866 276618 492102 276854
rect 491546 240938 491782 241174
rect 491866 240938 492102 241174
rect 491546 240618 491782 240854
rect 491866 240618 492102 240854
rect 491546 204938 491782 205174
rect 491866 204938 492102 205174
rect 491546 204618 491782 204854
rect 491866 204618 492102 204854
rect 491546 168938 491782 169174
rect 491866 168938 492102 169174
rect 491546 168618 491782 168854
rect 491866 168618 492102 168854
rect 491546 132938 491782 133174
rect 491866 132938 492102 133174
rect 491546 132618 491782 132854
rect 491866 132618 492102 132854
rect 491546 96938 491782 97174
rect 491866 96938 492102 97174
rect 491546 96618 491782 96854
rect 491866 96618 492102 96854
rect 491546 60938 491782 61174
rect 491866 60938 492102 61174
rect 491546 60618 491782 60854
rect 491866 60618 492102 60854
rect 491546 24938 491782 25174
rect 491866 24938 492102 25174
rect 491546 24618 491782 24854
rect 491866 24618 492102 24854
rect 491546 -3462 491782 -3226
rect 491866 -3462 492102 -3226
rect 491546 -3782 491782 -3546
rect 491866 -3782 492102 -3546
rect 495266 676658 495502 676894
rect 495586 676658 495822 676894
rect 495266 676338 495502 676574
rect 495586 676338 495822 676574
rect 495266 640658 495502 640894
rect 495586 640658 495822 640894
rect 495266 640338 495502 640574
rect 495586 640338 495822 640574
rect 495266 604658 495502 604894
rect 495586 604658 495822 604894
rect 495266 604338 495502 604574
rect 495586 604338 495822 604574
rect 495266 568658 495502 568894
rect 495586 568658 495822 568894
rect 495266 568338 495502 568574
rect 495586 568338 495822 568574
rect 495266 532658 495502 532894
rect 495586 532658 495822 532894
rect 495266 532338 495502 532574
rect 495586 532338 495822 532574
rect 495266 496658 495502 496894
rect 495586 496658 495822 496894
rect 495266 496338 495502 496574
rect 495586 496338 495822 496574
rect 495266 460658 495502 460894
rect 495586 460658 495822 460894
rect 495266 460338 495502 460574
rect 495586 460338 495822 460574
rect 495266 424658 495502 424894
rect 495586 424658 495822 424894
rect 495266 424338 495502 424574
rect 495586 424338 495822 424574
rect 495266 388658 495502 388894
rect 495586 388658 495822 388894
rect 495266 388338 495502 388574
rect 495586 388338 495822 388574
rect 495266 352658 495502 352894
rect 495586 352658 495822 352894
rect 495266 352338 495502 352574
rect 495586 352338 495822 352574
rect 495266 316658 495502 316894
rect 495586 316658 495822 316894
rect 495266 316338 495502 316574
rect 495586 316338 495822 316574
rect 495266 280658 495502 280894
rect 495586 280658 495822 280894
rect 495266 280338 495502 280574
rect 495586 280338 495822 280574
rect 495266 244658 495502 244894
rect 495586 244658 495822 244894
rect 495266 244338 495502 244574
rect 495586 244338 495822 244574
rect 495266 208658 495502 208894
rect 495586 208658 495822 208894
rect 495266 208338 495502 208574
rect 495586 208338 495822 208574
rect 495266 172658 495502 172894
rect 495586 172658 495822 172894
rect 495266 172338 495502 172574
rect 495586 172338 495822 172574
rect 495266 136658 495502 136894
rect 495586 136658 495822 136894
rect 495266 136338 495502 136574
rect 495586 136338 495822 136574
rect 495266 100658 495502 100894
rect 495586 100658 495822 100894
rect 495266 100338 495502 100574
rect 495586 100338 495822 100574
rect 495266 64658 495502 64894
rect 495586 64658 495822 64894
rect 495266 64338 495502 64574
rect 495586 64338 495822 64574
rect 495266 28658 495502 28894
rect 495586 28658 495822 28894
rect 495266 28338 495502 28574
rect 495586 28338 495822 28574
rect 495266 -5382 495502 -5146
rect 495586 -5382 495822 -5146
rect 495266 -5702 495502 -5466
rect 495586 -5702 495822 -5466
rect 516986 710362 517222 710598
rect 517306 710362 517542 710598
rect 516986 710042 517222 710278
rect 517306 710042 517542 710278
rect 513266 708442 513502 708678
rect 513586 708442 513822 708678
rect 513266 708122 513502 708358
rect 513586 708122 513822 708358
rect 509546 706522 509782 706758
rect 509866 706522 510102 706758
rect 509546 706202 509782 706438
rect 509866 706202 510102 706438
rect 498986 680378 499222 680614
rect 499306 680378 499542 680614
rect 498986 680058 499222 680294
rect 499306 680058 499542 680294
rect 498986 644378 499222 644614
rect 499306 644378 499542 644614
rect 498986 644058 499222 644294
rect 499306 644058 499542 644294
rect 498986 608378 499222 608614
rect 499306 608378 499542 608614
rect 498986 608058 499222 608294
rect 499306 608058 499542 608294
rect 498986 572378 499222 572614
rect 499306 572378 499542 572614
rect 498986 572058 499222 572294
rect 499306 572058 499542 572294
rect 498986 536378 499222 536614
rect 499306 536378 499542 536614
rect 498986 536058 499222 536294
rect 499306 536058 499542 536294
rect 498986 500378 499222 500614
rect 499306 500378 499542 500614
rect 498986 500058 499222 500294
rect 499306 500058 499542 500294
rect 498986 464378 499222 464614
rect 499306 464378 499542 464614
rect 498986 464058 499222 464294
rect 499306 464058 499542 464294
rect 498986 428378 499222 428614
rect 499306 428378 499542 428614
rect 498986 428058 499222 428294
rect 499306 428058 499542 428294
rect 498986 392378 499222 392614
rect 499306 392378 499542 392614
rect 498986 392058 499222 392294
rect 499306 392058 499542 392294
rect 498986 356378 499222 356614
rect 499306 356378 499542 356614
rect 498986 356058 499222 356294
rect 499306 356058 499542 356294
rect 498986 320378 499222 320614
rect 499306 320378 499542 320614
rect 498986 320058 499222 320294
rect 499306 320058 499542 320294
rect 498986 284378 499222 284614
rect 499306 284378 499542 284614
rect 498986 284058 499222 284294
rect 499306 284058 499542 284294
rect 498986 248378 499222 248614
rect 499306 248378 499542 248614
rect 498986 248058 499222 248294
rect 499306 248058 499542 248294
rect 498986 212378 499222 212614
rect 499306 212378 499542 212614
rect 498986 212058 499222 212294
rect 499306 212058 499542 212294
rect 498986 176378 499222 176614
rect 499306 176378 499542 176614
rect 498986 176058 499222 176294
rect 499306 176058 499542 176294
rect 498986 140378 499222 140614
rect 499306 140378 499542 140614
rect 498986 140058 499222 140294
rect 499306 140058 499542 140294
rect 498986 104378 499222 104614
rect 499306 104378 499542 104614
rect 498986 104058 499222 104294
rect 499306 104058 499542 104294
rect 498986 68378 499222 68614
rect 499306 68378 499542 68614
rect 498986 68058 499222 68294
rect 499306 68058 499542 68294
rect 498986 32378 499222 32614
rect 499306 32378 499542 32614
rect 498986 32058 499222 32294
rect 499306 32058 499542 32294
rect 480986 -6342 481222 -6106
rect 481306 -6342 481542 -6106
rect 480986 -6662 481222 -6426
rect 481306 -6662 481542 -6426
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 509546 654938 509782 655174
rect 509866 654938 510102 655174
rect 509546 654618 509782 654854
rect 509866 654618 510102 654854
rect 509546 618938 509782 619174
rect 509866 618938 510102 619174
rect 509546 618618 509782 618854
rect 509866 618618 510102 618854
rect 509546 582938 509782 583174
rect 509866 582938 510102 583174
rect 509546 582618 509782 582854
rect 509866 582618 510102 582854
rect 509546 546938 509782 547174
rect 509866 546938 510102 547174
rect 509546 546618 509782 546854
rect 509866 546618 510102 546854
rect 509546 510938 509782 511174
rect 509866 510938 510102 511174
rect 509546 510618 509782 510854
rect 509866 510618 510102 510854
rect 509546 474938 509782 475174
rect 509866 474938 510102 475174
rect 509546 474618 509782 474854
rect 509866 474618 510102 474854
rect 509546 438938 509782 439174
rect 509866 438938 510102 439174
rect 509546 438618 509782 438854
rect 509866 438618 510102 438854
rect 509546 402938 509782 403174
rect 509866 402938 510102 403174
rect 509546 402618 509782 402854
rect 509866 402618 510102 402854
rect 509546 366938 509782 367174
rect 509866 366938 510102 367174
rect 509546 366618 509782 366854
rect 509866 366618 510102 366854
rect 509546 330938 509782 331174
rect 509866 330938 510102 331174
rect 509546 330618 509782 330854
rect 509866 330618 510102 330854
rect 509546 294938 509782 295174
rect 509866 294938 510102 295174
rect 509546 294618 509782 294854
rect 509866 294618 510102 294854
rect 509546 258938 509782 259174
rect 509866 258938 510102 259174
rect 509546 258618 509782 258854
rect 509866 258618 510102 258854
rect 509546 222938 509782 223174
rect 509866 222938 510102 223174
rect 509546 222618 509782 222854
rect 509866 222618 510102 222854
rect 509546 186938 509782 187174
rect 509866 186938 510102 187174
rect 509546 186618 509782 186854
rect 509866 186618 510102 186854
rect 509546 150938 509782 151174
rect 509866 150938 510102 151174
rect 509546 150618 509782 150854
rect 509866 150618 510102 150854
rect 509546 114938 509782 115174
rect 509866 114938 510102 115174
rect 509546 114618 509782 114854
rect 509866 114618 510102 114854
rect 509546 78938 509782 79174
rect 509866 78938 510102 79174
rect 509546 78618 509782 78854
rect 509866 78618 510102 78854
rect 509546 42938 509782 43174
rect 509866 42938 510102 43174
rect 509546 42618 509782 42854
rect 509866 42618 510102 42854
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -2502 509782 -2266
rect 509866 -2502 510102 -2266
rect 509546 -2822 509782 -2586
rect 509866 -2822 510102 -2586
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 513266 658658 513502 658894
rect 513586 658658 513822 658894
rect 513266 658338 513502 658574
rect 513586 658338 513822 658574
rect 513266 622658 513502 622894
rect 513586 622658 513822 622894
rect 513266 622338 513502 622574
rect 513586 622338 513822 622574
rect 513266 586658 513502 586894
rect 513586 586658 513822 586894
rect 513266 586338 513502 586574
rect 513586 586338 513822 586574
rect 513266 550658 513502 550894
rect 513586 550658 513822 550894
rect 513266 550338 513502 550574
rect 513586 550338 513822 550574
rect 513266 514658 513502 514894
rect 513586 514658 513822 514894
rect 513266 514338 513502 514574
rect 513586 514338 513822 514574
rect 513266 478658 513502 478894
rect 513586 478658 513822 478894
rect 513266 478338 513502 478574
rect 513586 478338 513822 478574
rect 513266 442658 513502 442894
rect 513586 442658 513822 442894
rect 513266 442338 513502 442574
rect 513586 442338 513822 442574
rect 513266 406658 513502 406894
rect 513586 406658 513822 406894
rect 513266 406338 513502 406574
rect 513586 406338 513822 406574
rect 513266 370658 513502 370894
rect 513586 370658 513822 370894
rect 513266 370338 513502 370574
rect 513586 370338 513822 370574
rect 513266 334658 513502 334894
rect 513586 334658 513822 334894
rect 513266 334338 513502 334574
rect 513586 334338 513822 334574
rect 513266 298658 513502 298894
rect 513586 298658 513822 298894
rect 513266 298338 513502 298574
rect 513586 298338 513822 298574
rect 513266 262658 513502 262894
rect 513586 262658 513822 262894
rect 513266 262338 513502 262574
rect 513586 262338 513822 262574
rect 513266 226658 513502 226894
rect 513586 226658 513822 226894
rect 513266 226338 513502 226574
rect 513586 226338 513822 226574
rect 513266 190658 513502 190894
rect 513586 190658 513822 190894
rect 513266 190338 513502 190574
rect 513586 190338 513822 190574
rect 513266 154658 513502 154894
rect 513586 154658 513822 154894
rect 513266 154338 513502 154574
rect 513586 154338 513822 154574
rect 513266 118658 513502 118894
rect 513586 118658 513822 118894
rect 513266 118338 513502 118574
rect 513586 118338 513822 118574
rect 513266 82658 513502 82894
rect 513586 82658 513822 82894
rect 513266 82338 513502 82574
rect 513586 82338 513822 82574
rect 513266 46658 513502 46894
rect 513586 46658 513822 46894
rect 513266 46338 513502 46574
rect 513586 46338 513822 46574
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -4422 513502 -4186
rect 513586 -4422 513822 -4186
rect 513266 -4742 513502 -4506
rect 513586 -4742 513822 -4506
rect 534986 711322 535222 711558
rect 535306 711322 535542 711558
rect 534986 711002 535222 711238
rect 535306 711002 535542 711238
rect 531266 709402 531502 709638
rect 531586 709402 531822 709638
rect 531266 709082 531502 709318
rect 531586 709082 531822 709318
rect 527546 707482 527782 707718
rect 527866 707482 528102 707718
rect 527546 707162 527782 707398
rect 527866 707162 528102 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 516986 662378 517222 662614
rect 517306 662378 517542 662614
rect 516986 662058 517222 662294
rect 517306 662058 517542 662294
rect 516986 626378 517222 626614
rect 517306 626378 517542 626614
rect 516986 626058 517222 626294
rect 517306 626058 517542 626294
rect 516986 590378 517222 590614
rect 517306 590378 517542 590614
rect 516986 590058 517222 590294
rect 517306 590058 517542 590294
rect 516986 554378 517222 554614
rect 517306 554378 517542 554614
rect 516986 554058 517222 554294
rect 517306 554058 517542 554294
rect 516986 518378 517222 518614
rect 517306 518378 517542 518614
rect 516986 518058 517222 518294
rect 517306 518058 517542 518294
rect 516986 482378 517222 482614
rect 517306 482378 517542 482614
rect 516986 482058 517222 482294
rect 517306 482058 517542 482294
rect 516986 446378 517222 446614
rect 517306 446378 517542 446614
rect 516986 446058 517222 446294
rect 517306 446058 517542 446294
rect 516986 410378 517222 410614
rect 517306 410378 517542 410614
rect 516986 410058 517222 410294
rect 517306 410058 517542 410294
rect 516986 374378 517222 374614
rect 517306 374378 517542 374614
rect 516986 374058 517222 374294
rect 517306 374058 517542 374294
rect 516986 338378 517222 338614
rect 517306 338378 517542 338614
rect 516986 338058 517222 338294
rect 517306 338058 517542 338294
rect 516986 302378 517222 302614
rect 517306 302378 517542 302614
rect 516986 302058 517222 302294
rect 517306 302058 517542 302294
rect 516986 266378 517222 266614
rect 517306 266378 517542 266614
rect 516986 266058 517222 266294
rect 517306 266058 517542 266294
rect 516986 230378 517222 230614
rect 517306 230378 517542 230614
rect 516986 230058 517222 230294
rect 517306 230058 517542 230294
rect 516986 194378 517222 194614
rect 517306 194378 517542 194614
rect 516986 194058 517222 194294
rect 517306 194058 517542 194294
rect 516986 158378 517222 158614
rect 517306 158378 517542 158614
rect 516986 158058 517222 158294
rect 517306 158058 517542 158294
rect 516986 122378 517222 122614
rect 517306 122378 517542 122614
rect 516986 122058 517222 122294
rect 517306 122058 517542 122294
rect 516986 86378 517222 86614
rect 517306 86378 517542 86614
rect 516986 86058 517222 86294
rect 517306 86058 517542 86294
rect 516986 50378 517222 50614
rect 517306 50378 517542 50614
rect 516986 50058 517222 50294
rect 517306 50058 517542 50294
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 498986 -7302 499222 -7066
rect 499306 -7302 499542 -7066
rect 498986 -7622 499222 -7386
rect 499306 -7622 499542 -7386
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -1542 524062 -1306
rect 524146 -1542 524382 -1306
rect 523826 -1862 524062 -1626
rect 524146 -1862 524382 -1626
rect 527546 672938 527782 673174
rect 527866 672938 528102 673174
rect 527546 672618 527782 672854
rect 527866 672618 528102 672854
rect 527546 636938 527782 637174
rect 527866 636938 528102 637174
rect 527546 636618 527782 636854
rect 527866 636618 528102 636854
rect 527546 600938 527782 601174
rect 527866 600938 528102 601174
rect 527546 600618 527782 600854
rect 527866 600618 528102 600854
rect 527546 564938 527782 565174
rect 527866 564938 528102 565174
rect 527546 564618 527782 564854
rect 527866 564618 528102 564854
rect 527546 528938 527782 529174
rect 527866 528938 528102 529174
rect 527546 528618 527782 528854
rect 527866 528618 528102 528854
rect 527546 492938 527782 493174
rect 527866 492938 528102 493174
rect 527546 492618 527782 492854
rect 527866 492618 528102 492854
rect 527546 456938 527782 457174
rect 527866 456938 528102 457174
rect 527546 456618 527782 456854
rect 527866 456618 528102 456854
rect 527546 420938 527782 421174
rect 527866 420938 528102 421174
rect 527546 420618 527782 420854
rect 527866 420618 528102 420854
rect 527546 384938 527782 385174
rect 527866 384938 528102 385174
rect 527546 384618 527782 384854
rect 527866 384618 528102 384854
rect 527546 348938 527782 349174
rect 527866 348938 528102 349174
rect 527546 348618 527782 348854
rect 527866 348618 528102 348854
rect 527546 312938 527782 313174
rect 527866 312938 528102 313174
rect 527546 312618 527782 312854
rect 527866 312618 528102 312854
rect 527546 276938 527782 277174
rect 527866 276938 528102 277174
rect 527546 276618 527782 276854
rect 527866 276618 528102 276854
rect 527546 240938 527782 241174
rect 527866 240938 528102 241174
rect 527546 240618 527782 240854
rect 527866 240618 528102 240854
rect 527546 204938 527782 205174
rect 527866 204938 528102 205174
rect 527546 204618 527782 204854
rect 527866 204618 528102 204854
rect 527546 168938 527782 169174
rect 527866 168938 528102 169174
rect 527546 168618 527782 168854
rect 527866 168618 528102 168854
rect 527546 132938 527782 133174
rect 527866 132938 528102 133174
rect 527546 132618 527782 132854
rect 527866 132618 528102 132854
rect 527546 96938 527782 97174
rect 527866 96938 528102 97174
rect 527546 96618 527782 96854
rect 527866 96618 528102 96854
rect 527546 60938 527782 61174
rect 527866 60938 528102 61174
rect 527546 60618 527782 60854
rect 527866 60618 528102 60854
rect 527546 24938 527782 25174
rect 527866 24938 528102 25174
rect 527546 24618 527782 24854
rect 527866 24618 528102 24854
rect 527546 -3462 527782 -3226
rect 527866 -3462 528102 -3226
rect 527546 -3782 527782 -3546
rect 527866 -3782 528102 -3546
rect 531266 676658 531502 676894
rect 531586 676658 531822 676894
rect 531266 676338 531502 676574
rect 531586 676338 531822 676574
rect 531266 640658 531502 640894
rect 531586 640658 531822 640894
rect 531266 640338 531502 640574
rect 531586 640338 531822 640574
rect 531266 604658 531502 604894
rect 531586 604658 531822 604894
rect 531266 604338 531502 604574
rect 531586 604338 531822 604574
rect 531266 568658 531502 568894
rect 531586 568658 531822 568894
rect 531266 568338 531502 568574
rect 531586 568338 531822 568574
rect 531266 532658 531502 532894
rect 531586 532658 531822 532894
rect 531266 532338 531502 532574
rect 531586 532338 531822 532574
rect 531266 496658 531502 496894
rect 531586 496658 531822 496894
rect 531266 496338 531502 496574
rect 531586 496338 531822 496574
rect 531266 460658 531502 460894
rect 531586 460658 531822 460894
rect 531266 460338 531502 460574
rect 531586 460338 531822 460574
rect 531266 424658 531502 424894
rect 531586 424658 531822 424894
rect 531266 424338 531502 424574
rect 531586 424338 531822 424574
rect 531266 388658 531502 388894
rect 531586 388658 531822 388894
rect 531266 388338 531502 388574
rect 531586 388338 531822 388574
rect 531266 352658 531502 352894
rect 531586 352658 531822 352894
rect 531266 352338 531502 352574
rect 531586 352338 531822 352574
rect 531266 316658 531502 316894
rect 531586 316658 531822 316894
rect 531266 316338 531502 316574
rect 531586 316338 531822 316574
rect 531266 280658 531502 280894
rect 531586 280658 531822 280894
rect 531266 280338 531502 280574
rect 531586 280338 531822 280574
rect 531266 244658 531502 244894
rect 531586 244658 531822 244894
rect 531266 244338 531502 244574
rect 531586 244338 531822 244574
rect 531266 208658 531502 208894
rect 531586 208658 531822 208894
rect 531266 208338 531502 208574
rect 531586 208338 531822 208574
rect 531266 172658 531502 172894
rect 531586 172658 531822 172894
rect 531266 172338 531502 172574
rect 531586 172338 531822 172574
rect 531266 136658 531502 136894
rect 531586 136658 531822 136894
rect 531266 136338 531502 136574
rect 531586 136338 531822 136574
rect 531266 100658 531502 100894
rect 531586 100658 531822 100894
rect 531266 100338 531502 100574
rect 531586 100338 531822 100574
rect 531266 64658 531502 64894
rect 531586 64658 531822 64894
rect 531266 64338 531502 64574
rect 531586 64338 531822 64574
rect 531266 28658 531502 28894
rect 531586 28658 531822 28894
rect 531266 28338 531502 28574
rect 531586 28338 531822 28574
rect 531266 -5382 531502 -5146
rect 531586 -5382 531822 -5146
rect 531266 -5702 531502 -5466
rect 531586 -5702 531822 -5466
rect 552986 710362 553222 710598
rect 553306 710362 553542 710598
rect 552986 710042 553222 710278
rect 553306 710042 553542 710278
rect 549266 708442 549502 708678
rect 549586 708442 549822 708678
rect 549266 708122 549502 708358
rect 549586 708122 549822 708358
rect 545546 706522 545782 706758
rect 545866 706522 546102 706758
rect 545546 706202 545782 706438
rect 545866 706202 546102 706438
rect 534986 680378 535222 680614
rect 535306 680378 535542 680614
rect 534986 680058 535222 680294
rect 535306 680058 535542 680294
rect 534986 644378 535222 644614
rect 535306 644378 535542 644614
rect 534986 644058 535222 644294
rect 535306 644058 535542 644294
rect 534986 608378 535222 608614
rect 535306 608378 535542 608614
rect 534986 608058 535222 608294
rect 535306 608058 535542 608294
rect 534986 572378 535222 572614
rect 535306 572378 535542 572614
rect 534986 572058 535222 572294
rect 535306 572058 535542 572294
rect 534986 536378 535222 536614
rect 535306 536378 535542 536614
rect 534986 536058 535222 536294
rect 535306 536058 535542 536294
rect 534986 500378 535222 500614
rect 535306 500378 535542 500614
rect 534986 500058 535222 500294
rect 535306 500058 535542 500294
rect 534986 464378 535222 464614
rect 535306 464378 535542 464614
rect 534986 464058 535222 464294
rect 535306 464058 535542 464294
rect 534986 428378 535222 428614
rect 535306 428378 535542 428614
rect 534986 428058 535222 428294
rect 535306 428058 535542 428294
rect 534986 392378 535222 392614
rect 535306 392378 535542 392614
rect 534986 392058 535222 392294
rect 535306 392058 535542 392294
rect 534986 356378 535222 356614
rect 535306 356378 535542 356614
rect 534986 356058 535222 356294
rect 535306 356058 535542 356294
rect 534986 320378 535222 320614
rect 535306 320378 535542 320614
rect 534986 320058 535222 320294
rect 535306 320058 535542 320294
rect 534986 284378 535222 284614
rect 535306 284378 535542 284614
rect 534986 284058 535222 284294
rect 535306 284058 535542 284294
rect 534986 248378 535222 248614
rect 535306 248378 535542 248614
rect 534986 248058 535222 248294
rect 535306 248058 535542 248294
rect 534986 212378 535222 212614
rect 535306 212378 535542 212614
rect 534986 212058 535222 212294
rect 535306 212058 535542 212294
rect 534986 176378 535222 176614
rect 535306 176378 535542 176614
rect 534986 176058 535222 176294
rect 535306 176058 535542 176294
rect 534986 140378 535222 140614
rect 535306 140378 535542 140614
rect 534986 140058 535222 140294
rect 535306 140058 535542 140294
rect 534986 104378 535222 104614
rect 535306 104378 535542 104614
rect 534986 104058 535222 104294
rect 535306 104058 535542 104294
rect 534986 68378 535222 68614
rect 535306 68378 535542 68614
rect 534986 68058 535222 68294
rect 535306 68058 535542 68294
rect 534986 32378 535222 32614
rect 535306 32378 535542 32614
rect 534986 32058 535222 32294
rect 535306 32058 535542 32294
rect 516986 -6342 517222 -6106
rect 517306 -6342 517542 -6106
rect 516986 -6662 517222 -6426
rect 517306 -6662 517542 -6426
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 545546 546938 545782 547174
rect 545866 546938 546102 547174
rect 545546 546618 545782 546854
rect 545866 546618 546102 546854
rect 545546 510938 545782 511174
rect 545866 510938 546102 511174
rect 545546 510618 545782 510854
rect 545866 510618 546102 510854
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 545546 402938 545782 403174
rect 545866 402938 546102 403174
rect 545546 402618 545782 402854
rect 545866 402618 546102 402854
rect 545546 366938 545782 367174
rect 545866 366938 546102 367174
rect 545546 366618 545782 366854
rect 545866 366618 546102 366854
rect 545546 330938 545782 331174
rect 545866 330938 546102 331174
rect 545546 330618 545782 330854
rect 545866 330618 546102 330854
rect 545546 294938 545782 295174
rect 545866 294938 546102 295174
rect 545546 294618 545782 294854
rect 545866 294618 546102 294854
rect 545546 258938 545782 259174
rect 545866 258938 546102 259174
rect 545546 258618 545782 258854
rect 545866 258618 546102 258854
rect 545546 222938 545782 223174
rect 545866 222938 546102 223174
rect 545546 222618 545782 222854
rect 545866 222618 546102 222854
rect 545546 186938 545782 187174
rect 545866 186938 546102 187174
rect 545546 186618 545782 186854
rect 545866 186618 546102 186854
rect 545546 150938 545782 151174
rect 545866 150938 546102 151174
rect 545546 150618 545782 150854
rect 545866 150618 546102 150854
rect 545546 114938 545782 115174
rect 545866 114938 546102 115174
rect 545546 114618 545782 114854
rect 545866 114618 546102 114854
rect 545546 78938 545782 79174
rect 545866 78938 546102 79174
rect 545546 78618 545782 78854
rect 545866 78618 546102 78854
rect 545546 42938 545782 43174
rect 545866 42938 546102 43174
rect 545546 42618 545782 42854
rect 545866 42618 546102 42854
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -2502 545782 -2266
rect 545866 -2502 546102 -2266
rect 545546 -2822 545782 -2586
rect 545866 -2822 546102 -2586
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 549266 658658 549502 658894
rect 549586 658658 549822 658894
rect 549266 658338 549502 658574
rect 549586 658338 549822 658574
rect 549266 622658 549502 622894
rect 549586 622658 549822 622894
rect 549266 622338 549502 622574
rect 549586 622338 549822 622574
rect 549266 586658 549502 586894
rect 549586 586658 549822 586894
rect 549266 586338 549502 586574
rect 549586 586338 549822 586574
rect 549266 550658 549502 550894
rect 549586 550658 549822 550894
rect 549266 550338 549502 550574
rect 549586 550338 549822 550574
rect 549266 514658 549502 514894
rect 549586 514658 549822 514894
rect 549266 514338 549502 514574
rect 549586 514338 549822 514574
rect 549266 478658 549502 478894
rect 549586 478658 549822 478894
rect 549266 478338 549502 478574
rect 549586 478338 549822 478574
rect 549266 442658 549502 442894
rect 549586 442658 549822 442894
rect 549266 442338 549502 442574
rect 549586 442338 549822 442574
rect 549266 406658 549502 406894
rect 549586 406658 549822 406894
rect 549266 406338 549502 406574
rect 549586 406338 549822 406574
rect 549266 370658 549502 370894
rect 549586 370658 549822 370894
rect 549266 370338 549502 370574
rect 549586 370338 549822 370574
rect 549266 334658 549502 334894
rect 549586 334658 549822 334894
rect 549266 334338 549502 334574
rect 549586 334338 549822 334574
rect 549266 298658 549502 298894
rect 549586 298658 549822 298894
rect 549266 298338 549502 298574
rect 549586 298338 549822 298574
rect 549266 262658 549502 262894
rect 549586 262658 549822 262894
rect 549266 262338 549502 262574
rect 549586 262338 549822 262574
rect 549266 226658 549502 226894
rect 549586 226658 549822 226894
rect 549266 226338 549502 226574
rect 549586 226338 549822 226574
rect 549266 190658 549502 190894
rect 549586 190658 549822 190894
rect 549266 190338 549502 190574
rect 549586 190338 549822 190574
rect 549266 154658 549502 154894
rect 549586 154658 549822 154894
rect 549266 154338 549502 154574
rect 549586 154338 549822 154574
rect 549266 118658 549502 118894
rect 549586 118658 549822 118894
rect 549266 118338 549502 118574
rect 549586 118338 549822 118574
rect 549266 82658 549502 82894
rect 549586 82658 549822 82894
rect 549266 82338 549502 82574
rect 549586 82338 549822 82574
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -4422 549502 -4186
rect 549586 -4422 549822 -4186
rect 549266 -4742 549502 -4506
rect 549586 -4742 549822 -4506
rect 570986 711322 571222 711558
rect 571306 711322 571542 711558
rect 570986 711002 571222 711238
rect 571306 711002 571542 711238
rect 567266 709402 567502 709638
rect 567586 709402 567822 709638
rect 567266 709082 567502 709318
rect 567586 709082 567822 709318
rect 563546 707482 563782 707718
rect 563866 707482 564102 707718
rect 563546 707162 563782 707398
rect 563866 707162 564102 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 552986 626378 553222 626614
rect 553306 626378 553542 626614
rect 552986 626058 553222 626294
rect 553306 626058 553542 626294
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 552986 554378 553222 554614
rect 553306 554378 553542 554614
rect 552986 554058 553222 554294
rect 553306 554058 553542 554294
rect 552986 518378 553222 518614
rect 553306 518378 553542 518614
rect 552986 518058 553222 518294
rect 553306 518058 553542 518294
rect 552986 482378 553222 482614
rect 553306 482378 553542 482614
rect 552986 482058 553222 482294
rect 553306 482058 553542 482294
rect 552986 446378 553222 446614
rect 553306 446378 553542 446614
rect 552986 446058 553222 446294
rect 553306 446058 553542 446294
rect 552986 410378 553222 410614
rect 553306 410378 553542 410614
rect 552986 410058 553222 410294
rect 553306 410058 553542 410294
rect 552986 374378 553222 374614
rect 553306 374378 553542 374614
rect 552986 374058 553222 374294
rect 553306 374058 553542 374294
rect 552986 338378 553222 338614
rect 553306 338378 553542 338614
rect 552986 338058 553222 338294
rect 553306 338058 553542 338294
rect 552986 302378 553222 302614
rect 553306 302378 553542 302614
rect 552986 302058 553222 302294
rect 553306 302058 553542 302294
rect 552986 266378 553222 266614
rect 553306 266378 553542 266614
rect 552986 266058 553222 266294
rect 553306 266058 553542 266294
rect 552986 230378 553222 230614
rect 553306 230378 553542 230614
rect 552986 230058 553222 230294
rect 553306 230058 553542 230294
rect 552986 194378 553222 194614
rect 553306 194378 553542 194614
rect 552986 194058 553222 194294
rect 553306 194058 553542 194294
rect 552986 158378 553222 158614
rect 553306 158378 553542 158614
rect 552986 158058 553222 158294
rect 553306 158058 553542 158294
rect 552986 122378 553222 122614
rect 553306 122378 553542 122614
rect 552986 122058 553222 122294
rect 553306 122058 553542 122294
rect 552986 86378 553222 86614
rect 553306 86378 553542 86614
rect 552986 86058 553222 86294
rect 553306 86058 553542 86294
rect 552986 50378 553222 50614
rect 553306 50378 553542 50614
rect 552986 50058 553222 50294
rect 553306 50058 553542 50294
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 534986 -7302 535222 -7066
rect 535306 -7302 535542 -7066
rect 534986 -7622 535222 -7386
rect 535306 -7622 535542 -7386
rect 559826 705562 560062 705798
rect 560146 705562 560382 705798
rect 559826 705242 560062 705478
rect 560146 705242 560382 705478
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -1542 560062 -1306
rect 560146 -1542 560382 -1306
rect 559826 -1862 560062 -1626
rect 560146 -1862 560382 -1626
rect 563546 672938 563782 673174
rect 563866 672938 564102 673174
rect 563546 672618 563782 672854
rect 563866 672618 564102 672854
rect 563546 636938 563782 637174
rect 563866 636938 564102 637174
rect 563546 636618 563782 636854
rect 563866 636618 564102 636854
rect 563546 600938 563782 601174
rect 563866 600938 564102 601174
rect 563546 600618 563782 600854
rect 563866 600618 564102 600854
rect 563546 564938 563782 565174
rect 563866 564938 564102 565174
rect 563546 564618 563782 564854
rect 563866 564618 564102 564854
rect 563546 528938 563782 529174
rect 563866 528938 564102 529174
rect 563546 528618 563782 528854
rect 563866 528618 564102 528854
rect 563546 492938 563782 493174
rect 563866 492938 564102 493174
rect 563546 492618 563782 492854
rect 563866 492618 564102 492854
rect 563546 456938 563782 457174
rect 563866 456938 564102 457174
rect 563546 456618 563782 456854
rect 563866 456618 564102 456854
rect 563546 420938 563782 421174
rect 563866 420938 564102 421174
rect 563546 420618 563782 420854
rect 563866 420618 564102 420854
rect 563546 384938 563782 385174
rect 563866 384938 564102 385174
rect 563546 384618 563782 384854
rect 563866 384618 564102 384854
rect 563546 348938 563782 349174
rect 563866 348938 564102 349174
rect 563546 348618 563782 348854
rect 563866 348618 564102 348854
rect 563546 312938 563782 313174
rect 563866 312938 564102 313174
rect 563546 312618 563782 312854
rect 563866 312618 564102 312854
rect 563546 276938 563782 277174
rect 563866 276938 564102 277174
rect 563546 276618 563782 276854
rect 563866 276618 564102 276854
rect 563546 240938 563782 241174
rect 563866 240938 564102 241174
rect 563546 240618 563782 240854
rect 563866 240618 564102 240854
rect 563546 204938 563782 205174
rect 563866 204938 564102 205174
rect 563546 204618 563782 204854
rect 563866 204618 564102 204854
rect 563546 168938 563782 169174
rect 563866 168938 564102 169174
rect 563546 168618 563782 168854
rect 563866 168618 564102 168854
rect 563546 132938 563782 133174
rect 563866 132938 564102 133174
rect 563546 132618 563782 132854
rect 563866 132618 564102 132854
rect 563546 96938 563782 97174
rect 563866 96938 564102 97174
rect 563546 96618 563782 96854
rect 563866 96618 564102 96854
rect 563546 60938 563782 61174
rect 563866 60938 564102 61174
rect 563546 60618 563782 60854
rect 563866 60618 564102 60854
rect 563546 24938 563782 25174
rect 563866 24938 564102 25174
rect 563546 24618 563782 24854
rect 563866 24618 564102 24854
rect 563546 -3462 563782 -3226
rect 563866 -3462 564102 -3226
rect 563546 -3782 563782 -3546
rect 563866 -3782 564102 -3546
rect 567266 676658 567502 676894
rect 567586 676658 567822 676894
rect 567266 676338 567502 676574
rect 567586 676338 567822 676574
rect 567266 640658 567502 640894
rect 567586 640658 567822 640894
rect 567266 640338 567502 640574
rect 567586 640338 567822 640574
rect 567266 604658 567502 604894
rect 567586 604658 567822 604894
rect 567266 604338 567502 604574
rect 567586 604338 567822 604574
rect 567266 568658 567502 568894
rect 567586 568658 567822 568894
rect 567266 568338 567502 568574
rect 567586 568338 567822 568574
rect 567266 532658 567502 532894
rect 567586 532658 567822 532894
rect 567266 532338 567502 532574
rect 567586 532338 567822 532574
rect 567266 496658 567502 496894
rect 567586 496658 567822 496894
rect 567266 496338 567502 496574
rect 567586 496338 567822 496574
rect 567266 460658 567502 460894
rect 567586 460658 567822 460894
rect 567266 460338 567502 460574
rect 567586 460338 567822 460574
rect 567266 424658 567502 424894
rect 567586 424658 567822 424894
rect 567266 424338 567502 424574
rect 567586 424338 567822 424574
rect 567266 388658 567502 388894
rect 567586 388658 567822 388894
rect 567266 388338 567502 388574
rect 567586 388338 567822 388574
rect 567266 352658 567502 352894
rect 567586 352658 567822 352894
rect 567266 352338 567502 352574
rect 567586 352338 567822 352574
rect 567266 316658 567502 316894
rect 567586 316658 567822 316894
rect 567266 316338 567502 316574
rect 567586 316338 567822 316574
rect 567266 280658 567502 280894
rect 567586 280658 567822 280894
rect 567266 280338 567502 280574
rect 567586 280338 567822 280574
rect 567266 244658 567502 244894
rect 567586 244658 567822 244894
rect 567266 244338 567502 244574
rect 567586 244338 567822 244574
rect 567266 208658 567502 208894
rect 567586 208658 567822 208894
rect 567266 208338 567502 208574
rect 567586 208338 567822 208574
rect 567266 172658 567502 172894
rect 567586 172658 567822 172894
rect 567266 172338 567502 172574
rect 567586 172338 567822 172574
rect 567266 136658 567502 136894
rect 567586 136658 567822 136894
rect 567266 136338 567502 136574
rect 567586 136338 567822 136574
rect 567266 100658 567502 100894
rect 567586 100658 567822 100894
rect 567266 100338 567502 100574
rect 567586 100338 567822 100574
rect 567266 64658 567502 64894
rect 567586 64658 567822 64894
rect 567266 64338 567502 64574
rect 567586 64338 567822 64574
rect 567266 28658 567502 28894
rect 567586 28658 567822 28894
rect 567266 28338 567502 28574
rect 567586 28338 567822 28574
rect 567266 -5382 567502 -5146
rect 567586 -5382 567822 -5146
rect 567266 -5702 567502 -5466
rect 567586 -5702 567822 -5466
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 581546 706522 581782 706758
rect 581866 706522 582102 706758
rect 581546 706202 581782 706438
rect 581866 706202 582102 706438
rect 570986 680378 571222 680614
rect 571306 680378 571542 680614
rect 570986 680058 571222 680294
rect 571306 680058 571542 680294
rect 570986 644378 571222 644614
rect 571306 644378 571542 644614
rect 570986 644058 571222 644294
rect 571306 644058 571542 644294
rect 570986 608378 571222 608614
rect 571306 608378 571542 608614
rect 570986 608058 571222 608294
rect 571306 608058 571542 608294
rect 570986 572378 571222 572614
rect 571306 572378 571542 572614
rect 570986 572058 571222 572294
rect 571306 572058 571542 572294
rect 570986 536378 571222 536614
rect 571306 536378 571542 536614
rect 570986 536058 571222 536294
rect 571306 536058 571542 536294
rect 570986 500378 571222 500614
rect 571306 500378 571542 500614
rect 570986 500058 571222 500294
rect 571306 500058 571542 500294
rect 570986 464378 571222 464614
rect 571306 464378 571542 464614
rect 570986 464058 571222 464294
rect 571306 464058 571542 464294
rect 570986 428378 571222 428614
rect 571306 428378 571542 428614
rect 570986 428058 571222 428294
rect 571306 428058 571542 428294
rect 570986 392378 571222 392614
rect 571306 392378 571542 392614
rect 570986 392058 571222 392294
rect 571306 392058 571542 392294
rect 570986 356378 571222 356614
rect 571306 356378 571542 356614
rect 570986 356058 571222 356294
rect 571306 356058 571542 356294
rect 570986 320378 571222 320614
rect 571306 320378 571542 320614
rect 570986 320058 571222 320294
rect 571306 320058 571542 320294
rect 570986 284378 571222 284614
rect 571306 284378 571542 284614
rect 570986 284058 571222 284294
rect 571306 284058 571542 284294
rect 570986 248378 571222 248614
rect 571306 248378 571542 248614
rect 570986 248058 571222 248294
rect 571306 248058 571542 248294
rect 570986 212378 571222 212614
rect 571306 212378 571542 212614
rect 570986 212058 571222 212294
rect 571306 212058 571542 212294
rect 570986 176378 571222 176614
rect 571306 176378 571542 176614
rect 570986 176058 571222 176294
rect 571306 176058 571542 176294
rect 570986 140378 571222 140614
rect 571306 140378 571542 140614
rect 570986 140058 571222 140294
rect 571306 140058 571542 140294
rect 570986 104378 571222 104614
rect 571306 104378 571542 104614
rect 570986 104058 571222 104294
rect 571306 104058 571542 104294
rect 570986 68378 571222 68614
rect 571306 68378 571542 68614
rect 570986 68058 571222 68294
rect 571306 68058 571542 68294
rect 570986 32378 571222 32614
rect 571306 32378 571542 32614
rect 570986 32058 571222 32294
rect 571306 32058 571542 32294
rect 552986 -6342 553222 -6106
rect 553306 -6342 553542 -6106
rect 552986 -6662 553222 -6426
rect 553306 -6662 553542 -6426
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 690938 587498 691174
rect 587582 690938 587818 691174
rect 587262 690618 587498 690854
rect 587582 690618 587818 690854
rect 587262 654938 587498 655174
rect 587582 654938 587818 655174
rect 587262 654618 587498 654854
rect 587582 654618 587818 654854
rect 587262 618938 587498 619174
rect 587582 618938 587818 619174
rect 587262 618618 587498 618854
rect 587582 618618 587818 618854
rect 587262 582938 587498 583174
rect 587582 582938 587818 583174
rect 587262 582618 587498 582854
rect 587582 582618 587818 582854
rect 587262 546938 587498 547174
rect 587582 546938 587818 547174
rect 587262 546618 587498 546854
rect 587582 546618 587818 546854
rect 587262 510938 587498 511174
rect 587582 510938 587818 511174
rect 587262 510618 587498 510854
rect 587582 510618 587818 510854
rect 587262 474938 587498 475174
rect 587582 474938 587818 475174
rect 587262 474618 587498 474854
rect 587582 474618 587818 474854
rect 587262 438938 587498 439174
rect 587582 438938 587818 439174
rect 587262 438618 587498 438854
rect 587582 438618 587818 438854
rect 587262 402938 587498 403174
rect 587582 402938 587818 403174
rect 587262 402618 587498 402854
rect 587582 402618 587818 402854
rect 587262 366938 587498 367174
rect 587582 366938 587818 367174
rect 587262 366618 587498 366854
rect 587582 366618 587818 366854
rect 587262 330938 587498 331174
rect 587582 330938 587818 331174
rect 587262 330618 587498 330854
rect 587582 330618 587818 330854
rect 587262 294938 587498 295174
rect 587582 294938 587818 295174
rect 587262 294618 587498 294854
rect 587582 294618 587818 294854
rect 587262 258938 587498 259174
rect 587582 258938 587818 259174
rect 587262 258618 587498 258854
rect 587582 258618 587818 258854
rect 587262 222938 587498 223174
rect 587582 222938 587818 223174
rect 587262 222618 587498 222854
rect 587582 222618 587818 222854
rect 587262 186938 587498 187174
rect 587582 186938 587818 187174
rect 587262 186618 587498 186854
rect 587582 186618 587818 186854
rect 587262 150938 587498 151174
rect 587582 150938 587818 151174
rect 587262 150618 587498 150854
rect 587582 150618 587818 150854
rect 587262 114938 587498 115174
rect 587582 114938 587818 115174
rect 587262 114618 587498 114854
rect 587582 114618 587818 114854
rect 587262 78938 587498 79174
rect 587582 78938 587818 79174
rect 587262 78618 587498 78854
rect 587582 78618 587818 78854
rect 587262 42938 587498 43174
rect 587582 42938 587818 43174
rect 587262 42618 587498 42854
rect 587582 42618 587818 42854
rect 587262 6938 587498 7174
rect 587582 6938 587818 7174
rect 587262 6618 587498 6854
rect 587582 6618 587818 6854
rect 581546 -2502 581782 -2266
rect 581866 -2502 582102 -2266
rect 581546 -2822 581782 -2586
rect 581866 -2822 582102 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 672938 588458 673174
rect 588542 672938 588778 673174
rect 588222 672618 588458 672854
rect 588542 672618 588778 672854
rect 588222 636938 588458 637174
rect 588542 636938 588778 637174
rect 588222 636618 588458 636854
rect 588542 636618 588778 636854
rect 588222 600938 588458 601174
rect 588542 600938 588778 601174
rect 588222 600618 588458 600854
rect 588542 600618 588778 600854
rect 588222 564938 588458 565174
rect 588542 564938 588778 565174
rect 588222 564618 588458 564854
rect 588542 564618 588778 564854
rect 588222 528938 588458 529174
rect 588542 528938 588778 529174
rect 588222 528618 588458 528854
rect 588542 528618 588778 528854
rect 588222 492938 588458 493174
rect 588542 492938 588778 493174
rect 588222 492618 588458 492854
rect 588542 492618 588778 492854
rect 588222 456938 588458 457174
rect 588542 456938 588778 457174
rect 588222 456618 588458 456854
rect 588542 456618 588778 456854
rect 588222 420938 588458 421174
rect 588542 420938 588778 421174
rect 588222 420618 588458 420854
rect 588542 420618 588778 420854
rect 588222 384938 588458 385174
rect 588542 384938 588778 385174
rect 588222 384618 588458 384854
rect 588542 384618 588778 384854
rect 588222 348938 588458 349174
rect 588542 348938 588778 349174
rect 588222 348618 588458 348854
rect 588542 348618 588778 348854
rect 588222 312938 588458 313174
rect 588542 312938 588778 313174
rect 588222 312618 588458 312854
rect 588542 312618 588778 312854
rect 588222 276938 588458 277174
rect 588542 276938 588778 277174
rect 588222 276618 588458 276854
rect 588542 276618 588778 276854
rect 588222 240938 588458 241174
rect 588542 240938 588778 241174
rect 588222 240618 588458 240854
rect 588542 240618 588778 240854
rect 588222 204938 588458 205174
rect 588542 204938 588778 205174
rect 588222 204618 588458 204854
rect 588542 204618 588778 204854
rect 588222 168938 588458 169174
rect 588542 168938 588778 169174
rect 588222 168618 588458 168854
rect 588542 168618 588778 168854
rect 588222 132938 588458 133174
rect 588542 132938 588778 133174
rect 588222 132618 588458 132854
rect 588542 132618 588778 132854
rect 588222 96938 588458 97174
rect 588542 96938 588778 97174
rect 588222 96618 588458 96854
rect 588542 96618 588778 96854
rect 588222 60938 588458 61174
rect 588542 60938 588778 61174
rect 588222 60618 588458 60854
rect 588542 60618 588778 60854
rect 588222 24938 588458 25174
rect 588542 24938 588778 25174
rect 588222 24618 588458 24854
rect 588542 24618 588778 24854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 694658 589418 694894
rect 589502 694658 589738 694894
rect 589182 694338 589418 694574
rect 589502 694338 589738 694574
rect 589182 658658 589418 658894
rect 589502 658658 589738 658894
rect 589182 658338 589418 658574
rect 589502 658338 589738 658574
rect 589182 622658 589418 622894
rect 589502 622658 589738 622894
rect 589182 622338 589418 622574
rect 589502 622338 589738 622574
rect 589182 586658 589418 586894
rect 589502 586658 589738 586894
rect 589182 586338 589418 586574
rect 589502 586338 589738 586574
rect 589182 550658 589418 550894
rect 589502 550658 589738 550894
rect 589182 550338 589418 550574
rect 589502 550338 589738 550574
rect 589182 514658 589418 514894
rect 589502 514658 589738 514894
rect 589182 514338 589418 514574
rect 589502 514338 589738 514574
rect 589182 478658 589418 478894
rect 589502 478658 589738 478894
rect 589182 478338 589418 478574
rect 589502 478338 589738 478574
rect 589182 442658 589418 442894
rect 589502 442658 589738 442894
rect 589182 442338 589418 442574
rect 589502 442338 589738 442574
rect 589182 406658 589418 406894
rect 589502 406658 589738 406894
rect 589182 406338 589418 406574
rect 589502 406338 589738 406574
rect 589182 370658 589418 370894
rect 589502 370658 589738 370894
rect 589182 370338 589418 370574
rect 589502 370338 589738 370574
rect 589182 334658 589418 334894
rect 589502 334658 589738 334894
rect 589182 334338 589418 334574
rect 589502 334338 589738 334574
rect 589182 298658 589418 298894
rect 589502 298658 589738 298894
rect 589182 298338 589418 298574
rect 589502 298338 589738 298574
rect 589182 262658 589418 262894
rect 589502 262658 589738 262894
rect 589182 262338 589418 262574
rect 589502 262338 589738 262574
rect 589182 226658 589418 226894
rect 589502 226658 589738 226894
rect 589182 226338 589418 226574
rect 589502 226338 589738 226574
rect 589182 190658 589418 190894
rect 589502 190658 589738 190894
rect 589182 190338 589418 190574
rect 589502 190338 589738 190574
rect 589182 154658 589418 154894
rect 589502 154658 589738 154894
rect 589182 154338 589418 154574
rect 589502 154338 589738 154574
rect 589182 118658 589418 118894
rect 589502 118658 589738 118894
rect 589182 118338 589418 118574
rect 589502 118338 589738 118574
rect 589182 82658 589418 82894
rect 589502 82658 589738 82894
rect 589182 82338 589418 82574
rect 589502 82338 589738 82574
rect 589182 46658 589418 46894
rect 589502 46658 589738 46894
rect 589182 46338 589418 46574
rect 589502 46338 589738 46574
rect 589182 10658 589418 10894
rect 589502 10658 589738 10894
rect 589182 10338 589418 10574
rect 589502 10338 589738 10574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 676658 590378 676894
rect 590462 676658 590698 676894
rect 590142 676338 590378 676574
rect 590462 676338 590698 676574
rect 590142 640658 590378 640894
rect 590462 640658 590698 640894
rect 590142 640338 590378 640574
rect 590462 640338 590698 640574
rect 590142 604658 590378 604894
rect 590462 604658 590698 604894
rect 590142 604338 590378 604574
rect 590462 604338 590698 604574
rect 590142 568658 590378 568894
rect 590462 568658 590698 568894
rect 590142 568338 590378 568574
rect 590462 568338 590698 568574
rect 590142 532658 590378 532894
rect 590462 532658 590698 532894
rect 590142 532338 590378 532574
rect 590462 532338 590698 532574
rect 590142 496658 590378 496894
rect 590462 496658 590698 496894
rect 590142 496338 590378 496574
rect 590462 496338 590698 496574
rect 590142 460658 590378 460894
rect 590462 460658 590698 460894
rect 590142 460338 590378 460574
rect 590462 460338 590698 460574
rect 590142 424658 590378 424894
rect 590462 424658 590698 424894
rect 590142 424338 590378 424574
rect 590462 424338 590698 424574
rect 590142 388658 590378 388894
rect 590462 388658 590698 388894
rect 590142 388338 590378 388574
rect 590462 388338 590698 388574
rect 590142 352658 590378 352894
rect 590462 352658 590698 352894
rect 590142 352338 590378 352574
rect 590462 352338 590698 352574
rect 590142 316658 590378 316894
rect 590462 316658 590698 316894
rect 590142 316338 590378 316574
rect 590462 316338 590698 316574
rect 590142 280658 590378 280894
rect 590462 280658 590698 280894
rect 590142 280338 590378 280574
rect 590462 280338 590698 280574
rect 590142 244658 590378 244894
rect 590462 244658 590698 244894
rect 590142 244338 590378 244574
rect 590462 244338 590698 244574
rect 590142 208658 590378 208894
rect 590462 208658 590698 208894
rect 590142 208338 590378 208574
rect 590462 208338 590698 208574
rect 590142 172658 590378 172894
rect 590462 172658 590698 172894
rect 590142 172338 590378 172574
rect 590462 172338 590698 172574
rect 590142 136658 590378 136894
rect 590462 136658 590698 136894
rect 590142 136338 590378 136574
rect 590462 136338 590698 136574
rect 590142 100658 590378 100894
rect 590462 100658 590698 100894
rect 590142 100338 590378 100574
rect 590462 100338 590698 100574
rect 590142 64658 590378 64894
rect 590462 64658 590698 64894
rect 590142 64338 590378 64574
rect 590462 64338 590698 64574
rect 590142 28658 590378 28894
rect 590462 28658 590698 28894
rect 590142 28338 590378 28574
rect 590462 28338 590698 28574
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 698378 591338 698614
rect 591422 698378 591658 698614
rect 591102 698058 591338 698294
rect 591422 698058 591658 698294
rect 591102 662378 591338 662614
rect 591422 662378 591658 662614
rect 591102 662058 591338 662294
rect 591422 662058 591658 662294
rect 591102 626378 591338 626614
rect 591422 626378 591658 626614
rect 591102 626058 591338 626294
rect 591422 626058 591658 626294
rect 591102 590378 591338 590614
rect 591422 590378 591658 590614
rect 591102 590058 591338 590294
rect 591422 590058 591658 590294
rect 591102 554378 591338 554614
rect 591422 554378 591658 554614
rect 591102 554058 591338 554294
rect 591422 554058 591658 554294
rect 591102 518378 591338 518614
rect 591422 518378 591658 518614
rect 591102 518058 591338 518294
rect 591422 518058 591658 518294
rect 591102 482378 591338 482614
rect 591422 482378 591658 482614
rect 591102 482058 591338 482294
rect 591422 482058 591658 482294
rect 591102 446378 591338 446614
rect 591422 446378 591658 446614
rect 591102 446058 591338 446294
rect 591422 446058 591658 446294
rect 591102 410378 591338 410614
rect 591422 410378 591658 410614
rect 591102 410058 591338 410294
rect 591422 410058 591658 410294
rect 591102 374378 591338 374614
rect 591422 374378 591658 374614
rect 591102 374058 591338 374294
rect 591422 374058 591658 374294
rect 591102 338378 591338 338614
rect 591422 338378 591658 338614
rect 591102 338058 591338 338294
rect 591422 338058 591658 338294
rect 591102 302378 591338 302614
rect 591422 302378 591658 302614
rect 591102 302058 591338 302294
rect 591422 302058 591658 302294
rect 591102 266378 591338 266614
rect 591422 266378 591658 266614
rect 591102 266058 591338 266294
rect 591422 266058 591658 266294
rect 591102 230378 591338 230614
rect 591422 230378 591658 230614
rect 591102 230058 591338 230294
rect 591422 230058 591658 230294
rect 591102 194378 591338 194614
rect 591422 194378 591658 194614
rect 591102 194058 591338 194294
rect 591422 194058 591658 194294
rect 591102 158378 591338 158614
rect 591422 158378 591658 158614
rect 591102 158058 591338 158294
rect 591422 158058 591658 158294
rect 591102 122378 591338 122614
rect 591422 122378 591658 122614
rect 591102 122058 591338 122294
rect 591422 122058 591658 122294
rect 591102 86378 591338 86614
rect 591422 86378 591658 86614
rect 591102 86058 591338 86294
rect 591422 86058 591658 86294
rect 591102 50378 591338 50614
rect 591422 50378 591658 50614
rect 591102 50058 591338 50294
rect 591422 50058 591658 50294
rect 591102 14378 591338 14614
rect 591422 14378 591658 14614
rect 591102 14058 591338 14294
rect 591422 14058 591658 14294
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 680378 592298 680614
rect 592382 680378 592618 680614
rect 592062 680058 592298 680294
rect 592382 680058 592618 680294
rect 592062 644378 592298 644614
rect 592382 644378 592618 644614
rect 592062 644058 592298 644294
rect 592382 644058 592618 644294
rect 592062 608378 592298 608614
rect 592382 608378 592618 608614
rect 592062 608058 592298 608294
rect 592382 608058 592618 608294
rect 592062 572378 592298 572614
rect 592382 572378 592618 572614
rect 592062 572058 592298 572294
rect 592382 572058 592618 572294
rect 592062 536378 592298 536614
rect 592382 536378 592618 536614
rect 592062 536058 592298 536294
rect 592382 536058 592618 536294
rect 592062 500378 592298 500614
rect 592382 500378 592618 500614
rect 592062 500058 592298 500294
rect 592382 500058 592618 500294
rect 592062 464378 592298 464614
rect 592382 464378 592618 464614
rect 592062 464058 592298 464294
rect 592382 464058 592618 464294
rect 592062 428378 592298 428614
rect 592382 428378 592618 428614
rect 592062 428058 592298 428294
rect 592382 428058 592618 428294
rect 592062 392378 592298 392614
rect 592382 392378 592618 392614
rect 592062 392058 592298 392294
rect 592382 392058 592618 392294
rect 592062 356378 592298 356614
rect 592382 356378 592618 356614
rect 592062 356058 592298 356294
rect 592382 356058 592618 356294
rect 592062 320378 592298 320614
rect 592382 320378 592618 320614
rect 592062 320058 592298 320294
rect 592382 320058 592618 320294
rect 592062 284378 592298 284614
rect 592382 284378 592618 284614
rect 592062 284058 592298 284294
rect 592382 284058 592618 284294
rect 592062 248378 592298 248614
rect 592382 248378 592618 248614
rect 592062 248058 592298 248294
rect 592382 248058 592618 248294
rect 592062 212378 592298 212614
rect 592382 212378 592618 212614
rect 592062 212058 592298 212294
rect 592382 212058 592618 212294
rect 592062 176378 592298 176614
rect 592382 176378 592618 176614
rect 592062 176058 592298 176294
rect 592382 176058 592618 176294
rect 592062 140378 592298 140614
rect 592382 140378 592618 140614
rect 592062 140058 592298 140294
rect 592382 140058 592618 140294
rect 592062 104378 592298 104614
rect 592382 104378 592618 104614
rect 592062 104058 592298 104294
rect 592382 104058 592618 104294
rect 592062 68378 592298 68614
rect 592382 68378 592618 68614
rect 592062 68058 592298 68294
rect 592382 68058 592618 68294
rect 592062 32378 592298 32614
rect 592382 32378 592618 32614
rect 592062 32058 592298 32294
rect 592382 32058 592618 32294
rect 570986 -7302 571222 -7066
rect 571306 -7302 571542 -7066
rect 570986 -7622 571222 -7386
rect 571306 -7622 571542 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 592650 698294
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 590730 694894
rect -6806 694574 590730 694658
rect -6806 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 590730 694574
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 588810 691174
rect -4886 690854 588810 690938
rect -4886 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 588810 690854
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect -8726 680294 592650 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect -6806 676574 590730 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect -4886 672854 588810 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 592650 662294
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 590730 658894
rect -6806 658574 590730 658658
rect -6806 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 590730 658574
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 588810 655174
rect -4886 654854 588810 654938
rect -4886 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 588810 654854
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect -8726 644294 592650 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect -6806 640574 590730 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect -4886 636854 588810 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 592650 626294
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 590730 622894
rect -6806 622574 590730 622658
rect -6806 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 590730 622574
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 588810 619174
rect -4886 618854 588810 618938
rect -4886 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 588810 618854
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect -8726 608294 592650 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect -6806 604574 590730 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect -4886 600854 588810 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 592650 590294
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 590730 586894
rect -6806 586574 590730 586658
rect -6806 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 590730 586574
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 588810 583174
rect -4886 582854 588810 582938
rect -4886 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 588810 582854
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect -8726 572294 592650 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect -6806 568574 590730 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect -4886 564854 588810 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect -4886 564586 588810 564618
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 592650 554294
rect -8726 554026 592650 554058
rect -6806 550894 590730 550926
rect -6806 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 590730 550894
rect -6806 550574 590730 550658
rect -6806 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 590730 550574
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 588810 547174
rect -4886 546854 588810 546938
rect -4886 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 588810 546854
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect -8726 536294 592650 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect -6806 532574 590730 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect -4886 528854 588810 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 592650 518294
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 590730 514894
rect -6806 514574 590730 514658
rect -6806 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 590730 514574
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 588810 511174
rect -4886 510854 588810 510938
rect -4886 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 588810 510854
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect -8726 500294 592650 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect -6806 496574 590730 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect -4886 492854 588810 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 592650 482294
rect -8726 482026 592650 482058
rect -6806 478894 590730 478926
rect -6806 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 590730 478894
rect -6806 478574 590730 478658
rect -6806 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 590730 478574
rect -6806 478306 590730 478338
rect -4886 475174 588810 475206
rect -4886 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 588810 475174
rect -4886 474854 588810 474938
rect -4886 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 588810 474854
rect -4886 474586 588810 474618
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 61008 471454
rect 61244 471218 195376 471454
rect 195612 471218 221008 471454
rect 221244 471218 355376 471454
rect 355612 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 61008 471134
rect 61244 470898 195376 471134
rect 195612 470898 221008 471134
rect 221244 470898 355376 471134
rect 355612 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect -8726 464294 592650 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect -6806 460574 590730 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect -4886 456854 588810 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 60328 453454
rect 60564 453218 196056 453454
rect 196292 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 220328 453454
rect 220564 453218 356056 453454
rect 356292 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 60328 453134
rect 60564 452898 196056 453134
rect 196292 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 220328 453134
rect 220564 452898 356056 453134
rect 356292 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 592650 446294
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 590730 442894
rect -6806 442574 590730 442658
rect -6806 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 590730 442574
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 588810 439174
rect -4886 438854 588810 438938
rect -4886 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 588810 438854
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 61008 435454
rect 61244 435218 195376 435454
rect 195612 435218 221008 435454
rect 221244 435218 355376 435454
rect 355612 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 61008 435134
rect 61244 434898 195376 435134
rect 195612 434898 221008 435134
rect 221244 434898 355376 435134
rect 355612 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 390986 428614
rect 391222 428378 391306 428614
rect 391542 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect -8726 428294 592650 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 390986 428294
rect 391222 428058 391306 428294
rect 391542 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 387266 424894
rect 387502 424658 387586 424894
rect 387822 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect -6806 424574 590730 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 387266 424574
rect 387502 424338 387586 424574
rect 387822 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 383546 421174
rect 383782 420938 383866 421174
rect 384102 420938 419546 421174
rect 419782 420938 419866 421174
rect 420102 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect -4886 420854 588810 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 383546 420854
rect 383782 420618 383866 420854
rect 384102 420618 419546 420854
rect 419782 420618 419866 420854
rect 420102 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 60328 417454
rect 60564 417218 196056 417454
rect 196292 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 220328 417454
rect 220564 417218 356056 417454
rect 356292 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 60328 417134
rect 60564 416898 196056 417134
rect 196292 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 220328 417134
rect 220564 416898 356056 417134
rect 356292 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 592650 410294
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 590730 406894
rect -6806 406574 590730 406658
rect -6806 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 590730 406574
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 588810 403174
rect -4886 402854 588810 402938
rect -4886 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 588810 402854
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 66986 392614
rect 67222 392378 67306 392614
rect 67542 392378 102986 392614
rect 103222 392378 103306 392614
rect 103542 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 210986 392614
rect 211222 392378 211306 392614
rect 211542 392378 246986 392614
rect 247222 392378 247306 392614
rect 247542 392378 282986 392614
rect 283222 392378 283306 392614
rect 283542 392378 318986 392614
rect 319222 392378 319306 392614
rect 319542 392378 354986 392614
rect 355222 392378 355306 392614
rect 355542 392378 390986 392614
rect 391222 392378 391306 392614
rect 391542 392378 426986 392614
rect 427222 392378 427306 392614
rect 427542 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect -8726 392294 592650 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 66986 392294
rect 67222 392058 67306 392294
rect 67542 392058 102986 392294
rect 103222 392058 103306 392294
rect 103542 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 210986 392294
rect 211222 392058 211306 392294
rect 211542 392058 246986 392294
rect 247222 392058 247306 392294
rect 247542 392058 282986 392294
rect 283222 392058 283306 392294
rect 283542 392058 318986 392294
rect 319222 392058 319306 392294
rect 319542 392058 354986 392294
rect 355222 392058 355306 392294
rect 355542 392058 390986 392294
rect 391222 392058 391306 392294
rect 391542 392058 426986 392294
rect 427222 392058 427306 392294
rect 427542 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect -8726 392026 592650 392058
rect -6806 388894 590730 388926
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 99266 388894
rect 99502 388658 99586 388894
rect 99822 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 171266 388894
rect 171502 388658 171586 388894
rect 171822 388658 207266 388894
rect 207502 388658 207586 388894
rect 207822 388658 243266 388894
rect 243502 388658 243586 388894
rect 243822 388658 279266 388894
rect 279502 388658 279586 388894
rect 279822 388658 315266 388894
rect 315502 388658 315586 388894
rect 315822 388658 351266 388894
rect 351502 388658 351586 388894
rect 351822 388658 387266 388894
rect 387502 388658 387586 388894
rect 387822 388658 423266 388894
rect 423502 388658 423586 388894
rect 423822 388658 459266 388894
rect 459502 388658 459586 388894
rect 459822 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect -6806 388574 590730 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 99266 388574
rect 99502 388338 99586 388574
rect 99822 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 171266 388574
rect 171502 388338 171586 388574
rect 171822 388338 207266 388574
rect 207502 388338 207586 388574
rect 207822 388338 243266 388574
rect 243502 388338 243586 388574
rect 243822 388338 279266 388574
rect 279502 388338 279586 388574
rect 279822 388338 315266 388574
rect 315502 388338 315586 388574
rect 315822 388338 351266 388574
rect 351502 388338 351586 388574
rect 351822 388338 387266 388574
rect 387502 388338 387586 388574
rect 387822 388338 423266 388574
rect 423502 388338 423586 388574
rect 423822 388338 459266 388574
rect 459502 388338 459586 388574
rect 459822 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 95546 385174
rect 95782 384938 95866 385174
rect 96102 384938 131546 385174
rect 131782 384938 131866 385174
rect 132102 384938 167546 385174
rect 167782 384938 167866 385174
rect 168102 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 239546 385174
rect 239782 384938 239866 385174
rect 240102 384938 275546 385174
rect 275782 384938 275866 385174
rect 276102 384938 311546 385174
rect 311782 384938 311866 385174
rect 312102 384938 347546 385174
rect 347782 384938 347866 385174
rect 348102 384938 383546 385174
rect 383782 384938 383866 385174
rect 384102 384938 419546 385174
rect 419782 384938 419866 385174
rect 420102 384938 455546 385174
rect 455782 384938 455866 385174
rect 456102 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect -4886 384854 588810 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 95546 384854
rect 95782 384618 95866 384854
rect 96102 384618 131546 384854
rect 131782 384618 131866 384854
rect 132102 384618 167546 384854
rect 167782 384618 167866 384854
rect 168102 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 239546 384854
rect 239782 384618 239866 384854
rect 240102 384618 275546 384854
rect 275782 384618 275866 384854
rect 276102 384618 311546 384854
rect 311782 384618 311866 384854
rect 312102 384618 347546 384854
rect 347782 384618 347866 384854
rect 348102 384618 383546 384854
rect 383782 384618 383866 384854
rect 384102 384618 419546 384854
rect 419782 384618 419866 384854
rect 420102 384618 455546 384854
rect 455782 384618 455866 384854
rect 456102 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect -2966 381134 586890 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 592650 374294
rect -8726 374026 592650 374058
rect -6806 370894 590730 370926
rect -6806 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 590730 370894
rect -6806 370574 590730 370658
rect -6806 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 590730 370574
rect -6806 370306 590730 370338
rect -4886 367174 588810 367206
rect -4886 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 588810 367174
rect -4886 366854 588810 366938
rect -4886 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 588810 366854
rect -4886 366586 588810 366618
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect -8726 356614 592650 356646
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 102986 356614
rect 103222 356378 103306 356614
rect 103542 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 210986 356614
rect 211222 356378 211306 356614
rect 211542 356378 246986 356614
rect 247222 356378 247306 356614
rect 247542 356378 282986 356614
rect 283222 356378 283306 356614
rect 283542 356378 318986 356614
rect 319222 356378 319306 356614
rect 319542 356378 354986 356614
rect 355222 356378 355306 356614
rect 355542 356378 390986 356614
rect 391222 356378 391306 356614
rect 391542 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect -8726 356294 592650 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 102986 356294
rect 103222 356058 103306 356294
rect 103542 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 210986 356294
rect 211222 356058 211306 356294
rect 211542 356058 246986 356294
rect 247222 356058 247306 356294
rect 247542 356058 282986 356294
rect 283222 356058 283306 356294
rect 283542 356058 318986 356294
rect 319222 356058 319306 356294
rect 319542 356058 354986 356294
rect 355222 356058 355306 356294
rect 355542 356058 390986 356294
rect 391222 356058 391306 356294
rect 391542 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 99266 352894
rect 99502 352658 99586 352894
rect 99822 352658 135266 352894
rect 135502 352658 135586 352894
rect 135822 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 243266 352894
rect 243502 352658 243586 352894
rect 243822 352658 279266 352894
rect 279502 352658 279586 352894
rect 279822 352658 315266 352894
rect 315502 352658 315586 352894
rect 315822 352658 351266 352894
rect 351502 352658 351586 352894
rect 351822 352658 387266 352894
rect 387502 352658 387586 352894
rect 387822 352658 423266 352894
rect 423502 352658 423586 352894
rect 423822 352658 459266 352894
rect 459502 352658 459586 352894
rect 459822 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect -6806 352574 590730 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 99266 352574
rect 99502 352338 99586 352574
rect 99822 352338 135266 352574
rect 135502 352338 135586 352574
rect 135822 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 243266 352574
rect 243502 352338 243586 352574
rect 243822 352338 279266 352574
rect 279502 352338 279586 352574
rect 279822 352338 315266 352574
rect 315502 352338 315586 352574
rect 315822 352338 351266 352574
rect 351502 352338 351586 352574
rect 351822 352338 387266 352574
rect 387502 352338 387586 352574
rect 387822 352338 423266 352574
rect 423502 352338 423586 352574
rect 423822 352338 459266 352574
rect 459502 352338 459586 352574
rect 459822 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 95546 349174
rect 95782 348938 95866 349174
rect 96102 348938 131546 349174
rect 131782 348938 131866 349174
rect 132102 348938 167546 349174
rect 167782 348938 167866 349174
rect 168102 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 239546 349174
rect 239782 348938 239866 349174
rect 240102 348938 275546 349174
rect 275782 348938 275866 349174
rect 276102 348938 311546 349174
rect 311782 348938 311866 349174
rect 312102 348938 347546 349174
rect 347782 348938 347866 349174
rect 348102 348938 383546 349174
rect 383782 348938 383866 349174
rect 384102 348938 419546 349174
rect 419782 348938 419866 349174
rect 420102 348938 455546 349174
rect 455782 348938 455866 349174
rect 456102 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect -4886 348854 588810 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 95546 348854
rect 95782 348618 95866 348854
rect 96102 348618 131546 348854
rect 131782 348618 131866 348854
rect 132102 348618 167546 348854
rect 167782 348618 167866 348854
rect 168102 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 239546 348854
rect 239782 348618 239866 348854
rect 240102 348618 275546 348854
rect 275782 348618 275866 348854
rect 276102 348618 311546 348854
rect 311782 348618 311866 348854
rect 312102 348618 347546 348854
rect 347782 348618 347866 348854
rect 348102 348618 383546 348854
rect 383782 348618 383866 348854
rect 384102 348618 419546 348854
rect 419782 348618 419866 348854
rect 420102 348618 455546 348854
rect 455782 348618 455866 348854
rect 456102 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect -4886 348586 588810 348618
rect -2966 345454 586890 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect -2966 345134 586890 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect -2966 344866 586890 344898
rect -8726 338614 592650 338646
rect -8726 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 264986 338614
rect 265222 338378 265306 338614
rect 265542 338378 300986 338614
rect 301222 338378 301306 338614
rect 301542 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 264986 338294
rect 265222 338058 265306 338294
rect 265542 338058 300986 338294
rect 301222 338058 301306 338294
rect 301542 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 592650 338294
rect -8726 338026 592650 338058
rect -6806 334894 590730 334926
rect -6806 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 225266 334894
rect 225502 334658 225586 334894
rect 225822 334658 261266 334894
rect 261502 334658 261586 334894
rect 261822 334658 297266 334894
rect 297502 334658 297586 334894
rect 297822 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 590730 334894
rect -6806 334574 590730 334658
rect -6806 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 225266 334574
rect 225502 334338 225586 334574
rect 225822 334338 261266 334574
rect 261502 334338 261586 334574
rect 261822 334338 297266 334574
rect 297502 334338 297586 334574
rect 297822 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 590730 334574
rect -6806 334306 590730 334338
rect -4886 331174 588810 331206
rect -4886 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 257546 331174
rect 257782 330938 257866 331174
rect 258102 330938 293546 331174
rect 293782 330938 293866 331174
rect 294102 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 588810 331174
rect -4886 330854 588810 330938
rect -4886 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 257546 330854
rect 257782 330618 257866 330854
rect 258102 330618 293546 330854
rect 293782 330618 293866 330854
rect 294102 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 588810 330854
rect -4886 330586 588810 330618
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 66986 320614
rect 67222 320378 67306 320614
rect 67542 320378 102986 320614
rect 103222 320378 103306 320614
rect 103542 320378 138986 320614
rect 139222 320378 139306 320614
rect 139542 320378 174986 320614
rect 175222 320378 175306 320614
rect 175542 320378 210986 320614
rect 211222 320378 211306 320614
rect 211542 320378 246986 320614
rect 247222 320378 247306 320614
rect 247542 320378 282986 320614
rect 283222 320378 283306 320614
rect 283542 320378 318986 320614
rect 319222 320378 319306 320614
rect 319542 320378 354986 320614
rect 355222 320378 355306 320614
rect 355542 320378 390986 320614
rect 391222 320378 391306 320614
rect 391542 320378 426986 320614
rect 427222 320378 427306 320614
rect 427542 320378 462986 320614
rect 463222 320378 463306 320614
rect 463542 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect -8726 320294 592650 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 66986 320294
rect 67222 320058 67306 320294
rect 67542 320058 102986 320294
rect 103222 320058 103306 320294
rect 103542 320058 138986 320294
rect 139222 320058 139306 320294
rect 139542 320058 174986 320294
rect 175222 320058 175306 320294
rect 175542 320058 210986 320294
rect 211222 320058 211306 320294
rect 211542 320058 246986 320294
rect 247222 320058 247306 320294
rect 247542 320058 282986 320294
rect 283222 320058 283306 320294
rect 283542 320058 318986 320294
rect 319222 320058 319306 320294
rect 319542 320058 354986 320294
rect 355222 320058 355306 320294
rect 355542 320058 390986 320294
rect 391222 320058 391306 320294
rect 391542 320058 426986 320294
rect 427222 320058 427306 320294
rect 427542 320058 462986 320294
rect 463222 320058 463306 320294
rect 463542 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 99266 316894
rect 99502 316658 99586 316894
rect 99822 316658 135266 316894
rect 135502 316658 135586 316894
rect 135822 316658 171266 316894
rect 171502 316658 171586 316894
rect 171822 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 243266 316894
rect 243502 316658 243586 316894
rect 243822 316658 279266 316894
rect 279502 316658 279586 316894
rect 279822 316658 315266 316894
rect 315502 316658 315586 316894
rect 315822 316658 351266 316894
rect 351502 316658 351586 316894
rect 351822 316658 387266 316894
rect 387502 316658 387586 316894
rect 387822 316658 423266 316894
rect 423502 316658 423586 316894
rect 423822 316658 459266 316894
rect 459502 316658 459586 316894
rect 459822 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect -6806 316574 590730 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 99266 316574
rect 99502 316338 99586 316574
rect 99822 316338 135266 316574
rect 135502 316338 135586 316574
rect 135822 316338 171266 316574
rect 171502 316338 171586 316574
rect 171822 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 243266 316574
rect 243502 316338 243586 316574
rect 243822 316338 279266 316574
rect 279502 316338 279586 316574
rect 279822 316338 315266 316574
rect 315502 316338 315586 316574
rect 315822 316338 351266 316574
rect 351502 316338 351586 316574
rect 351822 316338 387266 316574
rect 387502 316338 387586 316574
rect 387822 316338 423266 316574
rect 423502 316338 423586 316574
rect 423822 316338 459266 316574
rect 459502 316338 459586 316574
rect 459822 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 95546 313174
rect 95782 312938 95866 313174
rect 96102 312938 131546 313174
rect 131782 312938 131866 313174
rect 132102 312938 167546 313174
rect 167782 312938 167866 313174
rect 168102 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 239546 313174
rect 239782 312938 239866 313174
rect 240102 312938 275546 313174
rect 275782 312938 275866 313174
rect 276102 312938 311546 313174
rect 311782 312938 311866 313174
rect 312102 312938 347546 313174
rect 347782 312938 347866 313174
rect 348102 312938 383546 313174
rect 383782 312938 383866 313174
rect 384102 312938 419546 313174
rect 419782 312938 419866 313174
rect 420102 312938 455546 313174
rect 455782 312938 455866 313174
rect 456102 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect -4886 312854 588810 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 95546 312854
rect 95782 312618 95866 312854
rect 96102 312618 131546 312854
rect 131782 312618 131866 312854
rect 132102 312618 167546 312854
rect 167782 312618 167866 312854
rect 168102 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 239546 312854
rect 239782 312618 239866 312854
rect 240102 312618 275546 312854
rect 275782 312618 275866 312854
rect 276102 312618 311546 312854
rect 311782 312618 311866 312854
rect 312102 312618 347546 312854
rect 347782 312618 347866 312854
rect 348102 312618 383546 312854
rect 383782 312618 383866 312854
rect 384102 312618 419546 312854
rect 419782 312618 419866 312854
rect 420102 312618 455546 312854
rect 455782 312618 455866 312854
rect 456102 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect -2966 309134 586890 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect -2966 308866 586890 308898
rect -8726 302614 592650 302646
rect -8726 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 192986 302614
rect 193222 302378 193306 302614
rect 193542 302378 228986 302614
rect 229222 302378 229306 302614
rect 229542 302378 264986 302614
rect 265222 302378 265306 302614
rect 265542 302378 300986 302614
rect 301222 302378 301306 302614
rect 301542 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 192986 302294
rect 193222 302058 193306 302294
rect 193542 302058 228986 302294
rect 229222 302058 229306 302294
rect 229542 302058 264986 302294
rect 265222 302058 265306 302294
rect 265542 302058 300986 302294
rect 301222 302058 301306 302294
rect 301542 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 592650 302294
rect -8726 302026 592650 302058
rect -6806 298894 590730 298926
rect -6806 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 81266 298894
rect 81502 298658 81586 298894
rect 81822 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 225266 298894
rect 225502 298658 225586 298894
rect 225822 298658 261266 298894
rect 261502 298658 261586 298894
rect 261822 298658 297266 298894
rect 297502 298658 297586 298894
rect 297822 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 590730 298894
rect -6806 298574 590730 298658
rect -6806 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 81266 298574
rect 81502 298338 81586 298574
rect 81822 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 225266 298574
rect 225502 298338 225586 298574
rect 225822 298338 261266 298574
rect 261502 298338 261586 298574
rect 261822 298338 297266 298574
rect 297502 298338 297586 298574
rect 297822 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 590730 298574
rect -6806 298306 590730 298338
rect -4886 295174 588810 295206
rect -4886 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 221546 295174
rect 221782 294938 221866 295174
rect 222102 294938 257546 295174
rect 257782 294938 257866 295174
rect 258102 294938 293546 295174
rect 293782 294938 293866 295174
rect 294102 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 588810 295174
rect -4886 294854 588810 294938
rect -4886 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 221546 294854
rect 221782 294618 221866 294854
rect 222102 294618 257546 294854
rect 257782 294618 257866 294854
rect 258102 294618 293546 294854
rect 293782 294618 293866 294854
rect 294102 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 588810 294854
rect -4886 294586 588810 294618
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 66986 284614
rect 67222 284378 67306 284614
rect 67542 284378 102986 284614
rect 103222 284378 103306 284614
rect 103542 284378 138986 284614
rect 139222 284378 139306 284614
rect 139542 284378 174986 284614
rect 175222 284378 175306 284614
rect 175542 284378 210986 284614
rect 211222 284378 211306 284614
rect 211542 284378 246986 284614
rect 247222 284378 247306 284614
rect 247542 284378 282986 284614
rect 283222 284378 283306 284614
rect 283542 284378 318986 284614
rect 319222 284378 319306 284614
rect 319542 284378 354986 284614
rect 355222 284378 355306 284614
rect 355542 284378 390986 284614
rect 391222 284378 391306 284614
rect 391542 284378 426986 284614
rect 427222 284378 427306 284614
rect 427542 284378 462986 284614
rect 463222 284378 463306 284614
rect 463542 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect -8726 284294 592650 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 66986 284294
rect 67222 284058 67306 284294
rect 67542 284058 102986 284294
rect 103222 284058 103306 284294
rect 103542 284058 138986 284294
rect 139222 284058 139306 284294
rect 139542 284058 174986 284294
rect 175222 284058 175306 284294
rect 175542 284058 210986 284294
rect 211222 284058 211306 284294
rect 211542 284058 246986 284294
rect 247222 284058 247306 284294
rect 247542 284058 282986 284294
rect 283222 284058 283306 284294
rect 283542 284058 318986 284294
rect 319222 284058 319306 284294
rect 319542 284058 354986 284294
rect 355222 284058 355306 284294
rect 355542 284058 390986 284294
rect 391222 284058 391306 284294
rect 391542 284058 426986 284294
rect 427222 284058 427306 284294
rect 427542 284058 462986 284294
rect 463222 284058 463306 284294
rect 463542 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 99266 280894
rect 99502 280658 99586 280894
rect 99822 280658 135266 280894
rect 135502 280658 135586 280894
rect 135822 280658 171266 280894
rect 171502 280658 171586 280894
rect 171822 280658 207266 280894
rect 207502 280658 207586 280894
rect 207822 280658 243266 280894
rect 243502 280658 243586 280894
rect 243822 280658 279266 280894
rect 279502 280658 279586 280894
rect 279822 280658 315266 280894
rect 315502 280658 315586 280894
rect 315822 280658 351266 280894
rect 351502 280658 351586 280894
rect 351822 280658 387266 280894
rect 387502 280658 387586 280894
rect 387822 280658 423266 280894
rect 423502 280658 423586 280894
rect 423822 280658 459266 280894
rect 459502 280658 459586 280894
rect 459822 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect -6806 280574 590730 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 99266 280574
rect 99502 280338 99586 280574
rect 99822 280338 135266 280574
rect 135502 280338 135586 280574
rect 135822 280338 171266 280574
rect 171502 280338 171586 280574
rect 171822 280338 207266 280574
rect 207502 280338 207586 280574
rect 207822 280338 243266 280574
rect 243502 280338 243586 280574
rect 243822 280338 279266 280574
rect 279502 280338 279586 280574
rect 279822 280338 315266 280574
rect 315502 280338 315586 280574
rect 315822 280338 351266 280574
rect 351502 280338 351586 280574
rect 351822 280338 387266 280574
rect 387502 280338 387586 280574
rect 387822 280338 423266 280574
rect 423502 280338 423586 280574
rect 423822 280338 459266 280574
rect 459502 280338 459586 280574
rect 459822 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 95546 277174
rect 95782 276938 95866 277174
rect 96102 276938 131546 277174
rect 131782 276938 131866 277174
rect 132102 276938 167546 277174
rect 167782 276938 167866 277174
rect 168102 276938 203546 277174
rect 203782 276938 203866 277174
rect 204102 276938 239546 277174
rect 239782 276938 239866 277174
rect 240102 276938 275546 277174
rect 275782 276938 275866 277174
rect 276102 276938 311546 277174
rect 311782 276938 311866 277174
rect 312102 276938 347546 277174
rect 347782 276938 347866 277174
rect 348102 276938 383546 277174
rect 383782 276938 383866 277174
rect 384102 276938 419546 277174
rect 419782 276938 419866 277174
rect 420102 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect -4886 276854 588810 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 95546 276854
rect 95782 276618 95866 276854
rect 96102 276618 131546 276854
rect 131782 276618 131866 276854
rect 132102 276618 167546 276854
rect 167782 276618 167866 276854
rect 168102 276618 203546 276854
rect 203782 276618 203866 276854
rect 204102 276618 239546 276854
rect 239782 276618 239866 276854
rect 240102 276618 275546 276854
rect 275782 276618 275866 276854
rect 276102 276618 311546 276854
rect 311782 276618 311866 276854
rect 312102 276618 347546 276854
rect 347782 276618 347866 276854
rect 348102 276618 383546 276854
rect 383782 276618 383866 276854
rect 384102 276618 419546 276854
rect 419782 276618 419866 276854
rect 420102 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect -4886 276586 588810 276618
rect -2966 273454 586890 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect -2966 273134 586890 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 84986 266614
rect 85222 266378 85306 266614
rect 85542 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 228986 266614
rect 229222 266378 229306 266614
rect 229542 266378 264986 266614
rect 265222 266378 265306 266614
rect 265542 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 84986 266294
rect 85222 266058 85306 266294
rect 85542 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 228986 266294
rect 229222 266058 229306 266294
rect 229542 266058 264986 266294
rect 265222 266058 265306 266294
rect 265542 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 592650 266294
rect -8726 266026 592650 266058
rect -6806 262894 590730 262926
rect -6806 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 81266 262894
rect 81502 262658 81586 262894
rect 81822 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 225266 262894
rect 225502 262658 225586 262894
rect 225822 262658 261266 262894
rect 261502 262658 261586 262894
rect 261822 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 590730 262894
rect -6806 262574 590730 262658
rect -6806 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 81266 262574
rect 81502 262338 81586 262574
rect 81822 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 225266 262574
rect 225502 262338 225586 262574
rect 225822 262338 261266 262574
rect 261502 262338 261586 262574
rect 261822 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 590730 262574
rect -6806 262306 590730 262338
rect -4886 259174 588810 259206
rect -4886 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 77546 259174
rect 77782 258938 77866 259174
rect 78102 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 221546 259174
rect 221782 258938 221866 259174
rect 222102 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 588810 259174
rect -4886 258854 588810 258938
rect -4886 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 77546 258854
rect 77782 258618 77866 258854
rect 78102 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 221546 258854
rect 221782 258618 221866 258854
rect 222102 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 588810 258854
rect -4886 258586 588810 258618
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -8726 248614 592650 248646
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 66986 248614
rect 67222 248378 67306 248614
rect 67542 248378 102986 248614
rect 103222 248378 103306 248614
rect 103542 248378 138986 248614
rect 139222 248378 139306 248614
rect 139542 248378 174986 248614
rect 175222 248378 175306 248614
rect 175542 248378 210986 248614
rect 211222 248378 211306 248614
rect 211542 248378 246986 248614
rect 247222 248378 247306 248614
rect 247542 248378 282986 248614
rect 283222 248378 283306 248614
rect 283542 248378 318986 248614
rect 319222 248378 319306 248614
rect 319542 248378 354986 248614
rect 355222 248378 355306 248614
rect 355542 248378 390986 248614
rect 391222 248378 391306 248614
rect 391542 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect -8726 248294 592650 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 66986 248294
rect 67222 248058 67306 248294
rect 67542 248058 102986 248294
rect 103222 248058 103306 248294
rect 103542 248058 138986 248294
rect 139222 248058 139306 248294
rect 139542 248058 174986 248294
rect 175222 248058 175306 248294
rect 175542 248058 210986 248294
rect 211222 248058 211306 248294
rect 211542 248058 246986 248294
rect 247222 248058 247306 248294
rect 247542 248058 282986 248294
rect 283222 248058 283306 248294
rect 283542 248058 318986 248294
rect 319222 248058 319306 248294
rect 319542 248058 354986 248294
rect 355222 248058 355306 248294
rect 355542 248058 390986 248294
rect 391222 248058 391306 248294
rect 391542 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 99266 244894
rect 99502 244658 99586 244894
rect 99822 244658 135266 244894
rect 135502 244658 135586 244894
rect 135822 244658 171266 244894
rect 171502 244658 171586 244894
rect 171822 244658 207266 244894
rect 207502 244658 207586 244894
rect 207822 244658 243266 244894
rect 243502 244658 243586 244894
rect 243822 244658 279266 244894
rect 279502 244658 279586 244894
rect 279822 244658 315266 244894
rect 315502 244658 315586 244894
rect 315822 244658 351266 244894
rect 351502 244658 351586 244894
rect 351822 244658 387266 244894
rect 387502 244658 387586 244894
rect 387822 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect -6806 244574 590730 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 99266 244574
rect 99502 244338 99586 244574
rect 99822 244338 135266 244574
rect 135502 244338 135586 244574
rect 135822 244338 171266 244574
rect 171502 244338 171586 244574
rect 171822 244338 207266 244574
rect 207502 244338 207586 244574
rect 207822 244338 243266 244574
rect 243502 244338 243586 244574
rect 243822 244338 279266 244574
rect 279502 244338 279586 244574
rect 279822 244338 315266 244574
rect 315502 244338 315586 244574
rect 315822 244338 351266 244574
rect 351502 244338 351586 244574
rect 351822 244338 387266 244574
rect 387502 244338 387586 244574
rect 387822 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 95546 241174
rect 95782 240938 95866 241174
rect 96102 240938 131546 241174
rect 131782 240938 131866 241174
rect 132102 240938 167546 241174
rect 167782 240938 167866 241174
rect 168102 240938 203546 241174
rect 203782 240938 203866 241174
rect 204102 240938 239546 241174
rect 239782 240938 239866 241174
rect 240102 240938 275546 241174
rect 275782 240938 275866 241174
rect 276102 240938 311546 241174
rect 311782 240938 311866 241174
rect 312102 240938 347546 241174
rect 347782 240938 347866 241174
rect 348102 240938 383546 241174
rect 383782 240938 383866 241174
rect 384102 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect -4886 240854 588810 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 95546 240854
rect 95782 240618 95866 240854
rect 96102 240618 131546 240854
rect 131782 240618 131866 240854
rect 132102 240618 167546 240854
rect 167782 240618 167866 240854
rect 168102 240618 203546 240854
rect 203782 240618 203866 240854
rect 204102 240618 239546 240854
rect 239782 240618 239866 240854
rect 240102 240618 275546 240854
rect 275782 240618 275866 240854
rect 276102 240618 311546 240854
rect 311782 240618 311866 240854
rect 312102 240618 347546 240854
rect 347782 240618 347866 240854
rect 348102 240618 383546 240854
rect 383782 240618 383866 240854
rect 384102 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect -2966 237134 586890 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 228986 230614
rect 229222 230378 229306 230614
rect 229542 230378 264986 230614
rect 265222 230378 265306 230614
rect 265542 230378 300986 230614
rect 301222 230378 301306 230614
rect 301542 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 228986 230294
rect 229222 230058 229306 230294
rect 229542 230058 264986 230294
rect 265222 230058 265306 230294
rect 265542 230058 300986 230294
rect 301222 230058 301306 230294
rect 301542 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 592650 230294
rect -8726 230026 592650 230058
rect -6806 226894 590730 226926
rect -6806 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 261266 226894
rect 261502 226658 261586 226894
rect 261822 226658 297266 226894
rect 297502 226658 297586 226894
rect 297822 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 590730 226894
rect -6806 226574 590730 226658
rect -6806 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 261266 226574
rect 261502 226338 261586 226574
rect 261822 226338 297266 226574
rect 297502 226338 297586 226574
rect 297822 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 590730 226574
rect -6806 226306 590730 226338
rect -4886 223174 588810 223206
rect -4886 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 257546 223174
rect 257782 222938 257866 223174
rect 258102 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 588810 223174
rect -4886 222854 588810 222938
rect -4886 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 257546 222854
rect 257782 222618 257866 222854
rect 258102 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 588810 222854
rect -4886 222586 588810 222618
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 64250 219454
rect 64486 219218 94970 219454
rect 95206 219218 125690 219454
rect 125926 219218 156410 219454
rect 156646 219218 187130 219454
rect 187366 219218 217850 219454
rect 218086 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 64250 219134
rect 64486 218898 94970 219134
rect 95206 218898 125690 219134
rect 125926 218898 156410 219134
rect 156646 218898 187130 219134
rect 187366 218898 217850 219134
rect 218086 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -8726 212614 592650 212646
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 246986 212614
rect 247222 212378 247306 212614
rect 247542 212378 282986 212614
rect 283222 212378 283306 212614
rect 283542 212378 318986 212614
rect 319222 212378 319306 212614
rect 319542 212378 354986 212614
rect 355222 212378 355306 212614
rect 355542 212378 390986 212614
rect 391222 212378 391306 212614
rect 391542 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect -8726 212294 592650 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 246986 212294
rect 247222 212058 247306 212294
rect 247542 212058 282986 212294
rect 283222 212058 283306 212294
rect 283542 212058 318986 212294
rect 319222 212058 319306 212294
rect 319542 212058 354986 212294
rect 355222 212058 355306 212294
rect 355542 212058 390986 212294
rect 391222 212058 391306 212294
rect 391542 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 243266 208894
rect 243502 208658 243586 208894
rect 243822 208658 279266 208894
rect 279502 208658 279586 208894
rect 279822 208658 315266 208894
rect 315502 208658 315586 208894
rect 315822 208658 351266 208894
rect 351502 208658 351586 208894
rect 351822 208658 387266 208894
rect 387502 208658 387586 208894
rect 387822 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect -6806 208574 590730 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 243266 208574
rect 243502 208338 243586 208574
rect 243822 208338 279266 208574
rect 279502 208338 279586 208574
rect 279822 208338 315266 208574
rect 315502 208338 315586 208574
rect 315822 208338 351266 208574
rect 351502 208338 351586 208574
rect 351822 208338 387266 208574
rect 387502 208338 387586 208574
rect 387822 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 239546 205174
rect 239782 204938 239866 205174
rect 240102 204938 275546 205174
rect 275782 204938 275866 205174
rect 276102 204938 311546 205174
rect 311782 204938 311866 205174
rect 312102 204938 347546 205174
rect 347782 204938 347866 205174
rect 348102 204938 383546 205174
rect 383782 204938 383866 205174
rect 384102 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect -4886 204854 588810 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 239546 204854
rect 239782 204618 239866 204854
rect 240102 204618 275546 204854
rect 275782 204618 275866 204854
rect 276102 204618 311546 204854
rect 311782 204618 311866 204854
rect 312102 204618 347546 204854
rect 347782 204618 347866 204854
rect 348102 204618 383546 204854
rect 383782 204618 383866 204854
rect 384102 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 79610 201454
rect 79846 201218 110330 201454
rect 110566 201218 141050 201454
rect 141286 201218 171770 201454
rect 172006 201218 202490 201454
rect 202726 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect -2966 201134 586890 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 79610 201134
rect 79846 200898 110330 201134
rect 110566 200898 141050 201134
rect 141286 200898 171770 201134
rect 172006 200898 202490 201134
rect 202726 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 264986 194614
rect 265222 194378 265306 194614
rect 265542 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 264986 194294
rect 265222 194058 265306 194294
rect 265542 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 592650 194294
rect -8726 194026 592650 194058
rect -6806 190894 590730 190926
rect -6806 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 261266 190894
rect 261502 190658 261586 190894
rect 261822 190658 297266 190894
rect 297502 190658 297586 190894
rect 297822 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 590730 190894
rect -6806 190574 590730 190658
rect -6806 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 261266 190574
rect 261502 190338 261586 190574
rect 261822 190338 297266 190574
rect 297502 190338 297586 190574
rect 297822 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 590730 190574
rect -6806 190306 590730 190338
rect -4886 187174 588810 187206
rect -4886 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 257546 187174
rect 257782 186938 257866 187174
rect 258102 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 588810 187174
rect -4886 186854 588810 186938
rect -4886 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 257546 186854
rect 257782 186618 257866 186854
rect 258102 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 588810 186854
rect -4886 186586 588810 186618
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 64250 183454
rect 64486 183218 94970 183454
rect 95206 183218 125690 183454
rect 125926 183218 156410 183454
rect 156646 183218 187130 183454
rect 187366 183218 217850 183454
rect 218086 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 64250 183134
rect 64486 182898 94970 183134
rect 95206 182898 125690 183134
rect 125926 182898 156410 183134
rect 156646 182898 187130 183134
rect 187366 182898 217850 183134
rect 218086 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect -8726 176614 592650 176646
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 246986 176614
rect 247222 176378 247306 176614
rect 247542 176378 282986 176614
rect 283222 176378 283306 176614
rect 283542 176378 318986 176614
rect 319222 176378 319306 176614
rect 319542 176378 354986 176614
rect 355222 176378 355306 176614
rect 355542 176378 390986 176614
rect 391222 176378 391306 176614
rect 391542 176378 426986 176614
rect 427222 176378 427306 176614
rect 427542 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect -8726 176294 592650 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 246986 176294
rect 247222 176058 247306 176294
rect 247542 176058 282986 176294
rect 283222 176058 283306 176294
rect 283542 176058 318986 176294
rect 319222 176058 319306 176294
rect 319542 176058 354986 176294
rect 355222 176058 355306 176294
rect 355542 176058 390986 176294
rect 391222 176058 391306 176294
rect 391542 176058 426986 176294
rect 427222 176058 427306 176294
rect 427542 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect -8726 176026 592650 176058
rect -6806 172894 590730 172926
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 243266 172894
rect 243502 172658 243586 172894
rect 243822 172658 279266 172894
rect 279502 172658 279586 172894
rect 279822 172658 315266 172894
rect 315502 172658 315586 172894
rect 315822 172658 351266 172894
rect 351502 172658 351586 172894
rect 351822 172658 387266 172894
rect 387502 172658 387586 172894
rect 387822 172658 423266 172894
rect 423502 172658 423586 172894
rect 423822 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect -6806 172574 590730 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 243266 172574
rect 243502 172338 243586 172574
rect 243822 172338 279266 172574
rect 279502 172338 279586 172574
rect 279822 172338 315266 172574
rect 315502 172338 315586 172574
rect 315822 172338 351266 172574
rect 351502 172338 351586 172574
rect 351822 172338 387266 172574
rect 387502 172338 387586 172574
rect 387822 172338 423266 172574
rect 423502 172338 423586 172574
rect 423822 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect -6806 172306 590730 172338
rect -4886 169174 588810 169206
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 239546 169174
rect 239782 168938 239866 169174
rect 240102 168938 275546 169174
rect 275782 168938 275866 169174
rect 276102 168938 311546 169174
rect 311782 168938 311866 169174
rect 312102 168938 347546 169174
rect 347782 168938 347866 169174
rect 348102 168938 383546 169174
rect 383782 168938 383866 169174
rect 384102 168938 419546 169174
rect 419782 168938 419866 169174
rect 420102 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect -4886 168854 588810 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 239546 168854
rect 239782 168618 239866 168854
rect 240102 168618 275546 168854
rect 275782 168618 275866 168854
rect 276102 168618 311546 168854
rect 311782 168618 311866 168854
rect 312102 168618 347546 168854
rect 347782 168618 347866 168854
rect 348102 168618 383546 168854
rect 383782 168618 383866 168854
rect 384102 168618 419546 168854
rect 419782 168618 419866 168854
rect 420102 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect -4886 168586 588810 168618
rect -2966 165454 586890 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 79610 165454
rect 79846 165218 110330 165454
rect 110566 165218 141050 165454
rect 141286 165218 171770 165454
rect 172006 165218 202490 165454
rect 202726 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect -2966 165134 586890 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 79610 165134
rect 79846 164898 110330 165134
rect 110566 164898 141050 165134
rect 141286 164898 171770 165134
rect 172006 164898 202490 165134
rect 202726 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect -2966 164866 586890 164898
rect -8726 158614 592650 158646
rect -8726 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 228986 158614
rect 229222 158378 229306 158614
rect 229542 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 228986 158294
rect 229222 158058 229306 158294
rect 229542 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 592650 158294
rect -8726 158026 592650 158058
rect -6806 154894 590730 154926
rect -6806 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 590730 154894
rect -6806 154574 590730 154658
rect -6806 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 590730 154574
rect -6806 154306 590730 154338
rect -4886 151174 588810 151206
rect -4886 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 588810 151174
rect -4886 150854 588810 150938
rect -4886 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 588810 150854
rect -4886 150586 588810 150618
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 64250 147454
rect 64486 147218 94970 147454
rect 95206 147218 125690 147454
rect 125926 147218 156410 147454
rect 156646 147218 187130 147454
rect 187366 147218 217850 147454
rect 218086 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 64250 147134
rect 64486 146898 94970 147134
rect 95206 146898 125690 147134
rect 125926 146898 156410 147134
rect 156646 146898 187130 147134
rect 187366 146898 217850 147134
rect 218086 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -8726 140614 592650 140646
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 246986 140614
rect 247222 140378 247306 140614
rect 247542 140378 282986 140614
rect 283222 140378 283306 140614
rect 283542 140378 318986 140614
rect 319222 140378 319306 140614
rect 319542 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 426986 140614
rect 427222 140378 427306 140614
rect 427542 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect -8726 140294 592650 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 246986 140294
rect 247222 140058 247306 140294
rect 247542 140058 282986 140294
rect 283222 140058 283306 140294
rect 283542 140058 318986 140294
rect 319222 140058 319306 140294
rect 319542 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 426986 140294
rect 427222 140058 427306 140294
rect 427542 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect -8726 140026 592650 140058
rect -6806 136894 590730 136926
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 243266 136894
rect 243502 136658 243586 136894
rect 243822 136658 279266 136894
rect 279502 136658 279586 136894
rect 279822 136658 315266 136894
rect 315502 136658 315586 136894
rect 315822 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 423266 136894
rect 423502 136658 423586 136894
rect 423822 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect -6806 136574 590730 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 243266 136574
rect 243502 136338 243586 136574
rect 243822 136338 279266 136574
rect 279502 136338 279586 136574
rect 279822 136338 315266 136574
rect 315502 136338 315586 136574
rect 315822 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 423266 136574
rect 423502 136338 423586 136574
rect 423822 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect -6806 136306 590730 136338
rect -4886 133174 588810 133206
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 239546 133174
rect 239782 132938 239866 133174
rect 240102 132938 275546 133174
rect 275782 132938 275866 133174
rect 276102 132938 311546 133174
rect 311782 132938 311866 133174
rect 312102 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 419546 133174
rect 419782 132938 419866 133174
rect 420102 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect -4886 132854 588810 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 239546 132854
rect 239782 132618 239866 132854
rect 240102 132618 275546 132854
rect 275782 132618 275866 132854
rect 276102 132618 311546 132854
rect 311782 132618 311866 132854
rect 312102 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 419546 132854
rect 419782 132618 419866 132854
rect 420102 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect -4886 132586 588810 132618
rect -2966 129454 586890 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 79610 129454
rect 79846 129218 110330 129454
rect 110566 129218 141050 129454
rect 141286 129218 171770 129454
rect 172006 129218 202490 129454
rect 202726 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect -2966 129134 586890 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 79610 129134
rect 79846 128898 110330 129134
rect 110566 128898 141050 129134
rect 141286 128898 171770 129134
rect 172006 128898 202490 129134
rect 202726 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect -2966 128866 586890 128898
rect -8726 122614 592650 122646
rect -8726 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 228986 122614
rect 229222 122378 229306 122614
rect 229542 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 228986 122294
rect 229222 122058 229306 122294
rect 229542 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 592650 122294
rect -8726 122026 592650 122058
rect -6806 118894 590730 118926
rect -6806 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 590730 118894
rect -6806 118574 590730 118658
rect -6806 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 590730 118574
rect -6806 118306 590730 118338
rect -4886 115174 588810 115206
rect -4886 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 588810 115174
rect -4886 114854 588810 114938
rect -4886 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 588810 114854
rect -4886 114586 588810 114618
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 64250 111454
rect 64486 111218 94970 111454
rect 95206 111218 125690 111454
rect 125926 111218 156410 111454
rect 156646 111218 187130 111454
rect 187366 111218 217850 111454
rect 218086 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 64250 111134
rect 64486 110898 94970 111134
rect 95206 110898 125690 111134
rect 125926 110898 156410 111134
rect 156646 110898 187130 111134
rect 187366 110898 217850 111134
rect 218086 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -8726 104614 592650 104646
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 246986 104614
rect 247222 104378 247306 104614
rect 247542 104378 282986 104614
rect 283222 104378 283306 104614
rect 283542 104378 318986 104614
rect 319222 104378 319306 104614
rect 319542 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 426986 104614
rect 427222 104378 427306 104614
rect 427542 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect -8726 104294 592650 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 246986 104294
rect 247222 104058 247306 104294
rect 247542 104058 282986 104294
rect 283222 104058 283306 104294
rect 283542 104058 318986 104294
rect 319222 104058 319306 104294
rect 319542 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 426986 104294
rect 427222 104058 427306 104294
rect 427542 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect -8726 104026 592650 104058
rect -6806 100894 590730 100926
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 243266 100894
rect 243502 100658 243586 100894
rect 243822 100658 279266 100894
rect 279502 100658 279586 100894
rect 279822 100658 315266 100894
rect 315502 100658 315586 100894
rect 315822 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 423266 100894
rect 423502 100658 423586 100894
rect 423822 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect -6806 100574 590730 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 243266 100574
rect 243502 100338 243586 100574
rect 243822 100338 279266 100574
rect 279502 100338 279586 100574
rect 279822 100338 315266 100574
rect 315502 100338 315586 100574
rect 315822 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 423266 100574
rect 423502 100338 423586 100574
rect 423822 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect -6806 100306 590730 100338
rect -4886 97174 588810 97206
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 239546 97174
rect 239782 96938 239866 97174
rect 240102 96938 275546 97174
rect 275782 96938 275866 97174
rect 276102 96938 311546 97174
rect 311782 96938 311866 97174
rect 312102 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect -4886 96854 588810 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 239546 96854
rect 239782 96618 239866 96854
rect 240102 96618 275546 96854
rect 275782 96618 275866 96854
rect 276102 96618 311546 96854
rect 311782 96618 311866 96854
rect 312102 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect -4886 96586 588810 96618
rect -2966 93454 586890 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 79610 93454
rect 79846 93218 110330 93454
rect 110566 93218 141050 93454
rect 141286 93218 171770 93454
rect 172006 93218 202490 93454
rect 202726 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect -2966 93134 586890 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 79610 93134
rect 79846 92898 110330 93134
rect 110566 92898 141050 93134
rect 141286 92898 171770 93134
rect 172006 92898 202490 93134
rect 202726 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect -2966 92866 586890 92898
rect -8726 86614 592650 86646
rect -8726 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 592650 86294
rect -8726 86026 592650 86058
rect -6806 82894 590730 82926
rect -6806 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 590730 82894
rect -6806 82574 590730 82658
rect -6806 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 590730 82574
rect -6806 82306 590730 82338
rect -4886 79174 588810 79206
rect -4886 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 588810 79174
rect -4886 78854 588810 78938
rect -4886 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 588810 78854
rect -4886 78586 588810 78618
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 64250 75454
rect 64486 75218 94970 75454
rect 95206 75218 125690 75454
rect 125926 75218 156410 75454
rect 156646 75218 187130 75454
rect 187366 75218 217850 75454
rect 218086 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 64250 75134
rect 64486 74898 94970 75134
rect 95206 74898 125690 75134
rect 125926 74898 156410 75134
rect 156646 74898 187130 75134
rect 187366 74898 217850 75134
rect 218086 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -8726 68614 592650 68646
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect -8726 68294 592650 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect -8726 68026 592650 68058
rect -6806 64894 590730 64926
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect -6806 64574 590730 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect -6806 64306 590730 64338
rect -4886 61174 588810 61206
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect -4886 60854 588810 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect -4886 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 592650 50294
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 590730 46894
rect -6806 46574 590730 46658
rect -6806 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 590730 46574
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 588810 43174
rect -4886 42854 588810 42938
rect -4886 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 588810 42854
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect -8726 32294 592650 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect -6806 28574 590730 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect -4886 24854 588810 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 592650 14294
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 590730 10894
rect -6806 10574 590730 10658
rect -6806 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 590730 10574
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 588810 7174
rect -4886 6854 588810 6938
rect -4886 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 588810 6854
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use sky130_sram_2kbyte_1rw1r_32x512_8  sram1
timestamp 1640373242
transform 1 0 220000 0 1 400000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  sram
timestamp 1640373242
transform 1 0 60000 0 1 400000
box 0 0 136620 83308
use user_proj  mprj
timestamp 1640373242
transform 1 0 60000 0 1 60000
box 0 0 164531 166675
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 -1894 74414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 -1894 110414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 -1894 146414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 -1894 182414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 -1894 218414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 228675 74414 398000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 228675 110414 398000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 228675 146414 398000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 228675 182414 398000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 228675 218414 398000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 -1894 254414 398000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 -1894 290414 398000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 -1894 326414 398000 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 -1894 38414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 485308 74414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 485308 110414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 485308 146414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 485308 182414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 485308 218414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 485308 254414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 485308 290414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 485308 326414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 -1894 362414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 -1894 398414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 -1894 434414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 -1894 470414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 -1894 506414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 -1894 542414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 -3814 78134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 -3814 114134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 -3814 150134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 -3814 186134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 -3814 222134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 228675 78134 398000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 228675 114134 398000 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 228675 150134 398000 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 228675 186134 398000 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 228675 222134 398000 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 -3814 258134 398000 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 -3814 294134 398000 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 -3814 330134 398000 6 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 -3814 42134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 485308 78134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 485308 114134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 485308 150134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 485308 186134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 485308 222134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 485308 258134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 485308 294134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 485308 330134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 -3814 366134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 -3814 402134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 -3814 438134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 -3814 474134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 -3814 510134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 -3814 546134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 581514 -3814 582134 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 -5734 81854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 -5734 117854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 -5734 153854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 -5734 189854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 -5734 225854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 228675 81854 398000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 228675 117854 398000 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 228675 153854 398000 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 228675 189854 398000 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 228675 225854 398000 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 -5734 261854 398000 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 -5734 297854 398000 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 -5734 333854 398000 6 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 -5734 45854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 485308 81854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 485308 117854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 485308 153854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 485308 189854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 485308 225854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 485308 261854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 485308 297854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 485308 333854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 -5734 369854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 -5734 405854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 -5734 441854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 -5734 477854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 -5734 513854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 -5734 549854 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 -7654 85574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 -7654 121574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 -7654 157574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 -7654 193574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 228675 85574 398000 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 228675 121574 398000 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 228675 157574 398000 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 228675 193574 398000 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 -7654 229574 398000 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 -7654 265574 398000 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 -7654 301574 398000 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 -7654 337574 398000 6 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 -7654 13574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 -7654 49574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 485308 85574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 485308 121574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 485308 157574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 485308 193574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 485308 229574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 485308 265574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 485308 301574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 485308 337574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 -7654 373574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 -7654 409574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 -7654 445574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 -7654 481574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 -7654 517574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 -7654 553574 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 -5734 63854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 -5734 99854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 -5734 135854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 -5734 171854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 -5734 207854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 228675 63854 398000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 228675 99854 398000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 228675 135854 398000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 228675 171854 398000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 -5734 243854 398000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 -5734 279854 398000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 -5734 315854 398000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 -5734 351854 398000 6 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 -5734 27854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 485308 63854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 485308 99854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 485308 135854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 485308 171854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 228675 207854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 485308 243854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 485308 279854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 485308 315854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 485308 351854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 -5734 387854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 -5734 423854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 -5734 459854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 -5734 495854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 -5734 531854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 -5734 567854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 -7654 67574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 -7654 103574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 -7654 139574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 -7654 175574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 -7654 211574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 228675 67574 398000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 228675 103574 398000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 228675 139574 398000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 228675 175574 398000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 -7654 247574 398000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 -7654 283574 398000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 -7654 319574 398000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 -7654 355574 398000 6 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 -7654 31574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 485308 67574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 485308 103574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 485308 139574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 485308 175574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 228675 211574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 485308 247574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 485308 283574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 485308 319574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 485308 355574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 -7654 391574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 -7654 427574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 -7654 463574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 -7654 499574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 -7654 535574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 -7654 571574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 -1894 92414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 -1894 128414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 -1894 164414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 -1894 200414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 228675 92414 398000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 228675 128414 398000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 228675 164414 398000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 -1894 236414 398000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 -1894 272414 398000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 -1894 308414 398000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 -1894 344414 398000 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 -1894 20414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 -1894 56414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 485308 92414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 485308 128414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 485308 164414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 228675 200414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 485308 236414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 485308 272414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 485308 308414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 485308 344414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 -1894 380414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 -1894 416414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 -1894 452414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 -1894 488414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 -1894 524414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 -1894 560414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 -3814 60134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 -3814 96134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 -3814 132134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 -3814 168134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 -3814 204134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 228675 60134 398000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 228675 96134 398000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 228675 132134 398000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 228675 168134 398000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 -3814 240134 398000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 -3814 276134 398000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 -3814 312134 398000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 -3814 348134 398000 6 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 -3814 24134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 485308 60134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 485308 96134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 485308 132134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 485308 168134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 228675 204134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 485308 240134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 485308 276134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 485308 312134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 485308 348134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 -3814 384134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 -3814 420134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 -3814 456134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 -3814 492134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 -3814 528134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 -3814 564134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
