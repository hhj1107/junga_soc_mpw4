magic
tech sky130A
magscale 1 2
timestamp 1639754316
<< locali >>
rect 50905 697595 50939 699397
rect 65625 698343 65659 699397
rect 80161 698411 80195 699397
rect 95157 698479 95191 699397
rect 109877 698547 109911 699397
rect 114569 698615 114603 699397
rect 124597 698683 124631 699397
rect 139317 698819 139351 699397
rect 144285 698751 144319 699397
rect 168849 698955 168883 699397
rect 173725 698887 173759 699397
rect 211261 699227 211295 699397
rect 394157 699023 394191 699329
rect 462881 697799 462915 699329
rect 492597 697731 492631 699329
rect 521853 697663 521887 699329
rect 7481 527 7515 697
rect 240517 595 240551 697
rect 255513 323 255547 629
rect 298419 629 298569 663
rect 279617 459 279651 561
rect 279709 391 279743 629
rect 307953 459 307987 629
rect 311449 595 311483 697
rect 312645 595 312679 765
rect 311173 255 311207 493
rect 334817 323 334851 561
rect 338681 119 338715 561
rect 338773 51 338807 561
rect 358737 391 358771 561
rect 362325 527 362359 629
rect 364717 459 364751 765
rect 370421 663 370455 901
rect 375205 663 375239 833
rect 364901 119 364935 561
rect 377505 527 377539 901
rect 388821 663 388855 1037
rect 393329 459 393363 833
rect 400045 663 400079 1105
rect 400229 595 400263 1037
rect 394191 561 394341 595
rect 404737 595 404771 765
rect 404829 595 404863 901
rect 394065 119 394099 493
rect 397745 187 397779 561
rect 399861 51 399895 425
rect 402161 119 402195 425
rect 403817 323 403851 425
rect 404921 391 404955 1105
rect 409245 663 409279 901
rect 412649 595 412683 833
rect 413753 595 413787 1309
rect 415501 595 415535 969
rect 418353 663 418387 969
rect 421021 663 421055 901
rect 425529 663 425563 1309
rect 425713 663 425747 969
rect 428381 595 428415 697
rect 431877 663 431911 1037
rect 435925 731 435959 969
rect 436477 663 436511 969
rect 414305 119 414339 561
rect 420929 187 420963 561
rect 423873 51 423907 561
rect 432061 119 432095 629
rect 434177 255 434211 629
rect 438685 595 438719 901
rect 439881 663 439915 1105
rect 440525 527 440559 765
rect 444481 595 444515 901
rect 445033 595 445067 1037
rect 446689 595 446723 765
rect 442641 255 442675 561
rect 449909 459 449943 629
rect 451657 459 451691 561
rect 451933 391 451967 561
rect 452301 391 452335 833
rect 453497 119 453531 1105
rect 453589 663 453623 1173
rect 454233 663 454267 969
rect 454509 51 454543 629
rect 454785 255 454819 629
rect 456073 595 456107 765
rect 458097 595 458131 901
rect 461501 595 461535 1105
rect 462145 663 462179 1241
rect 465641 459 465675 969
rect 466377 663 466411 1173
rect 467205 663 467239 1037
rect 468309 663 468343 1173
rect 470609 595 470643 901
rect 471713 595 471747 765
rect 474565 595 474599 969
rect 475761 595 475795 1105
rect 476957 595 476991 1241
rect 481741 595 481775 1037
rect 483029 663 483063 1173
rect 472265 323 472299 561
rect 484041 459 484075 629
rect 485145 187 485179 697
rect 485237 595 485271 901
rect 485329 663 485363 901
rect 486617 663 486651 833
rect 487445 663 487479 1309
rect 488273 663 488307 969
rect 487629 391 487663 629
rect 490941 595 490975 1037
rect 496829 663 496863 901
rect 498945 663 498979 901
rect 502349 663 502383 1241
rect 502993 663 503027 1309
rect 491125 51 491159 561
rect 503821 391 503855 561
rect 504005 391 504039 969
rect 504189 459 504223 697
rect 504649 459 504683 1309
rect 505753 663 505787 969
rect 506213 459 506247 1037
rect 507869 663 507903 1105
rect 509893 663 509927 833
rect 510261 187 510295 765
rect 510905 459 510939 697
rect 514401 663 514435 1173
rect 511181 323 511215 493
rect 513665 255 513699 561
rect 514493 119 514527 629
rect 514953 459 514987 901
rect 516977 663 517011 1037
rect 518173 935 518207 1241
rect 518265 663 518299 1241
rect 518357 663 518391 901
rect 520749 663 520783 1309
rect 521669 459 521703 697
rect 521761 51 521795 833
rect 521945 663 521979 969
rect 523049 595 523083 765
rect 523359 697 523727 731
rect 523693 527 523727 697
rect 524245 595 524279 1105
rect 531145 663 531179 1037
rect 525015 629 525165 663
rect 531329 663 531363 1173
rect 534549 119 534583 1241
rect 538229 595 538263 697
rect 538781 595 538815 833
rect 539793 527 539827 969
rect 540805 595 540839 901
rect 542001 595 542035 765
rect 538505 119 538539 493
rect 542369 323 542403 765
rect 542461 323 542495 833
rect 543381 595 543415 697
rect 544209 595 544243 1105
rect 545129 595 545163 1173
rect 544393 391 544427 561
rect 545497 51 545531 561
rect 549269 527 549303 697
rect 551109 663 551143 901
rect 551569 527 551603 765
rect 552489 391 552523 629
rect 554605 527 554639 1037
rect 558009 323 558043 969
rect 562057 595 562091 1105
rect 563253 595 563287 1173
<< viali >>
rect 50905 699397 50939 699431
rect 65625 699397 65659 699431
rect 80161 699397 80195 699431
rect 95157 699397 95191 699431
rect 109877 699397 109911 699431
rect 114569 699397 114603 699431
rect 124597 699397 124631 699431
rect 139317 699397 139351 699431
rect 139317 698785 139351 698819
rect 144285 699397 144319 699431
rect 168849 699397 168883 699431
rect 168849 698921 168883 698955
rect 173725 699397 173759 699431
rect 211261 699397 211295 699431
rect 211261 699193 211295 699227
rect 394157 699329 394191 699363
rect 394157 698989 394191 699023
rect 462881 699329 462915 699363
rect 173725 698853 173759 698887
rect 144285 698717 144319 698751
rect 124597 698649 124631 698683
rect 114569 698581 114603 698615
rect 109877 698513 109911 698547
rect 95157 698445 95191 698479
rect 80161 698377 80195 698411
rect 65625 698309 65659 698343
rect 462881 697765 462915 697799
rect 492597 699329 492631 699363
rect 492597 697697 492631 697731
rect 521853 699329 521887 699363
rect 521853 697629 521887 697663
rect 50905 697561 50939 697595
rect 413753 1309 413787 1343
rect 400045 1105 400079 1139
rect 388821 1037 388855 1071
rect 370421 901 370455 935
rect 312645 765 312679 799
rect 7481 697 7515 731
rect 240517 697 240551 731
rect 311449 697 311483 731
rect 240517 561 240551 595
rect 255513 629 255547 663
rect 7481 493 7515 527
rect 279709 629 279743 663
rect 298385 629 298419 663
rect 298569 629 298603 663
rect 307953 629 307987 663
rect 279617 561 279651 595
rect 279617 425 279651 459
rect 311449 561 311483 595
rect 364717 765 364751 799
rect 362325 629 362359 663
rect 312645 561 312679 595
rect 334817 561 334851 595
rect 307953 425 307987 459
rect 311173 493 311207 527
rect 279709 357 279743 391
rect 255513 289 255547 323
rect 334817 289 334851 323
rect 338681 561 338715 595
rect 311173 221 311207 255
rect 338681 85 338715 119
rect 338773 561 338807 595
rect 358737 561 358771 595
rect 362325 493 362359 527
rect 377505 901 377539 935
rect 370421 629 370455 663
rect 375205 833 375239 867
rect 375205 629 375239 663
rect 364717 425 364751 459
rect 364901 561 364935 595
rect 358737 357 358771 391
rect 388821 629 388855 663
rect 393329 833 393363 867
rect 377505 493 377539 527
rect 404921 1105 404955 1139
rect 400045 629 400079 663
rect 400229 1037 400263 1071
rect 404829 901 404863 935
rect 394157 561 394191 595
rect 394341 561 394375 595
rect 397745 561 397779 595
rect 400229 561 400263 595
rect 404737 765 404771 799
rect 404737 561 404771 595
rect 404829 561 404863 595
rect 393329 425 393363 459
rect 394065 493 394099 527
rect 364901 85 364935 119
rect 397745 153 397779 187
rect 399861 425 399895 459
rect 394065 85 394099 119
rect 338773 17 338807 51
rect 402161 425 402195 459
rect 403817 425 403851 459
rect 409245 901 409279 935
rect 409245 629 409279 663
rect 412649 833 412683 867
rect 412649 561 412683 595
rect 425529 1309 425563 1343
rect 415501 969 415535 1003
rect 418353 969 418387 1003
rect 418353 629 418387 663
rect 421021 901 421055 935
rect 421021 629 421055 663
rect 487445 1309 487479 1343
rect 462145 1241 462179 1275
rect 453589 1173 453623 1207
rect 439881 1105 439915 1139
rect 431877 1037 431911 1071
rect 425529 629 425563 663
rect 425713 969 425747 1003
rect 425713 629 425747 663
rect 428381 697 428415 731
rect 435925 969 435959 1003
rect 435925 697 435959 731
rect 436477 969 436511 1003
rect 431877 629 431911 663
rect 432061 629 432095 663
rect 413753 561 413787 595
rect 414305 561 414339 595
rect 415501 561 415535 595
rect 420929 561 420963 595
rect 404921 357 404955 391
rect 403817 289 403851 323
rect 402161 85 402195 119
rect 420929 153 420963 187
rect 423873 561 423907 595
rect 428381 561 428415 595
rect 414305 85 414339 119
rect 399861 17 399895 51
rect 434177 629 434211 663
rect 436477 629 436511 663
rect 438685 901 438719 935
rect 453497 1105 453531 1139
rect 445033 1037 445067 1071
rect 444481 901 444515 935
rect 439881 629 439915 663
rect 440525 765 440559 799
rect 438685 561 438719 595
rect 440525 493 440559 527
rect 442641 561 442675 595
rect 444481 561 444515 595
rect 452301 833 452335 867
rect 445033 561 445067 595
rect 446689 765 446723 799
rect 446689 561 446723 595
rect 449909 629 449943 663
rect 434177 221 434211 255
rect 449909 425 449943 459
rect 451657 561 451691 595
rect 451657 425 451691 459
rect 451933 561 451967 595
rect 451933 357 451967 391
rect 452301 357 452335 391
rect 442641 221 442675 255
rect 432061 85 432095 119
rect 461501 1105 461535 1139
rect 453589 629 453623 663
rect 454233 969 454267 1003
rect 458097 901 458131 935
rect 456073 765 456107 799
rect 454233 629 454267 663
rect 454509 629 454543 663
rect 453497 85 453531 119
rect 423873 17 423907 51
rect 454785 629 454819 663
rect 456073 561 456107 595
rect 458097 561 458131 595
rect 476957 1241 476991 1275
rect 466377 1173 466411 1207
rect 462145 629 462179 663
rect 465641 969 465675 1003
rect 461501 561 461535 595
rect 468309 1173 468343 1207
rect 466377 629 466411 663
rect 467205 1037 467239 1071
rect 467205 629 467239 663
rect 475761 1105 475795 1139
rect 474565 969 474599 1003
rect 468309 629 468343 663
rect 470609 901 470643 935
rect 470609 561 470643 595
rect 471713 765 471747 799
rect 471713 561 471747 595
rect 472265 561 472299 595
rect 474565 561 474599 595
rect 475761 561 475795 595
rect 483029 1173 483063 1207
rect 476957 561 476991 595
rect 481741 1037 481775 1071
rect 485237 901 485271 935
rect 485145 697 485179 731
rect 483029 629 483063 663
rect 484041 629 484075 663
rect 481741 561 481775 595
rect 465641 425 465675 459
rect 484041 425 484075 459
rect 472265 289 472299 323
rect 454785 221 454819 255
rect 485329 901 485363 935
rect 485329 629 485363 663
rect 486617 833 486651 867
rect 486617 629 486651 663
rect 502993 1309 503027 1343
rect 502349 1241 502383 1275
rect 490941 1037 490975 1071
rect 488273 969 488307 1003
rect 487445 629 487479 663
rect 487629 629 487663 663
rect 488273 629 488307 663
rect 485237 561 485271 595
rect 496829 901 496863 935
rect 496829 629 496863 663
rect 498945 901 498979 935
rect 498945 629 498979 663
rect 502349 629 502383 663
rect 504649 1309 504683 1343
rect 502993 629 503027 663
rect 504005 969 504039 1003
rect 490941 561 490975 595
rect 491125 561 491159 595
rect 487629 357 487663 391
rect 485145 153 485179 187
rect 454509 17 454543 51
rect 503821 561 503855 595
rect 503821 357 503855 391
rect 504189 697 504223 731
rect 504189 425 504223 459
rect 520749 1309 520783 1343
rect 518173 1241 518207 1275
rect 514401 1173 514435 1207
rect 507869 1105 507903 1139
rect 506213 1037 506247 1071
rect 505753 969 505787 1003
rect 505753 629 505787 663
rect 504649 425 504683 459
rect 507869 629 507903 663
rect 509893 833 509927 867
rect 509893 629 509927 663
rect 510261 765 510295 799
rect 506213 425 506247 459
rect 504005 357 504039 391
rect 510905 697 510939 731
rect 516977 1037 517011 1071
rect 514953 901 514987 935
rect 514401 629 514435 663
rect 514493 629 514527 663
rect 513665 561 513699 595
rect 510905 425 510939 459
rect 511181 493 511215 527
rect 511181 289 511215 323
rect 513665 221 513699 255
rect 510261 153 510295 187
rect 518173 901 518207 935
rect 518265 1241 518299 1275
rect 516977 629 517011 663
rect 518265 629 518299 663
rect 518357 901 518391 935
rect 518357 629 518391 663
rect 534549 1241 534583 1275
rect 531329 1173 531363 1207
rect 524245 1105 524279 1139
rect 521945 969 521979 1003
rect 521761 833 521795 867
rect 520749 629 520783 663
rect 521669 697 521703 731
rect 514953 425 514987 459
rect 521669 425 521703 459
rect 514493 85 514527 119
rect 491125 17 491159 51
rect 521945 629 521979 663
rect 523049 765 523083 799
rect 523325 697 523359 731
rect 523049 561 523083 595
rect 531145 1037 531179 1071
rect 524981 629 525015 663
rect 525165 629 525199 663
rect 531145 629 531179 663
rect 531329 629 531363 663
rect 524245 561 524279 595
rect 523693 493 523727 527
rect 545129 1173 545163 1207
rect 544209 1105 544243 1139
rect 539793 969 539827 1003
rect 538781 833 538815 867
rect 538229 697 538263 731
rect 538229 561 538263 595
rect 538781 561 538815 595
rect 540805 901 540839 935
rect 542461 833 542495 867
rect 540805 561 540839 595
rect 542001 765 542035 799
rect 542001 561 542035 595
rect 542369 765 542403 799
rect 534549 85 534583 119
rect 538505 493 538539 527
rect 539793 493 539827 527
rect 542369 289 542403 323
rect 543381 697 543415 731
rect 543381 561 543415 595
rect 563253 1173 563287 1207
rect 562057 1105 562091 1139
rect 554605 1037 554639 1071
rect 551109 901 551143 935
rect 549269 697 549303 731
rect 544209 561 544243 595
rect 544393 561 544427 595
rect 545129 561 545163 595
rect 545497 561 545531 595
rect 544393 357 544427 391
rect 542461 289 542495 323
rect 538505 85 538539 119
rect 521761 17 521795 51
rect 551109 629 551143 663
rect 551569 765 551603 799
rect 549269 493 549303 527
rect 551569 493 551603 527
rect 552489 629 552523 663
rect 554605 493 554639 527
rect 558009 969 558043 1003
rect 552489 357 552523 391
rect 562057 561 562091 595
rect 563253 561 563287 595
rect 558009 289 558043 323
rect 545497 17 545531 51
<< metal1 >>
rect 271782 703808 271788 703860
rect 271840 703848 271846 703860
rect 364702 703848 364708 703860
rect 271840 703820 364708 703848
rect 271840 703808 271846 703820
rect 364702 703808 364708 703820
rect 364760 703808 364766 703860
rect 257246 703740 257252 703792
rect 257304 703780 257310 703792
rect 371602 703780 371608 703792
rect 257304 703752 371608 703780
rect 257304 703740 257310 703752
rect 371602 703740 371608 703752
rect 371660 703740 371666 703792
rect 276842 703672 276848 703724
rect 276900 703712 276906 703724
rect 332318 703712 332324 703724
rect 276900 703684 332324 703712
rect 276900 703672 276906 703684
rect 332318 703672 332324 703684
rect 332376 703672 332382 703724
rect 300854 703644 300860 703656
rect 238726 703616 300860 703644
rect 235350 703536 235356 703588
rect 235408 703576 235414 703588
rect 238726 703576 238754 703616
rect 300854 703604 300860 703616
rect 300912 703604 300918 703656
rect 235408 703548 238754 703576
rect 235408 703536 235414 703548
rect 242434 703536 242440 703588
rect 242492 703576 242498 703588
rect 400858 703576 400864 703588
rect 242492 703548 400864 703576
rect 242492 703536 242498 703548
rect 400858 703536 400864 703548
rect 400916 703536 400922 703588
rect 315482 703508 315488 703520
rect 171106 703480 315488 703508
rect 170306 703400 170312 703452
rect 170364 703440 170370 703452
rect 171106 703440 171134 703480
rect 315482 703468 315488 703480
rect 315540 703468 315546 703520
rect 170364 703412 171134 703440
rect 170364 703400 170370 703412
rect 227622 703400 227628 703452
rect 227680 703440 227686 703452
rect 497458 703440 497464 703452
rect 227680 703412 497464 703440
rect 227680 703400 227686 703412
rect 497458 703400 497464 703412
rect 497516 703400 497522 703452
rect 1486 703332 1492 703384
rect 1544 703372 1550 703384
rect 359734 703372 359740 703384
rect 1544 703344 359740 703372
rect 1544 703332 1550 703344
rect 359734 703332 359740 703344
rect 359792 703332 359798 703384
rect 212994 703264 213000 703316
rect 213052 703304 213058 703316
rect 576394 703304 576400 703316
rect 213052 703276 576400 703304
rect 213052 703264 213058 703276
rect 576394 703264 576400 703276
rect 576452 703264 576458 703316
rect 1578 703196 1584 703248
rect 1636 703236 1642 703248
rect 374454 703236 374460 703248
rect 1636 703208 374460 703236
rect 1636 703196 1642 703208
rect 374454 703196 374460 703208
rect 374512 703196 374518 703248
rect 198274 703128 198280 703180
rect 198332 703168 198338 703180
rect 575106 703168 575112 703180
rect 198332 703140 575112 703168
rect 198332 703128 198338 703140
rect 575106 703128 575112 703140
rect 575164 703128 575170 703180
rect 1670 703060 1676 703112
rect 1728 703100 1734 703112
rect 389174 703100 389180 703112
rect 1728 703072 389180 703100
rect 1728 703060 1734 703072
rect 389174 703060 389180 703072
rect 389232 703060 389238 703112
rect 183370 702992 183376 703044
rect 183428 703032 183434 703044
rect 573726 703032 573732 703044
rect 183428 703004 573732 703032
rect 183428 702992 183434 703004
rect 573726 702992 573732 703004
rect 573784 702992 573790 703044
rect 1854 702924 1860 702976
rect 1912 702964 1918 702976
rect 403894 702964 403900 702976
rect 1912 702936 403900 702964
rect 1912 702924 1918 702936
rect 403894 702924 403900 702936
rect 403952 702924 403958 702976
rect 158622 702856 158628 702908
rect 158680 702896 158686 702908
rect 575014 702896 575020 702908
rect 158680 702868 575020 702896
rect 158680 702856 158686 702868
rect 575014 702856 575020 702868
rect 575072 702856 575078 702908
rect 750 702788 756 702840
rect 808 702828 814 702840
rect 423674 702828 423680 702840
rect 808 702800 423680 702828
rect 808 702788 814 702800
rect 423674 702788 423680 702800
rect 423732 702788 423738 702840
rect 2314 702720 2320 702772
rect 2372 702760 2378 702772
rect 477586 702760 477592 702772
rect 2372 702732 477592 702760
rect 2372 702720 2378 702732
rect 477586 702720 477592 702732
rect 477644 702720 477650 702772
rect 382 702652 388 702704
rect 440 702692 446 702704
rect 497274 702692 497280 702704
rect 440 702664 497280 702692
rect 440 702652 446 702664
rect 497274 702652 497280 702664
rect 497332 702652 497338 702704
rect 290 702584 296 702636
rect 348 702624 354 702636
rect 507118 702624 507124 702636
rect 348 702596 507124 702624
rect 348 702584 354 702596
rect 507118 702584 507124 702596
rect 507176 702584 507182 702636
rect 106 702516 112 702568
rect 164 702556 170 702568
rect 536834 702556 536840 702568
rect 164 702528 536840 702556
rect 164 702516 170 702528
rect 536834 702516 536840 702528
rect 536892 702516 536898 702568
rect 35802 702448 35808 702500
rect 35860 702488 35866 702500
rect 574738 702488 574744 702500
rect 35860 702460 574744 702488
rect 35860 702448 35866 702460
rect 574738 702448 574744 702460
rect 574796 702448 574802 702500
rect 154022 702380 154028 702432
rect 154080 702420 154086 702432
rect 311158 702420 311164 702432
rect 154080 702392 311164 702420
rect 154080 702380 154086 702392
rect 311158 702380 311164 702392
rect 311216 702380 311222 702432
rect 75454 702312 75460 702364
rect 75512 702352 75518 702364
rect 573450 702352 573456 702364
rect 75512 702324 573456 702352
rect 75512 702312 75518 702324
rect 573450 702312 573456 702324
rect 573508 702312 573514 702364
rect 237098 702244 237104 702296
rect 237156 702284 237162 702296
rect 305822 702284 305828 702296
rect 237156 702256 305828 702284
rect 237156 702244 237162 702256
rect 305822 702244 305828 702256
rect 305880 702244 305886 702296
rect 311066 702176 311072 702228
rect 311124 702216 311130 702228
rect 364610 702216 364616 702228
rect 311124 702188 364616 702216
rect 311124 702176 311130 702188
rect 364610 702176 364616 702188
rect 364668 702176 364674 702228
rect 178586 702108 178592 702160
rect 178644 702148 178650 702160
rect 339310 702148 339316 702160
rect 178644 702120 339316 702148
rect 178644 702108 178650 702120
rect 339310 702108 339316 702120
rect 339368 702108 339374 702160
rect 163866 702040 163872 702092
rect 163924 702080 163930 702092
rect 331306 702080 331312 702092
rect 163924 702052 331312 702080
rect 163924 702040 163930 702052
rect 331306 702040 331312 702052
rect 331364 702040 331370 702092
rect 335906 702040 335912 702092
rect 335964 702080 335970 702092
rect 467834 702080 467840 702092
rect 335964 702052 467840 702080
rect 335964 702040 335970 702052
rect 467834 702040 467840 702052
rect 467892 702040 467898 702092
rect 188430 701972 188436 702024
rect 188488 702012 188494 702024
rect 243354 702012 243360 702024
rect 188488 701984 243360 702012
rect 188488 701972 188494 701984
rect 243354 701972 243360 701984
rect 243412 701972 243418 702024
rect 262122 701972 262128 702024
rect 262180 702012 262186 702024
rect 482554 702012 482560 702024
rect 262180 701984 482560 702012
rect 262180 701972 262186 701984
rect 482554 701972 482560 701984
rect 482612 701972 482618 702024
rect 266354 701904 266360 701956
rect 266412 701944 266418 701956
rect 502334 701944 502340 701956
rect 266412 701916 502340 701944
rect 266412 701904 266418 701916
rect 502334 701904 502340 701916
rect 502392 701904 502398 701956
rect 70118 701836 70124 701888
rect 70176 701876 70182 701888
rect 329374 701876 329380 701888
rect 70176 701848 329380 701876
rect 70176 701836 70182 701848
rect 329374 701836 329380 701848
rect 329432 701836 329438 701888
rect 350534 701836 350540 701888
rect 350592 701876 350598 701888
rect 511994 701876 512000 701888
rect 350592 701848 512000 701876
rect 350592 701836 350598 701848
rect 511994 701836 512000 701848
rect 512052 701836 512058 701888
rect 1302 701768 1308 701820
rect 1360 701808 1366 701820
rect 414198 701808 414204 701820
rect 1360 701780 414204 701808
rect 1360 701768 1366 701780
rect 414198 701768 414204 701780
rect 414256 701768 414262 701820
rect 148962 701700 148968 701752
rect 149020 701740 149026 701752
rect 577498 701740 577504 701752
rect 149020 701712 577504 701740
rect 149020 701700 149026 701712
rect 577498 701700 577504 701712
rect 577556 701700 577562 701752
rect 4338 701632 4344 701684
rect 4396 701672 4402 701684
rect 443270 701672 443276 701684
rect 4396 701644 443276 701672
rect 4396 701632 4402 701644
rect 443270 701632 443276 701644
rect 443328 701632 443334 701684
rect 444282 701632 444288 701684
rect 444340 701672 444346 701684
rect 541526 701672 541532 701684
rect 444340 701644 541532 701672
rect 444340 701632 444346 701644
rect 541526 701632 541532 701644
rect 541584 701632 541590 701684
rect 129458 701564 129464 701616
rect 129516 701604 129522 701616
rect 574922 701604 574928 701616
rect 129516 701576 574928 701604
rect 129516 701564 129522 701576
rect 574922 701564 574928 701576
rect 574980 701564 574986 701616
rect 2590 701496 2596 701548
rect 2648 701536 2654 701548
rect 458174 701536 458180 701548
rect 2648 701508 458180 701536
rect 2648 701496 2654 701508
rect 458174 701496 458180 701508
rect 458232 701496 458238 701548
rect 119706 701428 119712 701480
rect 119764 701468 119770 701480
rect 576302 701468 576308 701480
rect 119764 701440 576308 701468
rect 119764 701428 119770 701440
rect 576302 701428 576308 701440
rect 576360 701428 576366 701480
rect 104802 701360 104808 701412
rect 104860 701400 104866 701412
rect 574830 701400 574836 701412
rect 104860 701372 574836 701400
rect 104860 701360 104866 701372
rect 574830 701360 574836 701372
rect 574888 701360 574894 701412
rect 100018 701292 100024 701344
rect 100076 701332 100082 701344
rect 576210 701332 576216 701344
rect 100076 701304 576216 701332
rect 100076 701292 100082 701304
rect 576210 701292 576216 701304
rect 576268 701292 576274 701344
rect 90174 701224 90180 701276
rect 90232 701264 90238 701276
rect 573542 701264 573548 701276
rect 90232 701236 573548 701264
rect 90232 701224 90238 701236
rect 573542 701224 573548 701236
rect 573600 701224 573606 701276
rect 85298 701156 85304 701208
rect 85356 701196 85362 701208
rect 569310 701196 569316 701208
rect 85356 701168 569316 701196
rect 85356 701156 85362 701168
rect 569310 701156 569316 701168
rect 569368 701156 569374 701208
rect 566 701088 572 701140
rect 624 701128 630 701140
rect 487430 701128 487436 701140
rect 624 701100 487436 701128
rect 624 701088 630 701100
rect 487430 701088 487436 701100
rect 487488 701088 487494 701140
rect 55766 701020 55772 701072
rect 55824 701060 55830 701072
rect 271506 701060 271512 701072
rect 55824 701032 271512 701060
rect 55824 701020 55830 701032
rect 271506 701020 271512 701032
rect 271564 701020 271570 701072
rect 282914 701020 282920 701072
rect 282972 701060 282978 701072
rect 291194 701060 291200 701072
rect 282972 701032 291200 701060
rect 282972 701020 282978 701032
rect 291194 701020 291200 701032
rect 291252 701020 291258 701072
rect 291378 701020 291384 701072
rect 291436 701060 291442 701072
rect 295886 701060 295892 701072
rect 291436 701032 295892 701060
rect 291436 701020 291442 701032
rect 295886 701020 295892 701032
rect 295944 701020 295950 701072
rect 331214 701020 331220 701072
rect 331272 701060 331278 701072
rect 335354 701060 335360 701072
rect 331272 701032 335360 701060
rect 331272 701020 331278 701032
rect 335354 701020 335360 701032
rect 335412 701020 335418 701072
rect 339402 701020 339408 701072
rect 339460 701060 339466 701072
rect 344922 701060 344928 701072
rect 339460 701032 344928 701060
rect 339460 701020 339466 701032
rect 344922 701020 344928 701032
rect 344980 701020 344986 701072
rect 349890 701060 349896 701072
rect 346320 701032 349896 701060
rect 8110 700952 8116 701004
rect 8168 700992 8174 701004
rect 346320 700992 346348 701032
rect 349890 701020 349896 701032
rect 349948 701020 349954 701072
rect 8168 700964 346348 700992
rect 8168 700952 8174 700964
rect 400858 700952 400864 701004
rect 400916 700992 400922 701004
rect 494790 700992 494796 701004
rect 400916 700964 494796 700992
rect 400916 700952 400922 700964
rect 494790 700952 494796 700964
rect 494848 700952 494854 701004
rect 497458 700952 497464 701004
rect 497516 700992 497522 701004
rect 559650 700992 559656 701004
rect 497516 700964 559656 700992
rect 497516 700952 497522 700964
rect 559650 700952 559656 700964
rect 559708 700952 559714 701004
rect 40494 700884 40500 700936
rect 40552 700924 40558 700936
rect 339402 700924 339408 700936
rect 40552 700896 339408 700924
rect 40552 700884 40558 700896
rect 339402 700884 339408 700896
rect 339460 700884 339466 700936
rect 371602 700884 371608 700936
rect 371660 700924 371666 700936
rect 429838 700924 429844 700936
rect 371660 700896 429844 700924
rect 371660 700884 371666 700896
rect 429838 700884 429844 700896
rect 429896 700884 429902 700936
rect 72970 700816 72976 700868
rect 73028 700856 73034 700868
rect 331214 700856 331220 700868
rect 73028 700828 331220 700856
rect 73028 700816 73034 700828
rect 331214 700816 331220 700828
rect 331272 700816 331278 700868
rect 202782 700748 202788 700800
rect 202840 700788 202846 700800
rect 305730 700788 305736 700800
rect 202840 700760 305736 700788
rect 202840 700748 202846 700760
rect 305730 700748 305736 700760
rect 305788 700748 305794 700800
rect 305822 700748 305828 700800
rect 305880 700788 305886 700800
rect 543458 700788 543464 700800
rect 305880 700760 543464 700788
rect 305880 700748 305886 700760
rect 543458 700748 543464 700760
rect 543516 700748 543522 700800
rect 137830 700680 137836 700732
rect 137888 700720 137894 700732
rect 320450 700720 320456 700732
rect 137888 700692 320456 700720
rect 137888 700680 137894 700692
rect 320450 700680 320456 700692
rect 320508 700680 320514 700732
rect 339310 700680 339316 700732
rect 339368 700720 339374 700732
rect 580718 700720 580724 700732
rect 339368 700692 580724 700720
rect 339368 700680 339374 700692
rect 580718 700680 580724 700692
rect 580776 700680 580782 700732
rect 105446 700612 105452 700664
rect 105504 700652 105510 700664
rect 330294 700652 330300 700664
rect 105504 700624 330300 700652
rect 105504 700612 105510 700624
rect 330294 700612 330300 700624
rect 330352 700612 330358 700664
rect 331306 700612 331312 700664
rect 331364 700652 331370 700664
rect 580626 700652 580632 700664
rect 331364 700624 580632 700652
rect 331364 700612 331370 700624
rect 580626 700612 580632 700624
rect 580684 700612 580690 700664
rect 89162 700544 89168 700596
rect 89220 700584 89226 700596
rect 340046 700584 340052 700596
rect 89220 700556 340052 700584
rect 89220 700544 89226 700556
rect 340046 700544 340052 700556
rect 340104 700544 340110 700596
rect 3878 700476 3884 700528
rect 3936 700516 3942 700528
rect 262122 700516 262128 700528
rect 3936 700488 262128 700516
rect 3936 700476 3942 700488
rect 262122 700476 262128 700488
rect 262180 700476 262186 700528
rect 281350 700476 281356 700528
rect 281408 700516 281414 700528
rect 348786 700516 348792 700528
rect 281408 700488 348792 700516
rect 281408 700476 281414 700488
rect 348786 700476 348792 700488
rect 348844 700476 348850 700528
rect 3694 700408 3700 700460
rect 3752 700448 3758 700460
rect 266354 700448 266360 700460
rect 3752 700420 266360 700448
rect 3752 700408 3758 700420
rect 266354 700408 266360 700420
rect 266412 700408 266418 700460
rect 267642 700408 267648 700460
rect 267700 700448 267706 700460
rect 282914 700448 282920 700460
rect 267700 700420 282920 700448
rect 267700 700408 267706 700420
rect 282914 700408 282920 700420
rect 282972 700408 282978 700460
rect 284110 700408 284116 700460
rect 284168 700448 284174 700460
rect 291378 700448 291384 700460
rect 284168 700420 291384 700448
rect 284168 700408 284174 700420
rect 291378 700408 291384 700420
rect 291436 700408 291442 700460
rect 291470 700408 291476 700460
rect 291528 700448 291534 700460
rect 300118 700448 300124 700460
rect 291528 700420 300124 700448
rect 291528 700408 291534 700420
rect 300118 700408 300124 700420
rect 300176 700408 300182 700460
rect 311158 700408 311164 700460
rect 311216 700448 311222 700460
rect 580534 700448 580540 700460
rect 311216 700420 580540 700448
rect 311216 700408 311222 700420
rect 580534 700408 580540 700420
rect 580592 700408 580598 700460
rect 232682 700340 232688 700392
rect 232740 700380 232746 700392
rect 527174 700380 527180 700392
rect 232740 700352 527180 700380
rect 232740 700340 232746 700352
rect 527174 700340 527180 700352
rect 527232 700340 527238 700392
rect 24302 700272 24308 700324
rect 24360 700312 24366 700324
rect 354950 700312 354956 700324
rect 24360 700284 354956 700312
rect 24360 700272 24366 700284
rect 354950 700272 354956 700284
rect 355008 700272 355014 700324
rect 252278 700204 252284 700256
rect 252336 700244 252342 700256
rect 478506 700244 478512 700256
rect 252336 700216 478512 700244
rect 252336 700204 252342 700216
rect 478506 700204 478512 700216
rect 478564 700204 478570 700256
rect 247080 700136 247086 700188
rect 247138 700176 247144 700188
rect 462314 700176 462320 700188
rect 247138 700148 462320 700176
rect 247138 700136 247144 700148
rect 462314 700136 462320 700148
rect 462372 700136 462378 700188
rect 154114 700068 154120 700120
rect 154172 700108 154178 700120
rect 325648 700108 325654 700120
rect 154172 700080 325654 700108
rect 154172 700068 154178 700080
rect 325648 700068 325654 700080
rect 325706 700068 325712 700120
rect 329374 700068 329380 700120
rect 329432 700108 329438 700120
rect 580350 700108 580356 700120
rect 329432 700080 580356 700108
rect 329432 700068 329438 700080
rect 580350 700068 580356 700080
rect 580408 700068 580414 700120
rect 266998 700000 267004 700052
rect 267056 700040 267062 700052
rect 413646 700040 413652 700052
rect 267056 700012 413652 700040
rect 267056 700000 267062 700012
rect 413646 700000 413652 700012
rect 413704 700000 413710 700052
rect 262122 699932 262128 699984
rect 262180 699972 262186 699984
rect 397454 699972 397460 699984
rect 262180 699944 397460 699972
rect 262180 699932 262186 699944
rect 397454 699932 397460 699944
rect 397512 699932 397518 699984
rect 218974 699864 218980 699916
rect 219032 699904 219038 699916
rect 310606 699904 310612 699916
rect 219032 699876 310612 699904
rect 219032 699864 219038 699876
rect 310606 699864 310612 699876
rect 310664 699864 310670 699916
rect 217870 699796 217876 699848
rect 217928 699836 217934 699848
rect 563514 699836 563520 699848
rect 217928 699808 563520 699836
rect 217928 699796 217934 699808
rect 563514 699796 563520 699808
rect 563572 699796 563578 699848
rect 3234 699728 3240 699780
rect 3292 699768 3298 699780
rect 369762 699768 369768 699780
rect 3292 699740 369768 699768
rect 3292 699728 3298 699740
rect 369762 699728 369768 699740
rect 369820 699728 369826 699780
rect 3786 699660 3792 699712
rect 3844 699700 3850 699712
rect 384298 699700 384304 699712
rect 3844 699672 384304 699700
rect 3844 699660 3850 699672
rect 384298 699660 384304 699672
rect 384356 699660 384362 699712
rect 3050 699592 3056 699644
rect 3108 699632 3114 699644
rect 311066 699632 311072 699644
rect 3108 699604 311072 699632
rect 3108 699592 3114 699604
rect 311066 699592 311072 699604
rect 311124 699592 311130 699644
rect 271506 699524 271512 699576
rect 271564 699564 271570 699576
rect 580258 699564 580264 699576
rect 271564 699536 580264 699564
rect 271564 699524 271570 699536
rect 580258 699524 580264 699536
rect 580316 699524 580322 699576
rect 3970 699456 3976 699508
rect 4028 699496 4034 699508
rect 335906 699496 335912 699508
rect 4028 699468 335912 699496
rect 4028 699456 4034 699468
rect 335906 699456 335912 699468
rect 335964 699456 335970 699508
rect 50890 699428 50896 699440
rect 50851 699400 50896 699428
rect 50890 699388 50896 699400
rect 50948 699388 50954 699440
rect 65610 699428 65616 699440
rect 65571 699400 65616 699428
rect 65610 699388 65616 699400
rect 65668 699388 65674 699440
rect 80146 699428 80152 699440
rect 80107 699400 80152 699428
rect 80146 699388 80152 699400
rect 80204 699388 80210 699440
rect 95142 699428 95148 699440
rect 95103 699400 95148 699428
rect 95142 699388 95148 699400
rect 95200 699388 95206 699440
rect 109862 699428 109868 699440
rect 109823 699400 109868 699428
rect 109862 699388 109868 699400
rect 109920 699388 109926 699440
rect 114554 699428 114560 699440
rect 114515 699400 114560 699428
rect 114554 699388 114560 699400
rect 114612 699388 114618 699440
rect 124582 699428 124588 699440
rect 124543 699400 124588 699428
rect 124582 699388 124588 699400
rect 124640 699388 124646 699440
rect 139302 699428 139308 699440
rect 139263 699400 139308 699428
rect 139302 699388 139308 699400
rect 139360 699388 139366 699440
rect 144270 699428 144276 699440
rect 144231 699400 144276 699428
rect 144270 699388 144276 699400
rect 144328 699388 144334 699440
rect 168834 699428 168840 699440
rect 168795 699400 168840 699428
rect 168834 699388 168840 699400
rect 168892 699388 168898 699440
rect 173710 699428 173716 699440
rect 173671 699400 173716 699428
rect 173710 699388 173716 699400
rect 173768 699388 173774 699440
rect 180766 699400 203104 699428
rect 3510 699320 3516 699372
rect 3568 699360 3574 699372
rect 180766 699360 180794 699400
rect 3568 699332 180794 699360
rect 3568 699320 3574 699332
rect 193214 699320 193220 699372
rect 193272 699360 193278 699372
rect 193272 699332 200114 699360
rect 193272 699320 193278 699332
rect 200086 699088 200114 699332
rect 202966 699320 202972 699372
rect 203024 699320 203030 699372
rect 203076 699360 203104 699400
rect 208118 699388 208124 699440
rect 208176 699428 208182 699440
rect 211249 699431 211307 699437
rect 211249 699428 211261 699431
rect 208176 699400 211261 699428
rect 208176 699388 208182 699400
rect 211249 699397 211261 699400
rect 211295 699397 211307 699431
rect 211249 699391 211307 699397
rect 219406 699400 229094 699428
rect 219406 699360 219434 699400
rect 203076 699332 219434 699360
rect 222838 699320 222844 699372
rect 222896 699320 222902 699372
rect 229066 699360 229094 699400
rect 243354 699388 243360 699440
rect 243412 699428 243418 699440
rect 580810 699428 580816 699440
rect 243412 699400 580816 699428
rect 243412 699388 243418 699400
rect 580810 699388 580816 699400
rect 580868 699388 580874 699440
rect 350534 699360 350540 699372
rect 229066 699332 350540 699360
rect 350534 699320 350540 699332
rect 350592 699320 350598 699372
rect 394142 699360 394148 699372
rect 394103 699332 394148 699360
rect 394142 699320 394148 699332
rect 394200 699320 394206 699372
rect 462866 699360 462872 699372
rect 462827 699332 462872 699360
rect 462866 699320 462872 699332
rect 462924 699320 462930 699372
rect 492582 699360 492588 699372
rect 492543 699332 492588 699360
rect 492582 699320 492588 699332
rect 492640 699320 492646 699372
rect 521838 699360 521844 699372
rect 521799 699332 521844 699360
rect 521838 699320 521844 699332
rect 521896 699320 521902 699372
rect 202984 699156 203012 699320
rect 222856 699292 222884 699320
rect 563698 699292 563704 699304
rect 222856 699264 563704 699292
rect 563698 699252 563704 699264
rect 563756 699252 563762 699304
rect 211249 699227 211307 699233
rect 211249 699193 211261 699227
rect 211295 699224 211307 699227
rect 567838 699224 567844 699236
rect 211295 699196 567844 699224
rect 211295 699193 211307 699196
rect 211249 699187 211307 699193
rect 567838 699184 567844 699196
rect 567896 699184 567902 699236
rect 578970 699156 578976 699168
rect 202984 699128 578976 699156
rect 578970 699116 578976 699128
rect 579028 699116 579034 699168
rect 572162 699088 572168 699100
rect 200086 699060 572168 699088
rect 572162 699048 572168 699060
rect 572220 699048 572226 699100
rect 842 698980 848 699032
rect 900 699020 906 699032
rect 394145 699023 394203 699029
rect 394145 699020 394157 699023
rect 900 698992 394157 699020
rect 900 698980 906 698992
rect 394145 698989 394157 698992
rect 394191 698989 394203 699023
rect 394145 698983 394203 698989
rect 168837 698955 168895 698961
rect 168837 698921 168849 698955
rect 168883 698952 168895 698955
rect 566826 698952 566832 698964
rect 168883 698924 566832 698952
rect 168883 698921 168895 698924
rect 168837 698915 168895 698921
rect 566826 698912 566832 698924
rect 566884 698912 566890 698964
rect 173713 698887 173771 698893
rect 173713 698853 173725 698887
rect 173759 698884 173771 698887
rect 573634 698884 573640 698896
rect 173759 698856 573640 698884
rect 173759 698853 173771 698856
rect 173713 698847 173771 698853
rect 573634 698844 573640 698856
rect 573692 698844 573698 698896
rect 139305 698819 139363 698825
rect 139305 698785 139317 698819
rect 139351 698816 139363 698819
rect 570690 698816 570696 698828
rect 139351 698788 570696 698816
rect 139351 698785 139363 698788
rect 139305 698779 139363 698785
rect 570690 698776 570696 698788
rect 570748 698776 570754 698828
rect 144273 698751 144331 698757
rect 144273 698717 144285 698751
rect 144319 698748 144331 698751
rect 578878 698748 578884 698760
rect 144319 698720 578884 698748
rect 144319 698717 144331 698720
rect 144273 698711 144331 698717
rect 578878 698708 578884 698720
rect 578936 698708 578942 698760
rect 124585 698683 124643 698689
rect 124585 698649 124597 698683
rect 124631 698680 124643 698683
rect 572070 698680 572076 698692
rect 124631 698652 572076 698680
rect 124631 698649 124643 698652
rect 124585 698643 124643 698649
rect 572070 698640 572076 698652
rect 572128 698640 572134 698692
rect 114557 698615 114615 698621
rect 114557 698581 114569 698615
rect 114603 698612 114615 698615
rect 570598 698612 570604 698624
rect 114603 698584 570604 698612
rect 114603 698581 114615 698584
rect 114557 698575 114615 698581
rect 570598 698572 570604 698584
rect 570656 698572 570662 698624
rect 109865 698547 109923 698553
rect 109865 698513 109877 698547
rect 109911 698544 109923 698547
rect 569494 698544 569500 698556
rect 109911 698516 569500 698544
rect 109911 698513 109923 698516
rect 109865 698507 109923 698513
rect 569494 698504 569500 698516
rect 569552 698504 569558 698556
rect 95145 698479 95203 698485
rect 95145 698445 95157 698479
rect 95191 698476 95203 698479
rect 565354 698476 565360 698488
rect 95191 698448 565360 698476
rect 95191 698445 95203 698448
rect 95145 698439 95203 698445
rect 565354 698436 565360 698448
rect 565412 698436 565418 698488
rect 80149 698411 80207 698417
rect 80149 698377 80161 698411
rect 80195 698408 80207 698411
rect 566734 698408 566740 698420
rect 80195 698380 566740 698408
rect 80195 698377 80207 698380
rect 80149 698371 80207 698377
rect 566734 698368 566740 698380
rect 566792 698368 566798 698420
rect 65613 698343 65671 698349
rect 65613 698309 65625 698343
rect 65659 698340 65671 698343
rect 566550 698340 566556 698352
rect 65659 698312 566556 698340
rect 65659 698309 65671 698312
rect 65613 698303 65671 698309
rect 566550 698300 566556 698312
rect 566608 698300 566614 698352
rect 563514 698232 563520 698284
rect 563572 698272 563578 698284
rect 580166 698272 580172 698284
rect 563572 698244 580172 698272
rect 563572 698232 563578 698244
rect 580166 698232 580172 698244
rect 580224 698232 580230 698284
rect 2406 697756 2412 697808
rect 2464 697796 2470 697808
rect 462869 697799 462927 697805
rect 462869 697796 462881 697799
rect 2464 697768 462881 697796
rect 2464 697756 2470 697768
rect 462869 697765 462881 697768
rect 462915 697765 462927 697799
rect 462869 697759 462927 697765
rect 474 697688 480 697740
rect 532 697728 538 697740
rect 492585 697731 492643 697737
rect 492585 697728 492597 697731
rect 532 697700 492597 697728
rect 532 697688 538 697700
rect 492585 697697 492597 697700
rect 492631 697697 492643 697731
rect 492585 697691 492643 697697
rect 198 697620 204 697672
rect 256 697660 262 697672
rect 521841 697663 521899 697669
rect 521841 697660 521853 697663
rect 256 697632 521853 697660
rect 256 697620 262 697632
rect 521841 697629 521853 697632
rect 521887 697629 521899 697663
rect 521841 697623 521899 697629
rect 50893 697595 50951 697601
rect 50893 697561 50905 697595
rect 50939 697592 50951 697595
rect 573358 697592 573364 697604
rect 50939 697564 573364 697592
rect 50939 697561 50951 697564
rect 50893 697555 50951 697561
rect 573358 697552 573364 697564
rect 573416 697552 573422 697604
rect 563698 684428 563704 684480
rect 563756 684468 563762 684480
rect 580166 684468 580172 684480
rect 563756 684440 580172 684468
rect 563756 684428 563762 684440
rect 580166 684428 580172 684440
rect 580224 684428 580230 684480
rect 576394 671984 576400 672036
rect 576452 672024 576458 672036
rect 580166 672024 580172 672036
rect 576452 671996 580172 672024
rect 576452 671984 576458 671996
rect 580166 671984 580172 671996
rect 580224 671984 580230 672036
rect 3234 661036 3240 661088
rect 3292 661076 3298 661088
rect 4338 661076 4344 661088
rect 3292 661048 4344 661076
rect 3292 661036 3298 661048
rect 4338 661036 4344 661048
rect 4396 661036 4402 661088
rect 567838 632000 567844 632052
rect 567896 632040 567902 632052
rect 580166 632040 580172 632052
rect 567896 632012 580172 632040
rect 567896 632000 567902 632012
rect 580166 632000 580172 632012
rect 580224 632000 580230 632052
rect 1302 619556 1308 619608
rect 1360 619596 1366 619608
rect 2774 619596 2780 619608
rect 1360 619568 2780 619596
rect 1360 619556 1366 619568
rect 2774 619556 2780 619568
rect 2832 619556 2838 619608
rect 575106 618196 575112 618248
rect 575164 618236 575170 618248
rect 580166 618236 580172 618248
rect 575164 618208 580172 618236
rect 575164 618196 575170 618208
rect 580166 618196 580172 618208
rect 580224 618196 580230 618248
rect 572162 578144 572168 578196
rect 572220 578184 572226 578196
rect 579798 578184 579804 578196
rect 572220 578156 579804 578184
rect 572220 578144 572226 578156
rect 579798 578144 579804 578156
rect 579856 578144 579862 578196
rect 3786 565836 3792 565888
rect 3844 565876 3850 565888
rect 4246 565876 4252 565888
rect 3844 565848 4252 565876
rect 3844 565836 3850 565848
rect 4246 565836 4252 565848
rect 4304 565836 4310 565888
rect 573726 564340 573732 564392
rect 573784 564380 573790 564392
rect 580166 564380 580172 564392
rect 573784 564352 580172 564380
rect 573784 564340 573790 564352
rect 580166 564340 580172 564352
rect 580224 564340 580230 564392
rect 573634 538160 573640 538212
rect 573692 538200 573698 538212
rect 580166 538200 580172 538212
rect 573692 538172 580172 538200
rect 573692 538160 573698 538172
rect 580166 538160 580172 538172
rect 580224 538160 580230 538212
rect 566826 511912 566832 511964
rect 566884 511952 566890 511964
rect 580166 511952 580172 511964
rect 566884 511924 580172 511952
rect 566884 511912 566890 511924
rect 580166 511912 580172 511924
rect 580224 511912 580230 511964
rect 575014 485732 575020 485784
rect 575072 485772 575078 485784
rect 579614 485772 579620 485784
rect 575072 485744 579620 485772
rect 575072 485732 575078 485744
rect 579614 485732 579620 485744
rect 579672 485732 579678 485784
rect 3326 463632 3332 463684
rect 3384 463672 3390 463684
rect 4430 463672 4436 463684
rect 3384 463644 4436 463672
rect 3384 463632 3390 463644
rect 4430 463632 4436 463644
rect 4488 463632 4494 463684
rect 577498 419432 577504 419484
rect 577556 419472 577562 419484
rect 579614 419472 579620 419484
rect 577556 419444 579620 419472
rect 577556 419432 577562 419444
rect 579614 419432 579620 419444
rect 579672 419432 579678 419484
rect 570690 405628 570696 405680
rect 570748 405668 570754 405680
rect 579798 405668 579804 405680
rect 570748 405640 579804 405668
rect 570748 405628 570754 405640
rect 579798 405628 579804 405640
rect 579856 405628 579862 405680
rect 574922 379448 574928 379500
rect 574980 379488 574986 379500
rect 579798 379488 579804 379500
rect 574980 379460 579804 379488
rect 574980 379448 574986 379460
rect 579798 379448 579804 379460
rect 579856 379448 579862 379500
rect 572070 353200 572076 353252
rect 572128 353240 572134 353252
rect 580166 353240 580172 353252
rect 572128 353212 580172 353240
rect 572128 353200 572134 353212
rect 580166 353200 580172 353212
rect 580224 353200 580230 353252
rect 570598 325592 570604 325644
rect 570656 325632 570662 325644
rect 580166 325632 580172 325644
rect 570656 325604 580172 325632
rect 570656 325592 570662 325604
rect 580166 325592 580172 325604
rect 580224 325592 580230 325644
rect 576302 313216 576308 313268
rect 576360 313256 576366 313268
rect 580166 313256 580172 313268
rect 576360 313228 580172 313256
rect 576360 313216 576366 313228
rect 580166 313216 580172 313228
rect 580224 313216 580230 313268
rect 569494 299412 569500 299464
rect 569552 299452 569558 299464
rect 580166 299452 580172 299464
rect 569552 299424 580172 299452
rect 569552 299412 569558 299424
rect 580166 299412 580172 299424
rect 580224 299412 580230 299464
rect 576210 273164 576216 273216
rect 576268 273204 576274 273216
rect 580166 273204 580172 273216
rect 576268 273176 580172 273204
rect 576268 273164 576274 273176
rect 580166 273164 580172 273176
rect 580224 273164 580230 273216
rect 574830 259360 574836 259412
rect 574888 259400 574894 259412
rect 579614 259400 579620 259412
rect 574888 259372 579620 259400
rect 574888 259360 574894 259372
rect 579614 259360 579620 259372
rect 579672 259360 579678 259412
rect 565354 245556 565360 245608
rect 565412 245596 565418 245608
rect 580166 245596 580172 245608
rect 565412 245568 580172 245596
rect 565412 245556 565418 245568
rect 580166 245556 580172 245568
rect 580224 245556 580230 245608
rect 569310 233180 569316 233232
rect 569368 233220 569374 233232
rect 580166 233220 580172 233232
rect 569368 233192 580172 233220
rect 569368 233180 569374 233192
rect 580166 233180 580172 233192
rect 580224 233180 580230 233232
rect 573542 219376 573548 219428
rect 573600 219416 573606 219428
rect 580166 219416 580172 219428
rect 573600 219388 580172 219416
rect 573600 219376 573606 219388
rect 580166 219376 580172 219388
rect 580224 219376 580230 219428
rect 566734 206932 566740 206984
rect 566792 206972 566798 206984
rect 579890 206972 579896 206984
rect 566792 206944 579896 206972
rect 566792 206932 566798 206944
rect 579890 206932 579896 206944
rect 579948 206932 579954 206984
rect 573450 179324 573456 179376
rect 573508 179364 573514 179376
rect 579982 179364 579988 179376
rect 573508 179336 579988 179364
rect 573508 179324 573514 179336
rect 579982 179324 579988 179336
rect 580040 179324 580046 179376
rect 566550 166948 566556 167000
rect 566608 166988 566614 167000
rect 580166 166988 580172 167000
rect 566608 166960 580172 166988
rect 566608 166948 566614 166960
rect 580166 166948 580172 166960
rect 580224 166948 580230 167000
rect 565170 139340 565176 139392
rect 565228 139380 565234 139392
rect 580166 139380 580172 139392
rect 565228 139352 580172 139380
rect 565228 139340 565234 139352
rect 580166 139340 580172 139352
rect 580224 139340 580230 139392
rect 573358 126896 573364 126948
rect 573416 126936 573422 126948
rect 580166 126936 580172 126948
rect 573416 126908 580172 126936
rect 573416 126896 573422 126908
rect 580166 126896 580172 126908
rect 580224 126896 580230 126948
rect 566642 113092 566648 113144
rect 566700 113132 566706 113144
rect 579798 113132 579804 113144
rect 566700 113104 579804 113132
rect 566700 113092 566706 113104
rect 579798 113092 579804 113104
rect 579856 113092 579862 113144
rect 571978 100648 571984 100700
rect 572036 100688 572042 100700
rect 580166 100688 580172 100700
rect 572036 100660 580172 100688
rect 572036 100648 572042 100660
rect 580166 100648 580172 100660
rect 580224 100648 580230 100700
rect 574738 86912 574744 86964
rect 574796 86952 574802 86964
rect 580166 86952 580172 86964
rect 574796 86924 580172 86952
rect 574796 86912 574802 86924
rect 580166 86912 580172 86924
rect 580224 86912 580230 86964
rect 565262 73108 565268 73160
rect 565320 73148 565326 73160
rect 580166 73148 580172 73160
rect 565320 73120 580172 73148
rect 565320 73108 565326 73120
rect 580166 73108 580172 73120
rect 580224 73108 580230 73160
rect 569402 60664 569408 60716
rect 569460 60704 569466 60716
rect 580166 60704 580172 60716
rect 569460 60676 580172 60704
rect 569460 60664 569466 60676
rect 580166 60664 580172 60676
rect 580224 60664 580230 60716
rect 576118 46860 576124 46912
rect 576176 46900 576182 46912
rect 580166 46900 580172 46912
rect 576176 46872 580172 46900
rect 576176 46860 576182 46872
rect 580166 46860 580172 46872
rect 580224 46860 580230 46912
rect 569218 33056 569224 33108
rect 569276 33096 569282 33108
rect 580166 33096 580172 33108
rect 569276 33068 580172 33096
rect 569276 33056 569282 33068
rect 580166 33056 580172 33068
rect 580224 33056 580230 33108
rect 566458 20612 566464 20664
rect 566516 20652 566522 20664
rect 579982 20652 579988 20664
rect 566516 20624 579988 20652
rect 566516 20612 566522 20624
rect 579982 20612 579988 20624
rect 580040 20612 580046 20664
rect 565078 6808 565084 6860
rect 565136 6848 565142 6860
rect 580166 6848 580172 6860
rect 565136 6820 580172 6848
rect 565136 6808 565142 6820
rect 580166 6808 580172 6820
rect 580224 6808 580230 6860
rect 563698 3000 563704 3052
rect 563756 3040 563762 3052
rect 583386 3040 583392 3052
rect 563756 3012 583392 3040
rect 563756 3000 563762 3012
rect 583386 3000 583392 3012
rect 583444 3000 583450 3052
rect 563514 2864 563520 2916
rect 563572 2904 563578 2916
rect 572714 2904 572720 2916
rect 563572 2876 572720 2904
rect 563572 2864 563578 2876
rect 572714 2864 572720 2876
rect 572772 2864 572778 2916
rect 569862 2796 569868 2848
rect 569920 2836 569926 2848
rect 576302 2836 576308 2848
rect 569920 2808 576308 2836
rect 569920 2796 569926 2808
rect 576302 2796 576308 2808
rect 576360 2796 576366 2848
rect 413741 1343 413799 1349
rect 413741 1309 413753 1343
rect 413787 1340 413799 1343
rect 425517 1343 425575 1349
rect 425517 1340 425529 1343
rect 413787 1312 425529 1340
rect 413787 1309 413799 1312
rect 413741 1303 413799 1309
rect 425517 1309 425529 1312
rect 425563 1309 425575 1343
rect 425517 1303 425575 1309
rect 487433 1343 487491 1349
rect 487433 1309 487445 1343
rect 487479 1340 487491 1343
rect 502981 1343 503039 1349
rect 502981 1340 502993 1343
rect 487479 1312 502993 1340
rect 487479 1309 487491 1312
rect 487433 1303 487491 1309
rect 502981 1309 502993 1312
rect 503027 1309 503039 1343
rect 502981 1303 503039 1309
rect 504637 1343 504695 1349
rect 504637 1309 504649 1343
rect 504683 1340 504695 1343
rect 520737 1343 520795 1349
rect 520737 1340 520749 1343
rect 504683 1312 520749 1340
rect 504683 1309 504695 1312
rect 504637 1303 504695 1309
rect 520737 1309 520749 1312
rect 520783 1309 520795 1343
rect 520737 1303 520795 1309
rect 462133 1275 462191 1281
rect 462133 1241 462145 1275
rect 462179 1272 462191 1275
rect 476945 1275 477003 1281
rect 476945 1272 476957 1275
rect 462179 1244 476957 1272
rect 462179 1241 462191 1244
rect 462133 1235 462191 1241
rect 476945 1241 476957 1244
rect 476991 1241 477003 1275
rect 476945 1235 477003 1241
rect 502337 1275 502395 1281
rect 502337 1241 502349 1275
rect 502383 1272 502395 1275
rect 518161 1275 518219 1281
rect 518161 1272 518173 1275
rect 502383 1244 518173 1272
rect 502383 1241 502395 1244
rect 502337 1235 502395 1241
rect 518161 1241 518173 1244
rect 518207 1241 518219 1275
rect 518161 1235 518219 1241
rect 518253 1275 518311 1281
rect 518253 1241 518265 1275
rect 518299 1272 518311 1275
rect 534537 1275 534595 1281
rect 534537 1272 534549 1275
rect 518299 1244 534549 1272
rect 518299 1241 518311 1244
rect 518253 1235 518311 1241
rect 534537 1241 534549 1244
rect 534583 1241 534595 1275
rect 534537 1235 534595 1241
rect 453577 1207 453635 1213
rect 453577 1173 453589 1207
rect 453623 1204 453635 1207
rect 466365 1207 466423 1213
rect 466365 1204 466377 1207
rect 453623 1176 466377 1204
rect 453623 1173 453635 1176
rect 453577 1167 453635 1173
rect 466365 1173 466377 1176
rect 466411 1173 466423 1207
rect 466365 1167 466423 1173
rect 468297 1207 468355 1213
rect 468297 1173 468309 1207
rect 468343 1204 468355 1207
rect 483017 1207 483075 1213
rect 483017 1204 483029 1207
rect 468343 1176 483029 1204
rect 468343 1173 468355 1176
rect 468297 1167 468355 1173
rect 483017 1173 483029 1176
rect 483063 1173 483075 1207
rect 483017 1167 483075 1173
rect 514389 1207 514447 1213
rect 514389 1173 514401 1207
rect 514435 1204 514447 1207
rect 531317 1207 531375 1213
rect 531317 1204 531329 1207
rect 514435 1176 531329 1204
rect 514435 1173 514447 1176
rect 514389 1167 514447 1173
rect 531317 1173 531329 1176
rect 531363 1173 531375 1207
rect 531317 1167 531375 1173
rect 545117 1207 545175 1213
rect 545117 1173 545129 1207
rect 545163 1204 545175 1207
rect 563241 1207 563299 1213
rect 563241 1204 563253 1207
rect 545163 1176 563253 1204
rect 545163 1173 545175 1176
rect 545117 1167 545175 1173
rect 563241 1173 563253 1176
rect 563287 1173 563299 1207
rect 563241 1167 563299 1173
rect 400033 1139 400091 1145
rect 400033 1105 400045 1139
rect 400079 1136 400091 1139
rect 404909 1139 404967 1145
rect 404909 1136 404921 1139
rect 400079 1108 404921 1136
rect 400079 1105 400091 1108
rect 400033 1099 400091 1105
rect 404909 1105 404921 1108
rect 404955 1105 404967 1139
rect 404909 1099 404967 1105
rect 439869 1139 439927 1145
rect 439869 1105 439881 1139
rect 439915 1136 439927 1139
rect 453485 1139 453543 1145
rect 453485 1136 453497 1139
rect 439915 1108 453497 1136
rect 439915 1105 439927 1108
rect 439869 1099 439927 1105
rect 453485 1105 453497 1108
rect 453531 1105 453543 1139
rect 453485 1099 453543 1105
rect 461489 1139 461547 1145
rect 461489 1105 461501 1139
rect 461535 1136 461547 1139
rect 475749 1139 475807 1145
rect 475749 1136 475761 1139
rect 461535 1108 475761 1136
rect 461535 1105 461547 1108
rect 461489 1099 461547 1105
rect 475749 1105 475761 1108
rect 475795 1105 475807 1139
rect 475749 1099 475807 1105
rect 507857 1139 507915 1145
rect 507857 1105 507869 1139
rect 507903 1136 507915 1139
rect 524233 1139 524291 1145
rect 524233 1136 524245 1139
rect 507903 1108 524245 1136
rect 507903 1105 507915 1108
rect 507857 1099 507915 1105
rect 524233 1105 524245 1108
rect 524279 1105 524291 1139
rect 524233 1099 524291 1105
rect 544197 1139 544255 1145
rect 544197 1105 544209 1139
rect 544243 1136 544255 1139
rect 562045 1139 562103 1145
rect 562045 1136 562057 1139
rect 544243 1108 562057 1136
rect 544243 1105 544255 1108
rect 544197 1099 544255 1105
rect 562045 1105 562057 1108
rect 562091 1105 562103 1139
rect 562045 1099 562103 1105
rect 388809 1071 388867 1077
rect 388809 1037 388821 1071
rect 388855 1068 388867 1071
rect 400217 1071 400275 1077
rect 400217 1068 400229 1071
rect 388855 1040 400229 1068
rect 388855 1037 388867 1040
rect 388809 1031 388867 1037
rect 400217 1037 400229 1040
rect 400263 1037 400275 1071
rect 400217 1031 400275 1037
rect 431865 1071 431923 1077
rect 431865 1037 431877 1071
rect 431911 1068 431923 1071
rect 445021 1071 445079 1077
rect 445021 1068 445033 1071
rect 431911 1040 445033 1068
rect 431911 1037 431923 1040
rect 431865 1031 431923 1037
rect 445021 1037 445033 1040
rect 445067 1037 445079 1071
rect 445021 1031 445079 1037
rect 467193 1071 467251 1077
rect 467193 1037 467205 1071
rect 467239 1068 467251 1071
rect 481729 1071 481787 1077
rect 481729 1068 481741 1071
rect 467239 1040 481741 1068
rect 467239 1037 467251 1040
rect 467193 1031 467251 1037
rect 481729 1037 481741 1040
rect 481775 1037 481787 1071
rect 481729 1031 481787 1037
rect 490929 1071 490987 1077
rect 490929 1037 490941 1071
rect 490975 1068 490987 1071
rect 506201 1071 506259 1077
rect 506201 1068 506213 1071
rect 490975 1040 506213 1068
rect 490975 1037 490987 1040
rect 490929 1031 490987 1037
rect 506201 1037 506213 1040
rect 506247 1037 506259 1071
rect 506201 1031 506259 1037
rect 516965 1071 517023 1077
rect 516965 1037 516977 1071
rect 517011 1068 517023 1071
rect 531133 1071 531191 1077
rect 531133 1068 531145 1071
rect 517011 1040 531145 1068
rect 517011 1037 517023 1040
rect 516965 1031 517023 1037
rect 531133 1037 531145 1040
rect 531179 1037 531191 1071
rect 531133 1031 531191 1037
rect 554593 1071 554651 1077
rect 554593 1037 554605 1071
rect 554639 1068 554651 1071
rect 563514 1068 563520 1080
rect 554639 1040 563520 1068
rect 554639 1037 554651 1040
rect 554593 1031 554651 1037
rect 563514 1028 563520 1040
rect 563572 1028 563578 1080
rect 415489 1003 415547 1009
rect 415489 1000 415501 1003
rect 408466 972 415501 1000
rect 370409 935 370467 941
rect 370409 901 370421 935
rect 370455 932 370467 935
rect 377493 935 377551 941
rect 377493 932 377505 935
rect 370455 904 377505 932
rect 370455 901 370467 904
rect 370409 895 370467 901
rect 377493 901 377505 904
rect 377539 901 377551 935
rect 404817 935 404875 941
rect 404817 932 404829 935
rect 377493 895 377551 901
rect 404556 904 404829 932
rect 375193 867 375251 873
rect 375193 833 375205 867
rect 375239 864 375251 867
rect 393317 867 393375 873
rect 375239 836 386000 864
rect 375239 833 375251 836
rect 375193 827 375251 833
rect 312633 799 312691 805
rect 312633 796 312645 799
rect 304966 768 312645 796
rect 7469 731 7527 737
rect 7469 697 7481 731
rect 7515 728 7527 731
rect 240505 731 240563 737
rect 240505 728 240517 731
rect 7515 700 11560 728
rect 7515 697 7527 700
rect 7469 691 7527 697
rect 11532 672 11560 700
rect 213886 700 218008 728
rect 213886 672 213914 700
rect 217980 672 218008 700
rect 237346 700 240517 728
rect 1670 620 1676 672
rect 1728 660 1734 672
rect 5350 660 5356 672
rect 1728 632 5356 660
rect 1728 620 1734 632
rect 5350 620 5356 632
rect 5408 620 5414 672
rect 6454 620 6460 672
rect 6512 660 6518 672
rect 10042 660 10048 672
rect 6512 632 10048 660
rect 6512 620 6518 632
rect 10042 620 10048 632
rect 10100 620 10106 672
rect 10152 632 11468 660
rect 566 552 572 604
rect 624 592 630 604
rect 4338 592 4344 604
rect 624 564 4344 592
rect 624 552 630 564
rect 4338 552 4344 564
rect 4396 552 4402 604
rect 5258 552 5264 604
rect 5316 592 5322 604
rect 8846 592 8852 604
rect 5316 564 8852 592
rect 5316 552 5322 564
rect 8846 552 8852 564
rect 8904 552 8910 604
rect 7466 524 7472 536
rect 7427 496 7472 524
rect 7466 484 7472 496
rect 7524 484 7530 536
rect 8570 484 8576 536
rect 8628 524 8634 536
rect 10152 524 10180 632
rect 11146 552 11152 604
rect 11204 552 11210 604
rect 11440 592 11468 632
rect 11514 620 11520 672
rect 11572 620 11578 672
rect 19426 620 19432 672
rect 19484 660 19490 672
rect 22370 660 22376 672
rect 19484 632 22376 660
rect 19484 620 19490 632
rect 22370 620 22376 632
rect 22428 620 22434 672
rect 24854 660 24860 672
rect 22480 632 24860 660
rect 11440 564 11836 592
rect 8628 496 10180 524
rect 11164 524 11192 552
rect 11808 524 11836 564
rect 12342 552 12348 604
rect 12400 592 12406 604
rect 15562 592 15568 604
rect 12400 564 15568 592
rect 12400 552 12406 564
rect 15562 552 15568 564
rect 15620 552 15626 604
rect 21818 552 21824 604
rect 21876 592 21882 604
rect 22480 592 22508 632
rect 24854 620 24860 632
rect 24912 620 24918 672
rect 25314 620 25320 672
rect 25372 660 25378 672
rect 28074 660 28080 672
rect 25372 632 28080 660
rect 25372 620 25378 632
rect 28074 620 28080 632
rect 28132 620 28138 672
rect 28718 620 28724 672
rect 28776 660 28782 672
rect 29178 660 29184 672
rect 28776 632 29184 660
rect 28776 620 28782 632
rect 29178 620 29184 632
rect 29236 620 29242 672
rect 31294 620 31300 672
rect 31352 660 31358 672
rect 33778 660 33784 672
rect 31352 632 33784 660
rect 31352 620 31358 632
rect 33778 620 33784 632
rect 33836 620 33842 672
rect 34790 620 34796 672
rect 34848 660 34854 672
rect 37274 660 37280 672
rect 34848 632 37280 660
rect 34848 620 34854 632
rect 37274 620 37280 632
rect 37332 620 37338 672
rect 38378 620 38384 672
rect 38436 660 38442 672
rect 38436 632 38654 660
rect 38436 620 38442 632
rect 21876 564 22508 592
rect 21876 552 21882 564
rect 23014 552 23020 604
rect 23072 592 23078 604
rect 25774 592 25780 604
rect 23072 564 25780 592
rect 23072 552 23078 564
rect 25774 552 25780 564
rect 25832 552 25838 604
rect 28810 552 28816 604
rect 28868 592 28874 604
rect 28868 564 29040 592
rect 28868 552 28874 564
rect 12618 524 12624 536
rect 11164 496 11284 524
rect 11808 496 12624 524
rect 8628 484 8634 496
rect 3234 416 3240 468
rect 3292 456 3298 468
rect 6638 456 6644 468
rect 3292 428 6644 456
rect 3292 416 3298 428
rect 6638 416 6644 428
rect 6696 416 6702 468
rect 11256 456 11284 496
rect 12618 484 12624 496
rect 12676 484 12682 536
rect 13262 484 13268 536
rect 13320 524 13326 536
rect 16666 524 16672 536
rect 13320 496 16672 524
rect 13320 484 13326 496
rect 16666 484 16672 496
rect 16724 484 16730 536
rect 17402 484 17408 536
rect 17460 524 17466 536
rect 20070 524 20076 536
rect 17460 496 20076 524
rect 17460 484 17466 496
rect 20070 484 20076 496
rect 20128 484 20134 536
rect 29012 524 29040 564
rect 30098 552 30104 604
rect 30156 592 30162 604
rect 32582 592 32588 604
rect 30156 564 32588 592
rect 30156 552 30162 564
rect 32582 552 32588 564
rect 32640 552 32646 604
rect 33594 552 33600 604
rect 33652 592 33658 604
rect 36078 592 36084 604
rect 33652 564 36084 592
rect 33652 552 33658 564
rect 36078 552 36084 564
rect 36136 552 36142 604
rect 37182 552 37188 604
rect 37240 552 37246 604
rect 38626 592 38654 632
rect 40678 620 40684 672
rect 40736 660 40742 672
rect 42794 660 42800 672
rect 40736 632 42800 660
rect 40736 620 40742 632
rect 42794 620 42800 632
rect 42852 620 42858 672
rect 46658 620 46664 672
rect 46716 660 46722 672
rect 48498 660 48504 672
rect 46716 632 48504 660
rect 46716 620 46722 632
rect 48498 620 48504 632
rect 48556 620 48562 672
rect 48958 620 48964 672
rect 49016 660 49022 672
rect 50798 660 50804 672
rect 49016 632 50804 660
rect 49016 620 49022 632
rect 50798 620 50804 632
rect 50856 620 50862 672
rect 53742 620 53748 672
rect 53800 660 53806 672
rect 55398 660 55404 672
rect 53800 632 55404 660
rect 53800 620 53806 632
rect 55398 620 55404 632
rect 55456 620 55462 672
rect 64322 620 64328 672
rect 64380 660 64386 672
rect 65610 660 65616 672
rect 64380 632 65616 660
rect 64380 620 64386 632
rect 65610 620 65616 632
rect 65668 620 65674 672
rect 66714 620 66720 672
rect 66772 660 66778 672
rect 68002 660 68008 672
rect 66772 632 68008 660
rect 66772 620 66778 632
rect 68002 620 68008 632
rect 68060 620 68066 672
rect 69106 620 69112 672
rect 69164 660 69170 672
rect 70578 660 70584 672
rect 69164 632 70584 660
rect 69164 620 69170 632
rect 70578 620 70584 632
rect 70636 620 70642 672
rect 133230 620 133236 672
rect 133288 660 133294 672
rect 134150 660 134156 672
rect 133288 632 134156 660
rect 133288 620 133294 632
rect 134150 620 134156 632
rect 134208 620 134214 672
rect 136174 620 136180 672
rect 136232 660 136238 672
rect 137646 660 137652 672
rect 136232 632 137652 660
rect 136232 620 136238 632
rect 137646 620 137652 632
rect 137704 620 137710 672
rect 138750 620 138756 672
rect 138808 660 138814 672
rect 140038 660 140044 672
rect 138808 632 140044 660
rect 138808 620 138814 632
rect 140038 620 140044 632
rect 140096 620 140102 672
rect 151354 620 151360 672
rect 151412 660 151418 672
rect 153010 660 153016 672
rect 151412 632 153016 660
rect 151412 620 151418 632
rect 153010 620 153016 632
rect 153068 620 153074 672
rect 153654 620 153660 672
rect 153712 660 153718 672
rect 155402 660 155408 672
rect 153712 632 155408 660
rect 153712 620 153718 632
rect 155402 620 155408 632
rect 155460 620 155466 672
rect 162762 620 162768 672
rect 162820 660 162826 672
rect 164878 660 164884 672
rect 162820 632 164884 660
rect 162820 620 162826 632
rect 164878 620 164884 632
rect 164936 620 164942 672
rect 166074 660 166080 672
rect 165908 632 166080 660
rect 40770 592 40776 604
rect 38626 564 40776 592
rect 40770 552 40776 564
rect 40828 552 40834 604
rect 41874 552 41880 604
rect 41932 592 41938 604
rect 43990 592 43996 604
rect 41932 564 43996 592
rect 41932 552 41938 564
rect 43990 552 43996 564
rect 44048 552 44054 604
rect 47854 552 47860 604
rect 47912 592 47918 604
rect 49602 592 49608 604
rect 47912 564 49608 592
rect 47912 552 47918 564
rect 49602 552 49608 564
rect 49660 552 49666 604
rect 50154 552 50160 604
rect 50212 552 50218 604
rect 51350 552 51356 604
rect 51408 592 51414 604
rect 53006 592 53012 604
rect 51408 564 53012 592
rect 51408 552 51414 564
rect 53006 552 53012 564
rect 53064 552 53070 604
rect 54938 552 54944 604
rect 54996 592 55002 604
rect 56410 592 56416 604
rect 54996 564 56416 592
rect 54996 552 55002 564
rect 56410 552 56416 564
rect 56468 552 56474 604
rect 60826 552 60832 604
rect 60884 592 60890 604
rect 62114 592 62120 604
rect 60884 564 62120 592
rect 60884 552 60890 564
rect 62114 552 62120 564
rect 62172 552 62178 604
rect 65518 552 65524 604
rect 65576 592 65582 604
rect 66806 592 66812 604
rect 65576 564 66812 592
rect 65576 552 65582 564
rect 66806 552 66812 564
rect 66864 552 66870 604
rect 70302 552 70308 604
rect 70360 592 70366 604
rect 71222 592 71228 604
rect 70360 564 71228 592
rect 70360 552 70366 564
rect 71222 552 71228 564
rect 71280 552 71286 604
rect 76190 552 76196 604
rect 76248 592 76254 604
rect 76926 592 76932 604
rect 76248 564 76932 592
rect 76248 552 76254 564
rect 76926 552 76932 564
rect 76984 552 76990 604
rect 77386 552 77392 604
rect 77444 592 77450 604
rect 78030 592 78036 604
rect 77444 564 78036 592
rect 77444 552 77450 564
rect 78030 552 78036 564
rect 78088 552 78094 604
rect 78582 552 78588 604
rect 78640 592 78646 604
rect 79134 592 79140 604
rect 78640 564 79140 592
rect 78640 552 78646 564
rect 79134 552 79140 564
rect 79192 552 79198 604
rect 79686 552 79692 604
rect 79744 592 79750 604
rect 80330 592 80336 604
rect 79744 564 80336 592
rect 79744 552 79750 564
rect 80330 552 80336 564
rect 80388 552 80394 604
rect 80882 552 80888 604
rect 80940 592 80946 604
rect 81434 592 81440 604
rect 80940 564 81440 592
rect 80940 552 80946 564
rect 81434 552 81440 564
rect 81492 552 81498 604
rect 82078 552 82084 604
rect 82136 592 82142 604
rect 82722 592 82728 604
rect 82136 564 82728 592
rect 82136 552 82142 564
rect 82722 552 82728 564
rect 82780 552 82786 604
rect 121822 552 121828 604
rect 121880 592 121886 604
rect 122282 592 122288 604
rect 121880 564 122288 592
rect 121880 552 121886 564
rect 122282 552 122288 564
rect 122340 552 122346 604
rect 124122 552 124128 604
rect 124180 592 124186 604
rect 124674 592 124680 604
rect 124180 564 124680 592
rect 124180 552 124186 564
rect 124674 552 124680 564
rect 124732 552 124738 604
rect 125226 552 125232 604
rect 125284 592 125290 604
rect 125870 592 125876 604
rect 125284 564 125876 592
rect 125284 552 125290 564
rect 125870 552 125876 564
rect 125928 552 125934 604
rect 126422 552 126428 604
rect 126480 592 126486 604
rect 126974 592 126980 604
rect 126480 564 126980 592
rect 126480 552 126486 564
rect 126974 552 126980 564
rect 127032 552 127038 604
rect 127526 552 127532 604
rect 127584 592 127590 604
rect 128170 592 128176 604
rect 127584 564 128176 592
rect 127584 552 127590 564
rect 128170 552 128176 564
rect 128228 552 128234 604
rect 128630 552 128636 604
rect 128688 592 128694 604
rect 129366 592 129372 604
rect 128688 564 129372 592
rect 128688 552 128694 564
rect 129366 552 129372 564
rect 129424 552 129430 604
rect 133874 552 133880 604
rect 133932 592 133938 604
rect 135254 592 135260 604
rect 133932 564 135260 592
rect 133932 552 133938 564
rect 135254 552 135260 564
rect 135312 552 135318 604
rect 136450 552 136456 604
rect 136508 552 136514 604
rect 137554 552 137560 604
rect 137612 592 137618 604
rect 138842 592 138848 604
rect 137612 564 138848 592
rect 137612 552 137618 564
rect 138842 552 138848 564
rect 138900 552 138906 604
rect 139946 552 139952 604
rect 140004 592 140010 604
rect 141234 592 141240 604
rect 140004 564 141240 592
rect 140004 552 140010 564
rect 141234 552 141240 564
rect 141292 552 141298 604
rect 144546 552 144552 604
rect 144604 592 144610 604
rect 145926 592 145932 604
rect 144604 564 145932 592
rect 144604 552 144610 564
rect 145926 552 145932 564
rect 145984 552 145990 604
rect 146846 552 146852 604
rect 146904 592 146910 604
rect 148318 592 148324 604
rect 146904 564 148324 592
rect 146904 552 146910 564
rect 148318 552 148324 564
rect 148376 552 148382 604
rect 152550 552 152556 604
rect 152608 592 152614 604
rect 154206 592 154212 604
rect 152608 564 154212 592
rect 152608 552 152614 564
rect 154206 552 154212 564
rect 154264 552 154270 604
rect 154758 552 154764 604
rect 154816 592 154822 604
rect 156598 592 156604 604
rect 154816 564 156604 592
rect 154816 552 154822 564
rect 156598 552 156604 564
rect 156656 552 156662 604
rect 157058 552 157064 604
rect 157116 592 157122 604
rect 158898 592 158904 604
rect 157116 564 158904 592
rect 157116 552 157122 564
rect 158898 552 158904 564
rect 158956 552 158962 604
rect 161566 552 161572 604
rect 161624 592 161630 604
rect 163682 592 163688 604
rect 161624 564 163688 592
rect 161624 552 161630 564
rect 163682 552 163688 564
rect 163740 552 163746 604
rect 31662 524 31668 536
rect 29012 496 31668 524
rect 31662 484 31668 496
rect 31720 484 31726 536
rect 33226 484 33232 536
rect 33284 524 33290 536
rect 34974 524 34980 536
rect 33284 496 34980 524
rect 33284 484 33290 496
rect 34974 484 34980 496
rect 35032 484 35038 536
rect 14458 456 14464 468
rect 11256 428 14464 456
rect 14458 416 14464 428
rect 14516 416 14522 468
rect 24394 416 24400 468
rect 24452 456 24458 468
rect 26878 456 26884 468
rect 24452 428 26884 456
rect 24452 416 24458 428
rect 26878 416 26884 428
rect 26936 416 26942 468
rect 37200 456 37228 552
rect 50172 524 50200 552
rect 51902 524 51908 536
rect 50172 496 51908 524
rect 51902 484 51908 496
rect 51960 484 51966 536
rect 63494 484 63500 536
rect 63552 524 63558 536
rect 64506 524 64512 536
rect 63552 496 64512 524
rect 63552 484 63558 496
rect 64506 484 64512 496
rect 64564 484 64570 536
rect 67726 484 67732 536
rect 67784 524 67790 536
rect 69382 524 69388 536
rect 67784 496 69388 524
rect 67784 484 67790 496
rect 69382 484 69388 496
rect 69440 484 69446 536
rect 134978 484 134984 536
rect 135036 524 135042 536
rect 136468 524 136496 552
rect 135036 496 136496 524
rect 135036 484 135042 496
rect 141050 484 141056 536
rect 141108 524 141114 536
rect 142062 524 142068 536
rect 141108 496 142068 524
rect 141108 484 141114 496
rect 142062 484 142068 496
rect 142120 484 142126 536
rect 158162 484 158168 536
rect 158220 524 158226 536
rect 159726 524 159732 536
rect 158220 496 159732 524
rect 158220 484 158226 496
rect 159726 484 159732 496
rect 159784 484 159790 536
rect 39850 456 39856 468
rect 37200 428 39856 456
rect 39850 416 39856 428
rect 39908 416 39914 468
rect 163406 416 163412 468
rect 163464 456 163470 468
rect 165908 456 165936 632
rect 166074 620 166080 632
rect 166132 620 166138 672
rect 167086 620 167092 672
rect 167144 660 167150 672
rect 169570 660 169576 672
rect 167144 632 169576 660
rect 167144 620 167150 632
rect 169570 620 169576 632
rect 169628 620 169634 672
rect 180886 620 180892 672
rect 180944 660 180950 672
rect 183738 660 183744 672
rect 180944 632 183744 660
rect 180944 620 180950 632
rect 183738 620 183744 632
rect 183796 620 183802 672
rect 189994 620 190000 672
rect 190052 660 190058 672
rect 193214 660 193220 672
rect 190052 632 193220 660
rect 190052 620 190058 632
rect 193214 620 193220 632
rect 193272 620 193278 672
rect 194318 620 194324 672
rect 194376 660 194382 672
rect 197906 660 197912 672
rect 194376 632 197912 660
rect 194376 620 194382 632
rect 197906 620 197912 632
rect 197964 620 197970 672
rect 213822 620 213828 672
rect 213880 632 213914 672
rect 215662 660 215668 672
rect 214392 632 215668 660
rect 213880 620 213886 632
rect 165982 552 165988 604
rect 166040 592 166046 604
rect 168374 592 168380 604
rect 166040 564 168380 592
rect 166040 552 166046 564
rect 168374 552 168380 564
rect 168432 552 168438 604
rect 170674 552 170680 604
rect 170732 592 170738 604
rect 173158 592 173164 604
rect 170732 564 173164 592
rect 170732 552 170738 564
rect 173158 552 173164 564
rect 173216 552 173222 604
rect 179782 552 179788 604
rect 179840 592 179846 604
rect 182542 592 182548 604
rect 179840 564 182548 592
rect 179840 552 179846 564
rect 182542 552 182548 564
rect 182600 552 182606 604
rect 183186 552 183192 604
rect 183244 592 183250 604
rect 186130 592 186136 604
rect 183244 564 186136 592
rect 183244 552 183250 564
rect 186130 552 186136 564
rect 186188 552 186194 604
rect 188798 552 188804 604
rect 188856 592 188862 604
rect 188856 564 192248 592
rect 188856 552 188862 564
rect 192220 536 192248 564
rect 192294 552 192300 604
rect 192352 592 192358 604
rect 195606 592 195612 604
rect 192352 564 195612 592
rect 192352 552 192358 564
rect 195606 552 195612 564
rect 195664 552 195670 604
rect 196894 552 196900 604
rect 196952 552 196958 604
rect 205726 552 205732 604
rect 205784 592 205790 604
rect 209774 592 209780 604
rect 205784 564 209780 592
rect 205784 552 205790 564
rect 209774 552 209780 564
rect 209832 552 209838 604
rect 210418 552 210424 604
rect 210476 592 210482 604
rect 210476 564 211154 592
rect 210476 552 210482 564
rect 187694 484 187700 536
rect 187752 524 187758 536
rect 191006 524 191012 536
rect 187752 496 191012 524
rect 187752 484 187758 496
rect 191006 484 191012 496
rect 191064 484 191070 536
rect 192202 484 192208 536
rect 192260 484 192266 536
rect 192938 484 192944 536
rect 192996 524 193002 536
rect 196912 524 196940 552
rect 192996 496 196940 524
rect 211126 524 211154 564
rect 211614 552 211620 604
rect 211672 592 211678 604
rect 214392 592 214420 632
rect 215662 620 215668 632
rect 215720 620 215726 672
rect 217962 620 217968 672
rect 218020 620 218026 672
rect 218422 620 218428 672
rect 218480 660 218486 672
rect 222746 660 222752 672
rect 218480 632 222752 660
rect 218480 620 218486 632
rect 222746 620 222752 632
rect 222804 620 222810 672
rect 226334 660 226340 672
rect 223868 632 226340 660
rect 211672 564 214420 592
rect 211672 552 211678 564
rect 214466 552 214472 604
rect 214524 552 214530 604
rect 220170 552 220176 604
rect 220228 592 220234 604
rect 220446 592 220452 604
rect 220228 564 220452 592
rect 220228 552 220234 564
rect 220446 552 220452 564
rect 220504 552 220510 604
rect 221826 552 221832 604
rect 221884 592 221890 604
rect 223868 592 223896 632
rect 226334 620 226340 632
rect 226392 620 226398 672
rect 231026 660 231032 672
rect 228192 632 231032 660
rect 221884 564 223896 592
rect 221884 552 221890 564
rect 223942 552 223948 604
rect 224000 552 224006 604
rect 226150 552 226156 604
rect 226208 592 226214 604
rect 228192 592 228220 632
rect 231026 620 231032 632
rect 231084 620 231090 672
rect 234614 660 234620 672
rect 231780 632 234620 660
rect 229830 592 229836 604
rect 226208 564 228220 592
rect 229066 564 229836 592
rect 226208 552 226214 564
rect 214484 524 214512 552
rect 211126 496 214512 524
rect 192996 484 193002 496
rect 219526 484 219532 536
rect 219584 524 219590 536
rect 223960 524 223988 552
rect 219584 496 223988 524
rect 219584 484 219590 496
rect 224770 484 224776 536
rect 224828 524 224834 536
rect 229066 524 229094 564
rect 229830 552 229836 564
rect 229888 552 229894 604
rect 224828 496 229094 524
rect 224828 484 224834 496
rect 229646 484 229652 536
rect 229704 524 229710 536
rect 231780 524 231808 632
rect 234614 620 234620 632
rect 234672 620 234678 672
rect 235442 620 235448 672
rect 235500 660 235506 672
rect 237346 660 237374 700
rect 240505 697 240517 700
rect 240551 697 240563 731
rect 304966 728 304994 768
rect 312633 765 312645 768
rect 312679 765 312691 799
rect 364705 799 364763 805
rect 312633 759 312691 765
rect 328472 768 333974 796
rect 311437 731 311495 737
rect 311437 728 311449 731
rect 240505 691 240563 697
rect 275986 700 279556 728
rect 235500 632 237374 660
rect 235500 620 235506 632
rect 237742 620 237748 672
rect 237800 660 237806 672
rect 242894 660 242900 672
rect 237800 632 242900 660
rect 237800 620 237806 632
rect 242894 620 242900 632
rect 242952 620 242958 672
rect 247954 620 247960 672
rect 248012 660 248018 672
rect 253474 660 253480 672
rect 248012 632 253480 660
rect 248012 620 248018 632
rect 253474 620 253480 632
rect 253532 620 253538 672
rect 255501 663 255559 669
rect 255501 629 255513 663
rect 255547 660 255559 663
rect 257062 660 257068 672
rect 255547 632 257068 660
rect 255547 629 255559 632
rect 255501 623 255559 629
rect 257062 620 257068 632
rect 257120 620 257126 672
rect 257246 620 257252 672
rect 257304 660 257310 672
rect 258258 660 258264 672
rect 257304 632 258264 660
rect 257304 620 257310 632
rect 258258 620 258264 632
rect 258316 620 258322 672
rect 260650 660 260656 672
rect 259288 632 260656 660
rect 231854 552 231860 604
rect 231912 592 231918 604
rect 237006 592 237012 604
rect 231912 564 237012 592
rect 231912 552 231918 564
rect 237006 552 237012 564
rect 237064 552 237070 604
rect 238110 552 238116 604
rect 238168 552 238174 604
rect 239306 592 239312 604
rect 238404 564 239312 592
rect 229704 496 231808 524
rect 229704 484 229710 496
rect 233142 484 233148 536
rect 233200 524 233206 536
rect 238128 524 238156 552
rect 233200 496 238156 524
rect 233200 484 233206 496
rect 163464 428 165936 456
rect 163464 416 163470 428
rect 212718 416 212724 468
rect 212776 456 212782 468
rect 216582 456 216588 468
rect 212776 428 216588 456
rect 212776 416 212782 428
rect 216582 416 216588 428
rect 216640 416 216646 468
rect 234338 416 234344 468
rect 234396 456 234402 468
rect 238404 456 238432 564
rect 239306 552 239312 564
rect 239364 552 239370 604
rect 240502 592 240508 604
rect 240463 564 240508 592
rect 240502 552 240508 564
rect 240560 552 240566 604
rect 241146 552 241152 604
rect 241204 592 241210 604
rect 246022 592 246028 604
rect 241204 564 246028 592
rect 241204 552 241210 564
rect 246022 552 246028 564
rect 246080 552 246086 604
rect 249978 552 249984 604
rect 250036 552 250042 604
rect 251174 552 251180 604
rect 251232 552 251238 604
rect 252370 552 252376 604
rect 252428 552 252434 604
rect 253382 552 253388 604
rect 253440 552 253446 604
rect 254578 552 254584 604
rect 254636 592 254642 604
rect 259288 592 259316 632
rect 260650 620 260656 632
rect 260708 620 260714 672
rect 262674 620 262680 672
rect 262732 660 262738 672
rect 268838 660 268844 672
rect 262732 632 268844 660
rect 262732 620 262738 632
rect 268838 620 268844 632
rect 268896 620 268902 672
rect 272886 620 272892 672
rect 272944 660 272950 672
rect 275986 660 276014 700
rect 272944 632 276014 660
rect 272944 620 272950 632
rect 279528 604 279556 700
rect 285646 700 287054 728
rect 279697 663 279755 669
rect 279697 629 279709 663
rect 279743 660 279755 663
rect 285398 660 285404 672
rect 279743 632 285404 660
rect 279743 629 279755 632
rect 279697 623 279755 629
rect 285398 620 285404 632
rect 285456 620 285462 672
rect 259454 592 259460 604
rect 254636 564 259316 592
rect 259380 564 259460 592
rect 254636 552 254642 564
rect 244550 484 244556 536
rect 244608 524 244614 536
rect 249996 524 250024 552
rect 251192 524 251220 552
rect 244608 496 250024 524
rect 251146 496 251220 524
rect 244608 484 244614 496
rect 234396 428 238432 456
rect 234396 416 234402 428
rect 239950 416 239956 468
rect 240008 456 240014 468
rect 244918 456 244924 468
rect 240008 428 244924 456
rect 240008 416 240014 428
rect 244918 416 244924 428
rect 244976 416 244982 468
rect 245654 416 245660 468
rect 245712 456 245718 468
rect 251146 456 251174 496
rect 245712 428 251174 456
rect 245712 416 245718 428
rect 14550 348 14556 400
rect 14608 388 14614 400
rect 17862 388 17868 400
rect 14608 360 17868 388
rect 14608 348 14614 360
rect 17862 348 17868 360
rect 17920 348 17926 400
rect 39298 348 39304 400
rect 39356 388 39362 400
rect 42150 388 42156 400
rect 39356 360 42156 388
rect 39356 348 39362 360
rect 42150 348 42156 360
rect 42208 348 42214 400
rect 42886 348 42892 400
rect 42944 388 42950 400
rect 45094 388 45100 400
rect 42944 360 45100 388
rect 42944 348 42950 360
rect 45094 348 45100 360
rect 45152 348 45158 400
rect 71314 348 71320 400
rect 71372 388 71378 400
rect 72326 388 72332 400
rect 71372 360 72332 388
rect 71372 348 71378 360
rect 72326 348 72332 360
rect 72384 348 72390 400
rect 72418 348 72424 400
rect 72476 388 72482 400
rect 73522 388 73528 400
rect 72476 360 73528 388
rect 72476 348 72482 360
rect 73522 348 73528 360
rect 73580 348 73586 400
rect 73614 348 73620 400
rect 73672 388 73678 400
rect 74626 388 74632 400
rect 73672 360 74632 388
rect 73672 348 73678 360
rect 74626 348 74632 360
rect 74684 348 74690 400
rect 130930 348 130936 400
rect 130988 388 130994 400
rect 131942 388 131948 400
rect 130988 360 131948 388
rect 130988 348 130994 360
rect 131942 348 131948 360
rect 132000 348 132006 400
rect 132034 348 132040 400
rect 132092 388 132098 400
rect 133138 388 133144 400
rect 132092 360 133144 388
rect 132092 348 132098 360
rect 133138 348 133144 360
rect 133196 348 133202 400
rect 160462 348 160468 400
rect 160520 388 160526 400
rect 162670 388 162676 400
rect 160520 360 162676 388
rect 160520 348 160526 360
rect 162670 348 162676 360
rect 162728 348 162734 400
rect 220170 348 220176 400
rect 220228 388 220234 400
rect 225322 388 225328 400
rect 220228 360 225328 388
rect 220228 348 220234 360
rect 225322 348 225328 360
rect 225380 348 225386 400
rect 246758 348 246764 400
rect 246816 388 246822 400
rect 252388 388 252416 552
rect 253400 524 253428 552
rect 259380 524 259408 564
rect 259454 552 259460 564
rect 259512 552 259518 604
rect 260466 552 260472 604
rect 260524 592 260530 604
rect 266538 592 266544 604
rect 260524 564 266544 592
rect 260524 552 260530 564
rect 266538 552 266544 564
rect 266596 552 266602 604
rect 270034 552 270040 604
rect 270092 552 270098 604
rect 274082 552 274088 604
rect 274140 592 274146 604
rect 274140 564 278084 592
rect 274140 552 274146 564
rect 253400 496 259408 524
rect 263686 484 263692 536
rect 263744 524 263750 536
rect 270052 524 270080 552
rect 263744 496 270080 524
rect 263744 484 263750 496
rect 270494 484 270500 536
rect 270552 524 270558 536
rect 276750 524 276756 536
rect 270552 496 276756 524
rect 270552 484 270558 496
rect 276750 484 276756 496
rect 276808 484 276814 536
rect 278056 524 278084 564
rect 279510 552 279516 604
rect 279568 552 279574 604
rect 279605 595 279663 601
rect 279605 561 279617 595
rect 279651 592 279663 595
rect 284294 592 284300 604
rect 279651 564 284300 592
rect 279651 561 279663 564
rect 279605 555 279663 561
rect 284294 552 284300 564
rect 284352 552 284358 604
rect 278056 496 280154 524
rect 257982 416 257988 468
rect 258040 456 258046 468
rect 258040 416 258074 456
rect 259270 416 259276 468
rect 259328 456 259334 468
rect 264974 456 264980 468
rect 259328 428 264980 456
rect 259328 416 259334 428
rect 264974 416 264980 428
rect 265032 416 265038 468
rect 268378 416 268384 468
rect 268436 456 268442 468
rect 274542 456 274548 468
rect 268436 428 274548 456
rect 268436 416 268442 428
rect 274542 416 274548 428
rect 274600 416 274606 468
rect 277486 416 277492 468
rect 277544 456 277550 468
rect 279605 459 279663 465
rect 279605 456 279617 459
rect 277544 428 279617 456
rect 277544 416 277550 428
rect 279605 425 279617 428
rect 279651 425 279663 459
rect 280126 456 280154 496
rect 281534 484 281540 536
rect 281592 524 281598 536
rect 285646 524 285674 700
rect 287026 660 287054 700
rect 292546 700 298508 728
rect 288986 660 288992 672
rect 287026 632 288992 660
rect 288986 620 288992 632
rect 289044 620 289050 672
rect 291102 620 291108 672
rect 291160 660 291166 672
rect 292546 660 292574 700
rect 298480 672 298508 700
rect 304736 700 304994 728
rect 307036 700 311449 728
rect 304736 672 304764 700
rect 291160 632 292574 660
rect 291160 620 291166 632
rect 293402 620 293408 672
rect 293460 660 293466 672
rect 298373 663 298431 669
rect 298373 660 298385 663
rect 293460 632 298385 660
rect 293460 620 293466 632
rect 298373 629 298385 632
rect 298419 629 298431 663
rect 298373 623 298431 629
rect 298462 620 298468 672
rect 298520 620 298526 672
rect 298557 663 298615 669
rect 298557 629 298569 663
rect 298603 660 298615 663
rect 300762 660 300768 672
rect 298603 632 300768 660
rect 298603 629 298615 632
rect 298557 623 298615 629
rect 300762 620 300768 632
rect 300820 620 300826 672
rect 301314 620 301320 672
rect 301372 660 301378 672
rect 301372 632 303568 660
rect 301372 620 301378 632
rect 288802 552 288808 604
rect 288860 592 288866 604
rect 296070 592 296076 604
rect 288860 564 296076 592
rect 288860 552 288866 564
rect 296070 552 296076 564
rect 296128 552 296134 604
rect 303154 552 303160 604
rect 303212 552 303218 604
rect 281592 496 285674 524
rect 281592 484 281598 496
rect 287606 484 287612 536
rect 287664 524 287670 536
rect 293862 524 293868 536
rect 287664 496 293868 524
rect 287664 484 287670 496
rect 293862 484 293868 496
rect 293920 484 293926 536
rect 295610 484 295616 536
rect 295668 524 295674 536
rect 303172 524 303200 552
rect 295668 496 303200 524
rect 303540 524 303568 632
rect 304718 620 304724 672
rect 304776 620 304782 672
rect 303614 552 303620 604
rect 303672 592 303678 604
rect 307036 592 307064 700
rect 311437 697 311449 700
rect 311483 697 311495 731
rect 311437 691 311495 697
rect 318720 700 326844 728
rect 318720 672 318748 700
rect 326816 672 326844 700
rect 328472 672 328500 768
rect 333946 728 333974 768
rect 364705 765 364717 799
rect 364751 796 364763 799
rect 364751 768 370728 796
rect 364751 765 364763 768
rect 364705 759 364763 765
rect 333946 700 337516 728
rect 337488 672 337516 700
rect 344986 700 350488 728
rect 307938 660 307944 672
rect 307899 632 307944 660
rect 307938 620 307944 632
rect 307996 620 308002 672
rect 309962 620 309968 672
rect 310020 660 310026 672
rect 318518 660 318524 672
rect 310020 632 314654 660
rect 310020 620 310026 632
rect 303672 564 307064 592
rect 303672 552 303678 564
rect 309042 552 309048 604
rect 309100 552 309106 604
rect 310238 552 310244 604
rect 310296 552 310302 604
rect 311434 592 311440 604
rect 311395 564 311440 592
rect 311434 552 311440 564
rect 311492 552 311498 604
rect 312630 592 312636 604
rect 312591 564 312636 592
rect 312630 552 312636 564
rect 312688 552 312694 604
rect 314626 592 314654 632
rect 315132 632 318524 660
rect 315132 592 315160 632
rect 318518 620 318524 632
rect 318576 620 318582 672
rect 318702 620 318708 672
rect 318760 620 318766 672
rect 319530 620 319536 672
rect 319588 660 319594 672
rect 319588 632 326752 660
rect 319588 620 319594 632
rect 314626 564 315160 592
rect 315942 552 315948 604
rect 316000 592 316006 604
rect 316000 564 316172 592
rect 316000 552 316006 564
rect 309060 524 309088 552
rect 303540 496 309088 524
rect 295668 484 295674 496
rect 280890 456 280896 468
rect 280126 428 280896 456
rect 279605 419 279663 425
rect 280890 416 280896 428
rect 280948 416 280954 468
rect 284110 416 284116 468
rect 284168 456 284174 468
rect 291194 456 291200 468
rect 284168 428 291200 456
rect 284168 416 284174 428
rect 291194 416 291200 428
rect 291252 416 291258 468
rect 300210 416 300216 468
rect 300268 456 300274 468
rect 307941 459 307999 465
rect 307941 456 307953 459
rect 300268 428 307953 456
rect 300268 416 300274 428
rect 307941 425 307953 428
rect 307987 425 307999 459
rect 307941 419 307999 425
rect 246816 360 252416 388
rect 258046 388 258074 416
rect 263134 388 263140 400
rect 258046 360 263140 388
rect 246816 348 246822 360
rect 263134 348 263140 360
rect 263192 348 263198 400
rect 269482 348 269488 400
rect 269540 388 269546 400
rect 276198 388 276204 400
rect 269540 360 276204 388
rect 269540 348 269546 360
rect 276198 348 276204 360
rect 276256 348 276262 400
rect 278590 348 278596 400
rect 278648 388 278654 400
rect 279697 391 279755 397
rect 279697 388 279709 391
rect 278648 360 279709 388
rect 278648 348 278654 360
rect 279697 357 279709 360
rect 279743 357 279755 391
rect 279697 351 279755 357
rect 294506 348 294512 400
rect 294564 388 294570 400
rect 301774 388 301780 400
rect 294564 360 301780 388
rect 294564 348 294570 360
rect 301774 348 301780 360
rect 301832 348 301838 400
rect 302418 348 302424 400
rect 302476 388 302482 400
rect 310256 388 310284 552
rect 311161 527 311219 533
rect 311161 493 311173 527
rect 311207 524 311219 527
rect 316034 524 316040 536
rect 311207 496 316040 524
rect 311207 493 311219 496
rect 311161 487 311219 493
rect 316034 484 316040 496
rect 316092 484 316098 536
rect 316144 524 316172 564
rect 317138 552 317144 604
rect 317196 592 317202 604
rect 325602 592 325608 604
rect 317196 564 325608 592
rect 317196 552 317202 564
rect 325602 552 325608 564
rect 325660 552 325666 604
rect 326724 592 326752 632
rect 326798 620 326804 672
rect 326856 620 326862 672
rect 328454 620 328460 672
rect 328512 620 328518 672
rect 331950 620 331956 672
rect 332008 660 332014 672
rect 332008 632 333974 660
rect 332008 620 332014 632
rect 327994 592 328000 604
rect 326724 564 328000 592
rect 327994 552 328000 564
rect 328052 552 328058 604
rect 330386 552 330392 604
rect 330444 552 330450 604
rect 316144 496 320220 524
rect 316586 456 316592 468
rect 302476 360 310284 388
rect 310992 428 316592 456
rect 302476 348 302482 360
rect 242250 280 242256 332
rect 242308 320 242314 332
rect 247310 320 247316 332
rect 242308 292 247316 320
rect 242308 280 242314 292
rect 247310 280 247316 292
rect 247368 280 247374 332
rect 250898 280 250904 332
rect 250956 320 250962 332
rect 255501 323 255559 329
rect 255501 320 255513 323
rect 250956 292 255513 320
rect 250956 280 250962 292
rect 255501 289 255513 292
rect 255547 289 255559 323
rect 255501 283 255559 289
rect 256878 280 256884 332
rect 256936 320 256942 332
rect 262766 320 262772 332
rect 256936 292 262772 320
rect 256936 280 256942 292
rect 262766 280 262772 292
rect 262824 280 262830 332
rect 271782 280 271788 332
rect 271840 320 271846 332
rect 278498 320 278504 332
rect 271840 292 278504 320
rect 271840 280 271846 292
rect 278498 280 278504 292
rect 278556 280 278562 332
rect 297910 280 297916 332
rect 297968 320 297974 332
rect 305730 320 305736 332
rect 297968 292 305736 320
rect 297968 280 297974 292
rect 305730 280 305736 292
rect 305788 280 305794 332
rect 308766 280 308772 332
rect 308824 320 308830 332
rect 310992 320 311020 428
rect 316586 416 316592 428
rect 316644 416 316650 468
rect 318334 416 318340 468
rect 318392 456 318398 468
rect 318702 456 318708 468
rect 318392 428 318708 456
rect 318392 416 318398 428
rect 318702 416 318708 428
rect 318760 416 318766 468
rect 320192 456 320220 496
rect 321554 484 321560 536
rect 321612 524 321618 536
rect 330404 524 330432 552
rect 321612 496 330432 524
rect 333946 524 333974 632
rect 337470 620 337476 672
rect 337528 620 337534 672
rect 342162 660 342168 672
rect 338500 632 342168 660
rect 334805 595 334863 601
rect 334805 561 334817 595
rect 334851 592 334863 595
rect 338500 592 338528 632
rect 342162 620 342168 632
rect 342220 620 342226 672
rect 344986 660 345014 700
rect 342824 632 345014 660
rect 338666 592 338672 604
rect 334851 564 338528 592
rect 338627 564 338672 592
rect 334851 561 334863 564
rect 334805 555 334863 561
rect 338666 552 338672 564
rect 338724 552 338730 604
rect 338761 595 338819 601
rect 338761 561 338773 595
rect 338807 592 338819 595
rect 339862 592 339868 604
rect 338807 564 339868 592
rect 338807 561 338819 564
rect 338761 555 338819 561
rect 339862 552 339868 564
rect 339920 552 339926 604
rect 340966 552 340972 604
rect 341024 552 341030 604
rect 342070 552 342076 604
rect 342128 592 342134 604
rect 342128 564 342254 592
rect 342128 552 342134 564
rect 340984 524 341012 552
rect 333946 496 341012 524
rect 342226 524 342254 564
rect 342824 524 342852 632
rect 348234 620 348240 672
rect 348292 660 348298 672
rect 349062 660 349068 672
rect 348292 632 349068 660
rect 348292 620 348298 632
rect 349062 620 349068 632
rect 349120 620 349126 672
rect 350460 660 350488 700
rect 356026 700 358814 728
rect 351638 660 351644 672
rect 350460 632 351644 660
rect 351638 620 351644 632
rect 351696 620 351702 672
rect 352466 620 352472 672
rect 352524 660 352530 672
rect 356026 660 356054 700
rect 352524 632 356054 660
rect 358786 660 358814 700
rect 370700 672 370728 768
rect 377232 768 382274 796
rect 372586 700 375512 728
rect 361942 660 361948 672
rect 358786 632 361948 660
rect 352524 620 352530 632
rect 361942 620 361948 632
rect 362000 620 362006 672
rect 362313 663 362371 669
rect 362313 629 362325 663
rect 362359 660 362371 663
rect 369578 660 369584 672
rect 362359 632 369584 660
rect 362359 629 362371 632
rect 362313 623 362371 629
rect 369578 620 369584 632
rect 369636 620 369642 672
rect 370406 660 370412 672
rect 370367 632 370412 660
rect 370406 620 370412 632
rect 370464 620 370470 672
rect 370682 620 370688 672
rect 370740 620 370746 672
rect 371602 620 371608 672
rect 371660 660 371666 672
rect 372586 660 372614 700
rect 375190 660 375196 672
rect 371660 632 372614 660
rect 375151 632 375196 660
rect 371660 620 371666 632
rect 375190 620 375196 632
rect 375248 620 375254 672
rect 375484 660 375512 700
rect 377232 660 377260 768
rect 382246 728 382274 768
rect 382246 700 382412 728
rect 382384 672 382412 700
rect 385972 672 386000 836
rect 393317 833 393329 867
rect 393363 864 393375 867
rect 404556 864 404584 904
rect 404817 901 404829 904
rect 404863 901 404875 935
rect 404817 895 404875 901
rect 408466 864 408494 972
rect 415489 969 415501 972
rect 415535 969 415547 1003
rect 415489 963 415547 969
rect 418341 1003 418399 1009
rect 418341 969 418353 1003
rect 418387 1000 418399 1003
rect 425701 1003 425759 1009
rect 425701 1000 425713 1003
rect 418387 972 425713 1000
rect 418387 969 418399 972
rect 418341 963 418399 969
rect 425701 969 425713 972
rect 425747 969 425759 1003
rect 435913 1003 435971 1009
rect 435913 1000 435925 1003
rect 425701 963 425759 969
rect 430546 972 435925 1000
rect 409233 935 409291 941
rect 409233 901 409245 935
rect 409279 932 409291 935
rect 421009 935 421067 941
rect 421009 932 421021 935
rect 409279 904 421021 932
rect 409279 901 409291 904
rect 409233 895 409291 901
rect 421009 901 421021 904
rect 421055 901 421067 935
rect 430546 932 430574 972
rect 435913 969 435925 972
rect 435959 969 435971 1003
rect 435913 963 435971 969
rect 436465 1003 436523 1009
rect 436465 969 436477 1003
rect 436511 1000 436523 1003
rect 454221 1003 454279 1009
rect 436511 972 440464 1000
rect 436511 969 436523 972
rect 436465 963 436523 969
rect 438673 935 438731 941
rect 438673 932 438685 935
rect 421009 895 421067 901
rect 425026 904 430574 932
rect 437446 904 438685 932
rect 393363 836 404584 864
rect 404648 836 408494 864
rect 412637 867 412695 873
rect 393363 833 393375 836
rect 393317 827 393375 833
rect 400186 768 401594 796
rect 400186 728 400214 768
rect 396644 700 400214 728
rect 401566 728 401594 768
rect 404648 728 404676 836
rect 412637 833 412649 867
rect 412683 864 412695 867
rect 412683 836 420914 864
rect 412683 833 412695 836
rect 412637 827 412695 833
rect 404725 799 404783 805
rect 404725 765 404737 799
rect 404771 796 404783 799
rect 404771 768 416728 796
rect 404771 765 404783 768
rect 404725 759 404783 765
rect 401566 700 402560 728
rect 375484 632 377260 660
rect 377398 620 377404 672
rect 377456 660 377462 672
rect 377456 632 382274 660
rect 377456 620 377462 632
rect 344462 552 344468 604
rect 344520 592 344526 604
rect 354030 592 354036 604
rect 344520 564 354036 592
rect 344520 552 344526 564
rect 354030 552 354036 564
rect 354088 552 354094 604
rect 356330 592 356336 604
rect 354600 564 356336 592
rect 342226 496 342852 524
rect 321612 484 321618 496
rect 343174 484 343180 536
rect 343232 524 343238 536
rect 351822 524 351828 536
rect 343232 496 351828 524
rect 343232 484 343238 496
rect 351822 484 351828 496
rect 351880 484 351886 536
rect 324222 456 324228 468
rect 320192 428 324228 456
rect 324222 416 324228 428
rect 324280 416 324286 468
rect 325142 416 325148 468
rect 325200 456 325206 468
rect 333606 456 333612 468
rect 325200 428 333612 456
rect 325200 416 325206 428
rect 333606 416 333612 428
rect 333664 416 333670 468
rect 346762 416 346768 468
rect 346820 456 346826 468
rect 354600 456 354628 564
rect 356330 552 356336 564
rect 356388 552 356394 604
rect 358722 592 358728 604
rect 358683 564 358728 592
rect 358722 552 358728 564
rect 358780 552 358786 604
rect 364794 592 364800 604
rect 359108 564 364800 592
rect 354674 484 354680 536
rect 354732 524 354738 536
rect 359108 524 359136 564
rect 364794 552 364800 564
rect 364852 552 364858 604
rect 364889 595 364947 601
rect 364889 561 364901 595
rect 364935 592 364947 595
rect 368198 592 368204 604
rect 364935 564 368204 592
rect 364935 561 364947 564
rect 364889 555 364947 561
rect 368198 552 368204 564
rect 368256 552 368262 604
rect 369302 552 369308 604
rect 369360 592 369366 604
rect 379974 592 379980 604
rect 369360 564 379980 592
rect 369360 552 369366 564
rect 379974 552 379980 564
rect 380032 552 380038 604
rect 381170 552 381176 604
rect 381228 552 381234 604
rect 382246 592 382274 632
rect 382366 620 382372 672
rect 382424 620 382430 672
rect 385954 620 385960 672
rect 386012 620 386018 672
rect 388806 660 388812 672
rect 388767 632 388812 660
rect 388806 620 388812 632
rect 388864 620 388870 672
rect 396534 660 396540 672
rect 389468 632 396540 660
rect 388254 592 388260 604
rect 382246 564 388260 592
rect 388254 552 388260 564
rect 388312 552 388318 604
rect 354732 496 359136 524
rect 354732 484 354738 496
rect 359274 484 359280 536
rect 359332 524 359338 536
rect 362313 527 362371 533
rect 362313 524 362325 527
rect 359332 496 362325 524
rect 359332 484 359338 496
rect 362313 493 362325 496
rect 362359 493 362371 527
rect 362313 487 362371 493
rect 362678 484 362684 536
rect 362736 524 362742 536
rect 373074 524 373080 536
rect 362736 496 373080 524
rect 362736 484 362742 496
rect 373074 484 373080 496
rect 373132 484 373138 536
rect 377398 524 377404 536
rect 373184 496 377404 524
rect 346820 428 354628 456
rect 346820 416 346826 428
rect 356974 416 356980 468
rect 357032 456 357038 468
rect 357032 428 359136 456
rect 357032 416 357038 428
rect 311066 348 311072 400
rect 311124 388 311130 400
rect 319898 388 319904 400
rect 311124 360 319904 388
rect 311124 348 311130 360
rect 319898 348 319904 360
rect 319956 348 319962 400
rect 327442 348 327448 400
rect 327500 388 327506 400
rect 336458 388 336464 400
rect 327500 360 336464 388
rect 327500 348 327506 360
rect 336458 348 336464 360
rect 336516 348 336522 400
rect 349062 348 349068 400
rect 349120 388 349126 400
rect 358725 391 358783 397
rect 358725 388 358737 391
rect 349120 360 358737 388
rect 349120 348 349126 360
rect 358725 357 358737 360
rect 358771 357 358783 391
rect 359108 388 359136 428
rect 360378 416 360384 468
rect 360436 456 360442 468
rect 364705 459 364763 465
rect 364705 456 364717 459
rect 360436 428 364717 456
rect 360436 416 360442 428
rect 364705 425 364717 428
rect 364751 425 364763 459
rect 364705 419 364763 425
rect 366726 416 366732 468
rect 366784 456 366790 468
rect 373184 456 373212 496
rect 377398 484 377404 496
rect 377456 484 377462 536
rect 377493 527 377551 533
rect 377493 493 377505 527
rect 377539 524 377551 527
rect 381188 524 381216 552
rect 377539 496 381216 524
rect 377539 493 377551 496
rect 377493 487 377551 493
rect 385402 484 385408 536
rect 385460 524 385466 536
rect 389468 524 389496 632
rect 396534 620 396540 632
rect 396592 620 396598 672
rect 391014 552 391020 604
rect 391072 592 391078 604
rect 394145 595 394203 601
rect 394145 592 394157 595
rect 391072 564 394157 592
rect 391072 552 391078 564
rect 394145 561 394157 564
rect 394191 561 394203 595
rect 394145 555 394203 561
rect 394329 595 394387 601
rect 394329 561 394341 595
rect 394375 592 394387 595
rect 396644 592 396672 700
rect 402532 672 402560 700
rect 403452 700 404676 728
rect 408466 700 410840 728
rect 403452 672 403480 700
rect 400030 660 400036 672
rect 399991 632 400036 660
rect 400030 620 400036 632
rect 400088 620 400094 672
rect 402514 620 402520 672
rect 402572 620 402578 672
rect 403434 620 403440 672
rect 403492 620 403498 672
rect 408466 660 408494 700
rect 410812 672 410840 700
rect 416700 672 416728 768
rect 420886 728 420914 836
rect 420886 700 421144 728
rect 421116 672 421144 700
rect 409230 660 409236 672
rect 403636 632 408494 660
rect 409191 632 409236 660
rect 397730 592 397736 604
rect 394375 564 396672 592
rect 397691 564 397736 592
rect 394375 561 394387 564
rect 394329 555 394387 561
rect 397730 552 397736 564
rect 397788 552 397794 604
rect 398834 552 398840 604
rect 398892 552 398898 604
rect 400214 592 400220 604
rect 400175 564 400220 592
rect 400214 552 400220 564
rect 400272 552 400278 604
rect 400306 552 400312 604
rect 400364 592 400370 604
rect 403526 592 403532 604
rect 400364 564 403532 592
rect 400364 552 400370 564
rect 403526 552 403532 564
rect 403584 552 403590 604
rect 385460 496 389496 524
rect 385460 484 385466 496
rect 389818 484 389824 536
rect 389876 524 389882 536
rect 394053 527 394111 533
rect 394053 524 394065 527
rect 389876 496 394065 524
rect 389876 484 389882 496
rect 394053 493 394065 496
rect 394099 493 394111 527
rect 398852 524 398880 552
rect 403636 524 403664 632
rect 409230 620 409236 632
rect 409288 620 409294 672
rect 410794 620 410800 672
rect 410852 620 410858 672
rect 411226 632 416636 660
rect 404722 592 404728 604
rect 404683 564 404728 592
rect 404722 552 404728 564
rect 404780 552 404786 604
rect 404814 552 404820 604
rect 404872 592 404878 604
rect 404872 564 404917 592
rect 404872 552 404878 564
rect 405642 552 405648 604
rect 405700 592 405706 604
rect 411226 592 411254 632
rect 412634 592 412640 604
rect 405700 564 411254 592
rect 412595 564 412640 592
rect 405700 552 405706 564
rect 412634 552 412640 564
rect 412692 552 412698 604
rect 413738 592 413744 604
rect 413699 564 413744 592
rect 413738 552 413744 564
rect 413796 552 413802 604
rect 414290 592 414296 604
rect 414251 564 414296 592
rect 414290 552 414296 564
rect 414348 552 414354 604
rect 415486 592 415492 604
rect 415447 564 415492 592
rect 415486 552 415492 564
rect 415544 552 415550 604
rect 416608 592 416636 632
rect 416682 620 416688 672
rect 416740 620 416746 672
rect 418338 660 418344 672
rect 418299 632 418344 660
rect 418338 620 418344 632
rect 418396 620 418402 672
rect 421006 660 421012 672
rect 420967 632 421012 660
rect 421006 620 421012 632
rect 421064 620 421070 672
rect 421098 620 421104 672
rect 421156 620 421162 672
rect 423490 620 423496 672
rect 423548 660 423554 672
rect 425026 660 425054 904
rect 437446 796 437474 904
rect 438673 901 438685 904
rect 438719 901 438731 935
rect 438673 895 438731 901
rect 425624 768 437474 796
rect 438504 836 440234 864
rect 425624 672 425652 768
rect 428369 731 428427 737
rect 428369 697 428381 731
rect 428415 728 428427 731
rect 435913 731 435971 737
rect 428415 700 435680 728
rect 428415 697 428427 700
rect 428369 691 428427 697
rect 425514 660 425520 672
rect 423548 632 425054 660
rect 425475 632 425520 660
rect 423548 620 423554 632
rect 425514 620 425520 632
rect 425572 620 425578 672
rect 425606 620 425612 672
rect 425664 620 425670 672
rect 425701 663 425759 669
rect 425701 629 425713 663
rect 425747 660 425759 663
rect 430850 660 430856 672
rect 425747 632 430856 660
rect 425747 629 425759 632
rect 425701 623 425759 629
rect 430850 620 430856 632
rect 430908 620 430914 672
rect 431862 660 431868 672
rect 431823 632 431868 660
rect 431862 620 431868 632
rect 431920 620 431926 672
rect 432046 660 432052 672
rect 432007 632 432052 660
rect 432046 620 432052 632
rect 432104 620 432110 672
rect 434165 663 434223 669
rect 434165 660 434177 663
rect 433168 632 434177 660
rect 417878 592 417884 604
rect 416608 564 417884 592
rect 417878 552 417884 564
rect 417936 552 417942 604
rect 420917 595 420975 601
rect 420917 561 420929 595
rect 420963 592 420975 595
rect 423766 592 423772 604
rect 420963 564 423772 592
rect 420963 561 420975 564
rect 420917 555 420975 561
rect 423766 552 423772 564
rect 423824 552 423830 604
rect 423861 595 423919 601
rect 423861 561 423873 595
rect 423907 592 423919 595
rect 427262 592 427268 604
rect 423907 564 427268 592
rect 423907 561 423919 564
rect 423861 555 423919 561
rect 427262 552 427268 564
rect 427320 552 427326 604
rect 428366 592 428372 604
rect 428327 564 428372 592
rect 428366 552 428372 564
rect 428424 552 428430 604
rect 429470 552 429476 604
rect 429528 592 429534 604
rect 433168 592 433196 632
rect 434165 629 434177 632
rect 434211 629 434223 663
rect 434165 623 434223 629
rect 429528 564 433196 592
rect 429528 552 429534 564
rect 433242 552 433248 604
rect 433300 552 433306 604
rect 434714 552 434720 604
rect 434772 592 434778 604
rect 435542 592 435548 604
rect 434772 564 435548 592
rect 434772 552 434778 564
rect 435542 552 435548 564
rect 435600 552 435606 604
rect 435652 592 435680 700
rect 435913 697 435925 731
rect 435959 728 435971 731
rect 435959 700 436784 728
rect 435959 697 435971 700
rect 435913 691 435971 697
rect 436756 672 436784 700
rect 436462 660 436468 672
rect 436423 632 436468 660
rect 436462 620 436468 632
rect 436520 620 436526 672
rect 436738 620 436744 672
rect 436796 620 436802 672
rect 437474 620 437480 672
rect 437532 660 437538 672
rect 438504 660 438532 836
rect 439866 660 439872 672
rect 437532 632 438532 660
rect 438596 632 439728 660
rect 439827 632 439872 660
rect 437532 620 437538 632
rect 438596 592 438624 632
rect 435652 564 438624 592
rect 438673 595 438731 601
rect 438673 561 438685 595
rect 438719 592 438731 595
rect 439130 592 439136 604
rect 438719 564 439136 592
rect 438719 561 438731 564
rect 438673 555 438731 561
rect 439130 552 439136 564
rect 439188 552 439194 604
rect 439700 592 439728 632
rect 439866 620 439872 632
rect 439924 620 439930 672
rect 440206 660 440234 836
rect 440436 728 440464 972
rect 454221 969 454233 1003
rect 454267 1000 454279 1003
rect 465629 1003 465687 1009
rect 454267 972 465488 1000
rect 454267 969 454279 972
rect 454221 963 454279 969
rect 444469 935 444527 941
rect 444469 901 444481 935
rect 444515 932 444527 935
rect 458085 935 458143 941
rect 458085 932 458097 935
rect 444515 904 458097 932
rect 444515 901 444527 904
rect 444469 895 444527 901
rect 458085 901 458097 904
rect 458131 901 458143 935
rect 458085 895 458143 901
rect 452289 867 452347 873
rect 452289 864 452301 867
rect 442966 836 452301 864
rect 440513 799 440571 805
rect 440513 765 440525 799
rect 440559 796 440571 799
rect 442966 796 442994 836
rect 452289 833 452301 836
rect 452335 833 452347 867
rect 452289 827 452347 833
rect 440559 768 442994 796
rect 446677 799 446735 805
rect 440559 765 440571 768
rect 440513 759 440571 765
rect 446677 765 446689 799
rect 446723 796 446735 799
rect 456061 799 456119 805
rect 446723 768 454034 796
rect 446723 765 446735 768
rect 446677 759 446735 765
rect 454006 728 454034 768
rect 456061 765 456073 799
rect 456107 796 456119 799
rect 456107 768 460704 796
rect 456107 765 456119 768
rect 456061 759 456119 765
rect 440436 700 450032 728
rect 454006 700 460428 728
rect 450004 672 450032 700
rect 460400 672 460428 700
rect 460676 672 460704 768
rect 465460 728 465488 972
rect 465629 969 465641 1003
rect 465675 1000 465687 1003
rect 474553 1003 474611 1009
rect 474553 1000 474565 1003
rect 465675 972 474565 1000
rect 465675 969 465687 972
rect 465629 963 465687 969
rect 474553 969 474565 972
rect 474599 969 474611 1003
rect 474553 963 474611 969
rect 488261 1003 488319 1009
rect 488261 969 488273 1003
rect 488307 1000 488319 1003
rect 503993 1003 504051 1009
rect 503993 1000 504005 1003
rect 488307 972 504005 1000
rect 488307 969 488319 972
rect 488261 963 488319 969
rect 503993 969 504005 972
rect 504039 969 504051 1003
rect 503993 963 504051 969
rect 505741 1003 505799 1009
rect 505741 969 505753 1003
rect 505787 1000 505799 1003
rect 521933 1003 521991 1009
rect 521933 1000 521945 1003
rect 505787 972 521945 1000
rect 505787 969 505799 972
rect 505741 963 505799 969
rect 521933 969 521945 972
rect 521979 969 521991 1003
rect 539781 1003 539839 1009
rect 539781 1000 539793 1003
rect 521933 963 521991 969
rect 523420 972 539793 1000
rect 470597 935 470655 941
rect 470597 901 470609 935
rect 470643 932 470655 935
rect 485225 935 485283 941
rect 485225 932 485237 935
rect 470643 904 485237 932
rect 470643 901 470655 904
rect 470597 895 470655 901
rect 485225 901 485237 904
rect 485271 901 485283 935
rect 485225 895 485283 901
rect 485317 935 485375 941
rect 485317 901 485329 935
rect 485363 932 485375 935
rect 496817 935 496875 941
rect 496817 932 496829 935
rect 485363 904 496829 932
rect 485363 901 485375 904
rect 485317 895 485375 901
rect 496817 901 496829 904
rect 496863 901 496875 935
rect 496817 895 496875 901
rect 498933 935 498991 941
rect 498933 901 498945 935
rect 498979 932 498991 935
rect 514941 935 514999 941
rect 514941 932 514953 935
rect 498979 904 514953 932
rect 498979 901 498991 904
rect 498933 895 498991 901
rect 514941 901 514953 904
rect 514987 901 514999 935
rect 514941 895 514999 901
rect 518161 935 518219 941
rect 518161 901 518173 935
rect 518207 932 518219 935
rect 518345 935 518403 941
rect 518345 932 518357 935
rect 518207 904 518357 932
rect 518207 901 518219 904
rect 518161 895 518219 901
rect 518345 901 518357 904
rect 518391 901 518403 935
rect 518345 895 518403 901
rect 486605 867 486663 873
rect 486605 864 486617 867
rect 482986 836 486617 864
rect 471701 799 471759 805
rect 471701 765 471713 799
rect 471747 796 471759 799
rect 482986 796 483014 836
rect 486605 833 486617 836
rect 486651 833 486663 867
rect 509881 867 509939 873
rect 486605 827 486663 833
rect 492646 836 498240 864
rect 492646 796 492674 836
rect 471747 768 483014 796
rect 485056 768 492674 796
rect 471747 765 471759 768
rect 471701 759 471759 765
rect 485056 728 485084 768
rect 465460 700 468708 728
rect 468680 672 468708 700
rect 482940 700 485084 728
rect 485133 731 485191 737
rect 482940 672 482968 700
rect 485133 697 485145 731
rect 485179 728 485191 731
rect 485179 700 489914 728
rect 485179 697 485191 700
rect 485133 691 485191 697
rect 449897 663 449955 669
rect 449897 660 449909 663
rect 440206 632 449909 660
rect 449897 629 449909 632
rect 449943 629 449955 663
rect 449897 623 449955 629
rect 449986 620 449992 672
rect 450044 620 450050 672
rect 453574 660 453580 672
rect 453535 632 453580 660
rect 453574 620 453580 632
rect 453632 620 453638 672
rect 454218 660 454224 672
rect 454179 632 454224 660
rect 454218 620 454224 632
rect 454276 620 454282 672
rect 454494 660 454500 672
rect 454455 632 454500 660
rect 454494 620 454500 632
rect 454552 620 454558 672
rect 454773 663 454831 669
rect 454773 629 454785 663
rect 454819 660 454831 663
rect 456886 660 456892 672
rect 454819 632 456892 660
rect 454819 629 454831 632
rect 454773 623 454831 629
rect 456886 620 456892 632
rect 456944 620 456950 672
rect 460382 620 460388 672
rect 460440 620 460446 672
rect 460658 620 460664 672
rect 460716 620 460722 672
rect 462130 660 462136 672
rect 462091 632 462136 660
rect 462130 620 462136 632
rect 462188 620 462194 672
rect 466362 660 466368 672
rect 466323 632 466368 660
rect 466362 620 466368 632
rect 466420 620 466426 672
rect 467190 660 467196 672
rect 467151 632 467196 660
rect 467190 620 467196 632
rect 467248 620 467254 672
rect 468294 660 468300 672
rect 468255 632 468300 660
rect 468294 620 468300 632
rect 468352 620 468358 672
rect 468662 620 468668 672
rect 468720 620 468726 672
rect 477862 660 477868 672
rect 469186 632 477868 660
rect 441522 592 441528 604
rect 439700 564 441528 592
rect 441522 552 441528 564
rect 441580 552 441586 604
rect 442626 592 442632 604
rect 442587 564 442632 592
rect 442626 552 442632 564
rect 442684 552 442690 604
rect 444466 592 444472 604
rect 444427 564 444472 592
rect 444466 552 444472 564
rect 444524 552 444530 604
rect 445018 592 445024 604
rect 444979 564 445024 592
rect 445018 552 445024 564
rect 445076 552 445082 604
rect 446214 592 446220 604
rect 445726 564 446220 592
rect 408218 524 408224 536
rect 398852 496 403664 524
rect 403728 496 408224 524
rect 394053 487 394111 493
rect 366784 428 373212 456
rect 366784 416 366790 428
rect 373902 416 373908 468
rect 373960 456 373966 468
rect 384574 456 384580 468
rect 373960 428 384580 456
rect 373960 416 373966 428
rect 384574 416 384580 428
rect 384632 416 384638 468
rect 393314 456 393320 468
rect 393275 428 393320 456
rect 393314 416 393320 428
rect 393372 416 393378 468
rect 395614 416 395620 468
rect 395672 456 395678 468
rect 399849 459 399907 465
rect 399849 456 399861 459
rect 395672 428 399861 456
rect 395672 416 395678 428
rect 399849 425 399861 428
rect 399895 425 399907 459
rect 399849 419 399907 425
rect 402149 459 402207 465
rect 402149 425 402161 459
rect 402195 456 402207 459
rect 403728 456 403756 496
rect 408218 484 408224 496
rect 408276 484 408282 536
rect 410334 484 410340 536
rect 410392 524 410398 536
rect 422754 524 422760 536
rect 410392 496 422760 524
rect 410392 484 410398 496
rect 422754 484 422760 496
rect 422812 484 422818 536
rect 433260 524 433288 552
rect 430546 496 433288 524
rect 402195 428 403756 456
rect 403805 459 403863 465
rect 402195 425 402207 428
rect 402149 419 402207 425
rect 403805 425 403817 459
rect 403851 456 403863 459
rect 405734 456 405740 468
rect 403851 428 405740 456
rect 403851 425 403863 428
rect 403805 419 403863 425
rect 405734 416 405740 428
rect 405792 416 405798 468
rect 408126 416 408132 468
rect 408184 456 408190 468
rect 419902 456 419908 468
rect 408184 428 419908 456
rect 408184 416 408190 428
rect 419902 416 419908 428
rect 419960 416 419966 468
rect 420546 416 420552 468
rect 420604 456 420610 468
rect 430546 456 430574 496
rect 438762 484 438768 536
rect 438820 524 438826 536
rect 440513 527 440571 533
rect 440513 524 440525 527
rect 438820 496 440525 524
rect 438820 484 438826 496
rect 440513 493 440525 496
rect 440559 493 440571 527
rect 440513 487 440571 493
rect 420604 428 430574 456
rect 420604 416 420610 428
rect 430666 416 430672 468
rect 430724 456 430730 468
rect 430724 428 433012 456
rect 430724 416 430730 428
rect 367278 388 367284 400
rect 359108 360 367284 388
rect 358725 351 358783 357
rect 367278 348 367284 360
rect 367336 348 367342 400
rect 372430 348 372436 400
rect 372488 388 372494 400
rect 372488 360 376616 388
rect 372488 348 372494 360
rect 308824 292 311020 320
rect 308824 280 308830 292
rect 312446 280 312452 332
rect 312504 320 312510 332
rect 320726 320 320732 332
rect 312504 292 320732 320
rect 312504 280 312510 292
rect 320726 280 320732 292
rect 320784 280 320790 332
rect 333146 280 333152 332
rect 333204 320 333210 332
rect 334805 323 334863 329
rect 334805 320 334817 323
rect 333204 292 334817 320
rect 333204 280 333210 292
rect 334805 289 334817 292
rect 334851 289 334863 323
rect 334805 283 334863 289
rect 340598 280 340604 332
rect 340656 320 340662 332
rect 347774 320 347780 332
rect 340656 292 347780 320
rect 340656 280 340662 292
rect 347774 280 347780 292
rect 347832 280 347838 332
rect 351270 280 351276 332
rect 351328 320 351334 332
rect 360838 320 360844 332
rect 351328 292 360844 320
rect 351328 280 351334 292
rect 360838 280 360844 292
rect 360896 280 360902 332
rect 363782 280 363788 332
rect 363840 320 363846 332
rect 374270 320 374276 332
rect 363840 292 374276 320
rect 363840 280 363846 292
rect 374270 280 374276 292
rect 374328 280 374334 332
rect 376588 320 376616 360
rect 378594 348 378600 400
rect 378652 388 378658 400
rect 389174 388 389180 400
rect 378652 360 389180 388
rect 378652 348 378658 360
rect 389174 348 389180 360
rect 389232 348 389238 400
rect 389910 348 389916 400
rect 389968 388 389974 400
rect 393774 388 393780 400
rect 389968 360 393780 388
rect 389968 348 389974 360
rect 393774 348 393780 360
rect 393832 348 393838 400
rect 396046 360 398604 388
rect 383286 320 383292 332
rect 376588 292 383292 320
rect 383286 280 383292 292
rect 383344 280 383350 332
rect 386966 280 386972 332
rect 387024 320 387030 332
rect 394418 320 394424 332
rect 387024 292 394424 320
rect 387024 280 387030 292
rect 394418 280 394424 292
rect 394476 280 394482 332
rect 233234 212 233240 264
rect 233292 212 233298 264
rect 236546 212 236552 264
rect 236604 252 236610 264
rect 241422 252 241428 264
rect 236604 224 241428 252
rect 236604 212 236610 224
rect 241422 212 241428 224
rect 241480 212 241486 264
rect 255682 212 255688 264
rect 255740 252 255746 264
rect 261478 252 261484 264
rect 255740 224 261484 252
rect 255740 212 255746 224
rect 261478 212 261484 224
rect 261536 212 261542 264
rect 261570 212 261576 264
rect 261628 252 261634 264
rect 267550 252 267556 264
rect 261628 224 267556 252
rect 261628 212 261634 224
rect 267550 212 267556 224
rect 267608 212 267614 264
rect 280430 212 280436 264
rect 280488 252 280494 264
rect 287054 252 287060 264
rect 280488 224 287060 252
rect 280488 212 280494 224
rect 287054 212 287060 224
rect 287112 212 287118 264
rect 296806 212 296812 264
rect 296864 252 296870 264
rect 303982 252 303988 264
rect 296864 224 303988 252
rect 296864 212 296870 224
rect 303982 212 303988 224
rect 304040 212 304046 264
rect 307662 212 307668 264
rect 307720 252 307726 264
rect 311161 255 311219 261
rect 311161 252 311173 255
rect 307720 224 311173 252
rect 307720 212 307726 224
rect 311161 221 311173 224
rect 311207 221 311219 255
rect 311161 215 311219 221
rect 313642 212 313648 264
rect 313700 252 313706 264
rect 321830 252 321836 264
rect 313700 224 321836 252
rect 313700 212 313706 224
rect 321830 212 321836 224
rect 321888 212 321894 264
rect 322842 212 322848 264
rect 322900 252 322906 264
rect 331214 252 331220 264
rect 322900 224 331220 252
rect 322900 212 322906 224
rect 331214 212 331220 224
rect 331272 212 331278 264
rect 337194 212 337200 264
rect 337252 252 337258 264
rect 337252 224 342254 252
rect 337252 212 337258 224
rect 186958 184 186964 196
rect 184906 156 186964 184
rect 16298 76 16304 128
rect 16356 116 16362 128
rect 18966 116 18972 128
rect 16356 88 18972 116
rect 16356 76 16362 88
rect 18966 76 18972 88
rect 19024 76 19030 128
rect 45738 76 45744 128
rect 45796 116 45802 128
rect 47394 116 47400 128
rect 45796 88 47400 116
rect 45796 76 45802 88
rect 47394 76 47400 88
rect 47452 76 47458 128
rect 129826 76 129832 128
rect 129884 116 129890 128
rect 130286 116 130292 128
rect 129884 88 130292 116
rect 129884 76 129890 88
rect 130286 76 130292 88
rect 130344 76 130350 128
rect 155954 76 155960 128
rect 156012 116 156018 128
rect 157518 116 157524 128
rect 156012 88 157524 116
rect 156012 76 156018 88
rect 157518 76 157524 88
rect 157576 76 157582 128
rect 159358 76 159364 128
rect 159416 116 159422 128
rect 161474 116 161480 128
rect 159416 88 161480 116
rect 159416 76 159422 88
rect 161474 76 161480 88
rect 161532 76 161538 128
rect 184290 76 184296 128
rect 184348 116 184354 128
rect 184906 116 184934 156
rect 186958 144 186964 156
rect 187016 144 187022 196
rect 228542 144 228548 196
rect 228600 184 228606 196
rect 233252 184 233280 212
rect 228600 156 233280 184
rect 228600 144 228606 156
rect 264882 144 264888 196
rect 264940 184 264946 196
rect 271046 184 271052 196
rect 264940 156 271052 184
rect 264940 144 264946 156
rect 271046 144 271052 156
rect 271104 144 271110 196
rect 282914 144 282920 196
rect 282972 184 282978 196
rect 289998 184 290004 196
rect 282972 156 290004 184
rect 282972 144 282978 156
rect 289998 144 290004 156
rect 290056 144 290062 196
rect 292206 144 292212 196
rect 292264 184 292270 196
rect 299382 184 299388 196
rect 292264 156 299388 184
rect 292264 144 292270 156
rect 299382 144 299388 156
rect 299440 144 299446 196
rect 324038 144 324044 196
rect 324096 184 324102 196
rect 332502 184 332508 196
rect 324096 156 332508 184
rect 324096 144 324102 156
rect 332502 144 332508 156
rect 332560 144 332566 196
rect 338298 144 338304 196
rect 338356 184 338362 196
rect 342226 184 342254 224
rect 345566 212 345572 264
rect 345624 252 345630 264
rect 354950 252 354956 264
rect 345624 224 354956 252
rect 345624 212 345630 224
rect 354950 212 354956 224
rect 355008 212 355014 264
rect 355870 212 355876 264
rect 355928 252 355934 264
rect 365990 252 365996 264
rect 355928 224 365996 252
rect 355928 212 355934 224
rect 365990 212 365996 224
rect 366048 212 366054 264
rect 381998 212 382004 264
rect 382056 252 382062 264
rect 393222 252 393228 264
rect 382056 224 393228 252
rect 382056 212 382062 224
rect 393222 212 393228 224
rect 393280 212 393286 264
rect 393958 212 393964 264
rect 394016 252 394022 264
rect 396046 252 396074 360
rect 398576 320 398604 360
rect 401134 348 401140 400
rect 401192 388 401198 400
rect 404909 391 404967 397
rect 401192 360 404768 388
rect 401192 348 401198 360
rect 403805 323 403863 329
rect 403805 320 403817 323
rect 398576 292 403817 320
rect 403805 289 403817 292
rect 403851 289 403863 323
rect 403805 283 403863 289
rect 394016 224 396074 252
rect 394016 212 394022 224
rect 397454 212 397460 264
rect 397512 252 397518 264
rect 404740 252 404768 360
rect 404909 357 404921 391
rect 404955 388 404967 391
rect 411714 388 411720 400
rect 404955 360 411720 388
rect 404955 357 404967 360
rect 404909 351 404967 357
rect 411714 348 411720 360
rect 411772 348 411778 400
rect 424686 348 424692 400
rect 424744 388 424750 400
rect 432984 388 433012 428
rect 433058 416 433064 468
rect 433116 456 433122 468
rect 445726 456 445754 564
rect 446214 552 446220 564
rect 446272 552 446278 604
rect 446674 592 446680 604
rect 446635 564 446680 592
rect 446674 552 446680 564
rect 446732 552 446738 604
rect 447870 552 447876 604
rect 447928 592 447934 604
rect 451645 595 451703 601
rect 451645 592 451657 595
rect 447928 564 451657 592
rect 447928 552 447934 564
rect 451645 561 451657 564
rect 451691 561 451703 595
rect 451645 555 451703 561
rect 451921 595 451979 601
rect 451921 561 451933 595
rect 451967 592 451979 595
rect 456061 595 456119 601
rect 456061 592 456073 595
rect 451967 564 456073 592
rect 451967 561 451979 564
rect 451921 555 451979 561
rect 456061 561 456073 564
rect 456107 561 456119 595
rect 458082 592 458088 604
rect 458043 564 458088 592
rect 456061 555 456119 561
rect 458082 552 458088 564
rect 458140 552 458146 604
rect 461486 592 461492 604
rect 461447 564 461492 592
rect 461486 552 461492 564
rect 461544 552 461550 604
rect 463602 552 463608 604
rect 463660 592 463666 604
rect 469186 592 469214 632
rect 477862 620 477868 632
rect 477920 620 477926 672
rect 482922 620 482928 672
rect 482980 620 482986 672
rect 483014 620 483020 672
rect 483072 660 483078 672
rect 484026 660 484032 672
rect 483072 632 483117 660
rect 483987 632 484032 660
rect 483072 620 483078 632
rect 484026 620 484032 632
rect 484084 620 484090 672
rect 485317 663 485375 669
rect 485317 660 485329 663
rect 485148 632 485329 660
rect 485148 604 485176 632
rect 485317 629 485329 632
rect 485363 629 485375 663
rect 486602 660 486608 672
rect 486563 632 486608 660
rect 485317 623 485375 629
rect 486602 620 486608 632
rect 486660 620 486666 672
rect 487430 660 487436 672
rect 487391 632 487436 660
rect 487430 620 487436 632
rect 487488 620 487494 672
rect 487614 660 487620 672
rect 487575 632 487620 660
rect 487614 620 487620 632
rect 487672 620 487678 672
rect 488258 660 488264 672
rect 488219 632 488264 660
rect 488258 620 488264 632
rect 488316 620 488322 672
rect 489886 660 489914 700
rect 498212 672 498240 836
rect 509881 833 509893 867
rect 509927 864 509939 867
rect 521749 867 521807 873
rect 521749 864 521761 867
rect 509927 836 521761 864
rect 509927 833 509939 836
rect 509881 827 509939 833
rect 521749 833 521761 836
rect 521795 833 521807 867
rect 521749 827 521807 833
rect 510249 799 510307 805
rect 510249 765 510261 799
rect 510295 796 510307 799
rect 523037 799 523095 805
rect 523037 796 523049 799
rect 510295 768 523049 796
rect 510295 765 510307 768
rect 510249 759 510307 765
rect 523037 765 523049 768
rect 523083 765 523095 799
rect 523037 759 523095 765
rect 504177 731 504235 737
rect 504177 697 504189 731
rect 504223 728 504235 731
rect 510893 731 510951 737
rect 510893 728 510905 731
rect 504223 700 510905 728
rect 504223 697 504235 700
rect 504177 691 504235 697
rect 510893 697 510905 700
rect 510939 697 510951 731
rect 521657 731 521715 737
rect 521657 728 521669 731
rect 510893 691 510951 697
rect 511000 700 521669 728
rect 511000 672 511028 700
rect 521657 697 521669 700
rect 521703 697 521715 731
rect 523313 731 523371 737
rect 523313 728 523325 731
rect 521657 691 521715 697
rect 522776 700 523325 728
rect 492674 660 492680 672
rect 489886 632 492680 660
rect 492674 620 492680 632
rect 492732 620 492738 672
rect 496814 660 496820 672
rect 496775 632 496820 660
rect 496814 620 496820 632
rect 496872 620 496878 672
rect 498194 620 498200 672
rect 498252 620 498258 672
rect 498930 660 498936 672
rect 498891 632 498936 660
rect 498930 620 498936 632
rect 498988 620 498994 672
rect 502334 660 502340 672
rect 502295 632 502340 660
rect 502334 620 502340 632
rect 502392 620 502398 672
rect 502978 660 502984 672
rect 502939 632 502984 660
rect 502978 620 502984 632
rect 503036 620 503042 672
rect 505738 660 505744 672
rect 505699 632 505744 660
rect 505738 620 505744 632
rect 505796 620 505802 672
rect 507854 620 507860 672
rect 507912 660 507918 672
rect 509878 660 509884 672
rect 507912 632 507957 660
rect 509839 632 509884 660
rect 507912 620 507918 632
rect 509878 620 509884 632
rect 509936 620 509942 672
rect 510982 620 510988 672
rect 511040 620 511046 672
rect 512454 660 512460 672
rect 511092 632 512460 660
rect 470594 592 470600 604
rect 463660 564 469214 592
rect 470555 564 470600 592
rect 463660 552 463666 564
rect 470594 552 470600 564
rect 470652 552 470658 604
rect 471698 592 471704 604
rect 471659 564 471704 592
rect 471698 552 471704 564
rect 471756 552 471762 604
rect 472250 592 472256 604
rect 472211 564 472256 592
rect 472250 552 472256 564
rect 472308 552 472314 604
rect 474550 592 474556 604
rect 474511 564 474556 592
rect 474550 552 474556 564
rect 474608 552 474614 604
rect 475746 592 475752 604
rect 475707 564 475752 592
rect 475746 552 475752 564
rect 475804 552 475810 604
rect 476942 592 476948 604
rect 476903 564 476948 592
rect 476942 552 476948 564
rect 477000 552 477006 604
rect 481726 592 481732 604
rect 481687 564 481732 592
rect 481726 552 481732 564
rect 481784 552 481790 604
rect 485130 552 485136 604
rect 485188 552 485194 604
rect 485225 595 485283 601
rect 485225 561 485237 595
rect 485271 592 485283 595
rect 485406 592 485412 604
rect 485271 564 485412 592
rect 485271 561 485283 564
rect 485225 555 485283 561
rect 485406 552 485412 564
rect 485464 552 485470 604
rect 486326 552 486332 604
rect 486384 592 486390 604
rect 490926 592 490932 604
rect 486384 564 490788 592
rect 490887 564 490932 592
rect 486384 552 486390 564
rect 455874 524 455880 536
rect 433116 428 445754 456
rect 449176 496 455880 524
rect 433116 416 433122 428
rect 443638 388 443644 400
rect 424744 360 432644 388
rect 432984 360 443644 388
rect 424744 348 424750 360
rect 406930 280 406936 332
rect 406988 320 406994 332
rect 406988 292 415164 320
rect 406988 280 406994 292
rect 412910 252 412916 264
rect 397512 224 403112 252
rect 404740 224 412916 252
rect 397512 212 397518 224
rect 345934 184 345940 196
rect 338356 156 340368 184
rect 342226 156 345940 184
rect 338356 144 338362 156
rect 184348 88 184934 116
rect 184348 76 184354 88
rect 185486 76 185492 128
rect 185544 116 185550 128
rect 188246 116 188252 128
rect 185544 88 188252 116
rect 185544 76 185550 88
rect 188246 76 188252 88
rect 188304 76 188310 128
rect 227346 76 227352 128
rect 227404 116 227410 128
rect 232038 116 232044 128
rect 227404 88 232044 116
rect 227404 76 227410 88
rect 232038 76 232044 88
rect 232096 76 232102 128
rect 252002 76 252008 128
rect 252060 116 252066 128
rect 257246 116 257252 128
rect 252060 88 257252 116
rect 252060 76 252066 88
rect 257246 76 257252 88
rect 257304 76 257310 128
rect 266078 76 266084 128
rect 266136 116 266142 128
rect 272150 116 272156 128
rect 266136 88 272156 116
rect 266136 76 266142 88
rect 272150 76 272156 88
rect 272208 76 272214 128
rect 286410 76 286416 128
rect 286468 116 286474 128
rect 291562 116 291568 128
rect 286468 88 291568 116
rect 286468 76 286474 88
rect 291562 76 291568 88
rect 291620 76 291626 128
rect 299014 76 299020 128
rect 299072 116 299078 128
rect 306926 116 306932 128
rect 299072 88 306932 116
rect 299072 76 299078 88
rect 306926 76 306932 88
rect 306984 76 306990 128
rect 320634 76 320640 128
rect 320692 116 320698 128
rect 329006 116 329012 128
rect 320692 88 329012 116
rect 320692 76 320698 88
rect 329006 76 329012 88
rect 329064 76 329070 128
rect 329742 76 329748 128
rect 329800 116 329806 128
rect 338669 119 338727 125
rect 338669 116 338681 119
rect 329800 88 338681 116
rect 329800 76 329806 88
rect 338669 85 338681 88
rect 338715 85 338727 119
rect 340340 116 340368 156
rect 345934 144 345940 156
rect 345992 144 345998 196
rect 347406 144 347412 196
rect 347464 184 347470 196
rect 357342 184 357348 196
rect 347464 156 357348 184
rect 347464 144 347470 156
rect 357342 144 357348 156
rect 357400 144 357406 196
rect 358078 144 358084 196
rect 358136 184 358142 196
rect 358136 156 360884 184
rect 358136 144 358142 156
rect 347682 116 347688 128
rect 340340 88 347688 116
rect 338669 79 338727 85
rect 347682 76 347688 88
rect 347740 76 347746 128
rect 350166 76 350172 128
rect 350224 116 350230 128
rect 359734 116 359740 128
rect 350224 88 359740 116
rect 350224 76 350230 88
rect 359734 76 359740 88
rect 359792 76 359798 128
rect 360856 116 360884 156
rect 361482 144 361488 196
rect 361540 184 361546 196
rect 371970 184 371976 196
rect 361540 156 371976 184
rect 361540 144 361546 156
rect 371970 144 371976 156
rect 372028 144 372034 196
rect 380802 144 380808 196
rect 380860 184 380866 196
rect 385770 184 385776 196
rect 380860 156 385776 184
rect 380860 144 380866 156
rect 385770 144 385776 156
rect 385828 144 385834 196
rect 386506 144 386512 196
rect 386564 184 386570 196
rect 397733 187 397791 193
rect 397733 184 397745 187
rect 386564 156 397745 184
rect 386564 144 386570 156
rect 397733 153 397745 156
rect 397779 153 397791 187
rect 403084 184 403112 224
rect 412910 212 412916 224
rect 412968 212 412974 264
rect 415136 252 415164 292
rect 416038 280 416044 332
rect 416096 320 416102 332
rect 428642 320 428648 332
rect 416096 292 428648 320
rect 416096 280 416102 292
rect 428642 280 428648 292
rect 428700 280 428706 332
rect 432616 320 432644 360
rect 443638 348 443644 360
rect 443696 348 443702 400
rect 437566 320 437572 332
rect 432616 292 437572 320
rect 437566 280 437572 292
rect 437624 280 437630 332
rect 442166 280 442172 332
rect 442224 320 442230 332
rect 449176 320 449204 496
rect 455874 484 455880 496
rect 455932 484 455938 536
rect 459002 484 459008 536
rect 459060 524 459066 536
rect 459060 496 465764 524
rect 459060 484 459066 496
rect 449897 459 449955 465
rect 449897 425 449909 459
rect 449943 456 449955 459
rect 450630 456 450636 468
rect 449943 428 450636 456
rect 449943 425 449955 428
rect 449897 419 449955 425
rect 450630 416 450636 428
rect 450688 416 450694 468
rect 451645 459 451703 465
rect 451645 425 451657 459
rect 451691 456 451703 459
rect 459554 456 459560 468
rect 451691 428 459560 456
rect 451691 425 451703 428
rect 451645 419 451703 425
rect 459554 416 459560 428
rect 459612 416 459618 468
rect 460198 416 460204 468
rect 460256 456 460262 468
rect 465629 459 465687 465
rect 465629 456 465641 459
rect 460256 428 465641 456
rect 460256 416 460262 428
rect 465629 425 465641 428
rect 465675 425 465687 459
rect 465629 419 465687 425
rect 449618 348 449624 400
rect 449676 388 449682 400
rect 451921 391 451979 397
rect 451921 388 451933 391
rect 449676 360 451933 388
rect 449676 348 449682 360
rect 451921 357 451933 360
rect 451967 357 451979 391
rect 452286 388 452292 400
rect 452247 360 452292 388
rect 451921 351 451979 357
rect 452286 348 452292 360
rect 452344 348 452350 400
rect 452378 348 452384 400
rect 452436 388 452442 400
rect 452436 360 456794 388
rect 452436 348 452442 360
rect 442224 292 449204 320
rect 442224 280 442230 292
rect 451274 280 451280 332
rect 451332 320 451338 332
rect 456766 320 456794 360
rect 457898 348 457904 400
rect 457956 388 457962 400
rect 465736 388 465764 496
rect 477402 484 477408 536
rect 477460 524 477466 536
rect 489270 524 489276 536
rect 477460 496 489276 524
rect 477460 484 477466 496
rect 489270 484 489276 496
rect 489328 484 489334 536
rect 490760 524 490788 564
rect 490926 552 490932 564
rect 490984 552 490990 604
rect 491110 592 491116 604
rect 491071 564 491116 592
rect 491110 552 491116 564
rect 491168 552 491174 604
rect 501782 592 501788 604
rect 495406 564 501788 592
rect 495406 524 495434 564
rect 501782 552 501788 564
rect 501840 552 501846 604
rect 503809 595 503867 601
rect 503809 561 503821 595
rect 503855 592 503867 595
rect 510246 592 510252 604
rect 503855 564 510252 592
rect 503855 561 503867 564
rect 503809 555 503867 561
rect 510246 552 510252 564
rect 510304 552 510310 604
rect 490760 496 495434 524
rect 496722 484 496728 536
rect 496780 524 496786 536
rect 511092 524 511120 632
rect 512454 620 512460 632
rect 512512 620 512518 672
rect 514386 660 514392 672
rect 514347 632 514392 660
rect 514386 620 514392 632
rect 514444 620 514450 672
rect 514481 663 514539 669
rect 514481 629 514493 663
rect 514527 660 514539 663
rect 515950 660 515956 672
rect 514527 632 515956 660
rect 514527 629 514539 632
rect 514481 623 514539 629
rect 515950 620 515956 632
rect 516008 620 516014 672
rect 516962 660 516968 672
rect 516923 632 516968 660
rect 516962 620 516968 632
rect 517020 620 517026 672
rect 518250 660 518256 672
rect 518211 632 518256 660
rect 518250 620 518256 632
rect 518308 620 518314 672
rect 518342 620 518348 672
rect 518400 660 518406 672
rect 518400 632 518445 660
rect 518400 620 518406 632
rect 519446 620 519452 672
rect 519504 660 519510 672
rect 520734 660 520740 672
rect 519504 632 520596 660
rect 520695 632 520740 660
rect 519504 620 519510 632
rect 513558 552 513564 604
rect 513616 552 513622 604
rect 513653 595 513711 601
rect 513653 561 513665 595
rect 513699 592 513711 595
rect 519538 592 519544 604
rect 513699 564 519544 592
rect 513699 561 513711 564
rect 513653 555 513711 561
rect 519538 552 519544 564
rect 519596 552 519602 604
rect 520568 592 520596 632
rect 520734 620 520740 632
rect 520792 620 520798 672
rect 521930 620 521936 672
rect 521988 660 521994 672
rect 521988 632 522033 660
rect 521988 620 521994 632
rect 522776 592 522804 700
rect 523313 697 523325 700
rect 523359 697 523371 731
rect 523313 691 523371 697
rect 522850 620 522856 672
rect 522908 660 522914 672
rect 523420 660 523448 972
rect 539781 969 539793 972
rect 539827 969 539839 1003
rect 539781 963 539839 969
rect 557997 1003 558055 1009
rect 557997 969 558009 1003
rect 558043 1000 558055 1003
rect 569862 1000 569868 1012
rect 558043 972 569868 1000
rect 558043 969 558055 972
rect 557997 963 558055 969
rect 569862 960 569868 972
rect 569920 960 569926 1012
rect 540793 935 540851 941
rect 540793 932 540805 935
rect 523512 904 540805 932
rect 523512 672 523540 904
rect 540793 901 540805 904
rect 540839 901 540851 935
rect 540793 895 540851 901
rect 551097 935 551155 941
rect 551097 901 551109 935
rect 551143 932 551155 935
rect 569126 932 569132 944
rect 551143 904 569132 932
rect 551143 901 551155 904
rect 551097 895 551155 901
rect 569126 892 569132 904
rect 569184 892 569190 944
rect 538769 867 538827 873
rect 538769 833 538781 867
rect 538815 864 538827 867
rect 542449 867 542507 873
rect 542449 864 542461 867
rect 538815 836 542461 864
rect 538815 833 538827 836
rect 538769 827 538827 833
rect 542449 833 542461 836
rect 542495 833 542507 867
rect 566826 864 566832 876
rect 542449 827 542507 833
rect 550606 836 566832 864
rect 541989 799 542047 805
rect 541989 796 542001 799
rect 527146 768 542001 796
rect 527146 728 527174 768
rect 541989 765 542001 768
rect 542035 765 542047 799
rect 541989 759 542047 765
rect 542357 799 542415 805
rect 542357 765 542369 799
rect 542403 796 542415 799
rect 542403 768 546494 796
rect 542403 765 542415 768
rect 542357 759 542415 765
rect 525076 700 527174 728
rect 538217 731 538275 737
rect 522908 632 523448 660
rect 522908 620 522914 632
rect 523494 620 523500 672
rect 523552 620 523558 672
rect 524969 663 525027 669
rect 524969 660 524981 663
rect 523604 632 524981 660
rect 523034 592 523040 604
rect 520568 564 522804 592
rect 522995 564 523040 592
rect 523034 552 523040 564
rect 523092 552 523098 604
rect 496780 496 511120 524
rect 511169 527 511227 533
rect 496780 484 496786 496
rect 511169 493 511181 527
rect 511215 524 511227 527
rect 513576 524 513604 552
rect 523604 524 523632 632
rect 524969 629 524981 632
rect 525015 629 525027 663
rect 524969 623 525027 629
rect 525076 604 525104 700
rect 538217 697 538229 731
rect 538263 728 538275 731
rect 543369 731 543427 737
rect 543369 728 543381 731
rect 538263 700 543381 728
rect 538263 697 538275 700
rect 538217 691 538275 697
rect 543369 697 543381 700
rect 543415 697 543427 731
rect 546466 728 546494 768
rect 549257 731 549315 737
rect 549257 728 549269 731
rect 546466 700 549269 728
rect 543369 691 543427 697
rect 549257 697 549269 700
rect 549303 697 549315 731
rect 549257 691 549315 697
rect 525153 663 525211 669
rect 525153 629 525165 663
rect 525199 660 525211 663
rect 530118 660 530124 672
rect 525199 632 530124 660
rect 525199 629 525211 632
rect 525153 623 525211 629
rect 530118 620 530124 632
rect 530176 620 530182 672
rect 531130 660 531136 672
rect 531091 632 531136 660
rect 531130 620 531136 632
rect 531188 620 531194 672
rect 531314 660 531320 672
rect 531275 632 531320 660
rect 531314 620 531320 632
rect 531372 620 531378 672
rect 531866 620 531872 672
rect 531924 660 531930 672
rect 548334 660 548340 672
rect 531924 632 548340 660
rect 531924 620 531930 632
rect 548334 620 548340 632
rect 548392 620 548398 672
rect 548978 620 548984 672
rect 549036 660 549042 672
rect 550606 660 550634 836
rect 566826 824 566832 836
rect 566884 824 566890 876
rect 551557 799 551615 805
rect 551557 765 551569 799
rect 551603 796 551615 799
rect 568022 796 568028 808
rect 551603 768 568028 796
rect 551603 765 551615 768
rect 551557 759 551615 765
rect 568022 756 568028 768
rect 568080 756 568086 808
rect 570322 728 570328 740
rect 552400 700 570328 728
rect 552400 672 552428 700
rect 570322 688 570328 700
rect 570380 688 570386 740
rect 551094 660 551100 672
rect 549036 632 550634 660
rect 551055 632 551100 660
rect 549036 620 549042 632
rect 551094 620 551100 632
rect 551152 620 551158 672
rect 551204 632 552336 660
rect 524230 592 524236 604
rect 524191 564 524236 592
rect 524230 552 524236 564
rect 524288 552 524294 604
rect 525058 552 525064 604
rect 525116 552 525122 604
rect 526254 552 526260 604
rect 526312 592 526318 604
rect 538217 595 538275 601
rect 538217 592 538229 595
rect 526312 564 538229 592
rect 526312 552 526318 564
rect 538217 561 538229 564
rect 538263 561 538275 595
rect 538766 592 538772 604
rect 538727 564 538772 592
rect 538217 555 538275 561
rect 538766 552 538772 564
rect 538824 552 538830 604
rect 540790 592 540796 604
rect 540751 564 540796 592
rect 540790 552 540796 564
rect 540848 552 540854 604
rect 541986 592 541992 604
rect 541947 564 541992 592
rect 541986 552 541992 564
rect 542044 552 542050 604
rect 543090 552 543096 604
rect 543148 552 543154 604
rect 543366 552 543372 604
rect 543424 592 543430 604
rect 544194 592 544200 604
rect 543424 564 543469 592
rect 544155 564 544200 592
rect 543424 552 543430 564
rect 544194 552 544200 564
rect 544252 552 544258 604
rect 544378 592 544384 604
rect 544339 564 544384 592
rect 544378 552 544384 564
rect 544436 552 544442 604
rect 545114 592 545120 604
rect 545075 564 545120 592
rect 545114 552 545120 564
rect 545172 552 545178 604
rect 545482 592 545488 604
rect 545443 564 545488 592
rect 545482 552 545488 564
rect 545540 552 545546 604
rect 551204 592 551232 632
rect 546466 564 551232 592
rect 552308 592 552336 632
rect 552382 620 552388 672
rect 552440 620 552446 672
rect 552477 663 552535 669
rect 552477 629 552489 663
rect 552523 660 552535 663
rect 565630 660 565636 672
rect 552523 632 565636 660
rect 552523 629 552535 632
rect 552477 623 552535 629
rect 565630 620 565636 632
rect 565688 620 565694 672
rect 560846 592 560852 604
rect 552308 564 560852 592
rect 511215 496 513604 524
rect 514726 496 523632 524
rect 523681 527 523739 533
rect 511215 493 511227 496
rect 511169 487 511227 493
rect 469214 416 469220 468
rect 469272 456 469278 468
rect 484029 459 484087 465
rect 484029 456 484041 459
rect 469272 428 484041 456
rect 469272 416 469278 428
rect 484029 425 484041 428
rect 484075 425 484087 459
rect 484029 419 484087 425
rect 495342 416 495348 468
rect 495400 456 495406 468
rect 504177 459 504235 465
rect 504177 456 504189 459
rect 495400 428 504189 456
rect 495400 416 495406 428
rect 504177 425 504189 428
rect 504223 425 504235 459
rect 504634 456 504640 468
rect 504595 428 504640 456
rect 504177 419 504235 425
rect 504634 416 504640 428
rect 504692 416 504698 468
rect 506198 456 506204 468
rect 506159 428 506204 456
rect 506198 416 506204 428
rect 506256 416 506262 468
rect 506934 416 506940 468
rect 506992 456 506998 468
rect 509694 456 509700 468
rect 506992 428 509700 456
rect 506992 416 506998 428
rect 509694 416 509700 428
rect 509752 416 509758 468
rect 510893 459 510951 465
rect 510893 425 510905 459
rect 510939 456 510951 459
rect 511442 456 511448 468
rect 510939 428 511448 456
rect 510939 425 510951 428
rect 510893 419 510951 425
rect 511442 416 511448 428
rect 511500 416 511506 468
rect 513282 416 513288 468
rect 513340 456 513346 468
rect 514726 456 514754 496
rect 523681 493 523693 527
rect 523727 524 523739 527
rect 523727 496 528554 524
rect 523727 493 523739 496
rect 523681 487 523739 493
rect 514938 456 514944 468
rect 513340 428 514754 456
rect 514899 428 514944 456
rect 513340 416 513346 428
rect 514938 416 514944 428
rect 514996 416 515002 468
rect 521657 459 521715 465
rect 521657 425 521669 459
rect 521703 456 521715 459
rect 527542 456 527548 468
rect 521703 428 527548 456
rect 521703 425 521715 428
rect 521657 419 521715 425
rect 527542 416 527548 428
rect 527600 416 527606 468
rect 528526 456 528554 496
rect 533062 484 533068 536
rect 533120 524 533126 536
rect 538493 527 538551 533
rect 538493 524 538505 527
rect 533120 496 538505 524
rect 533120 484 533126 496
rect 538493 493 538505 496
rect 538539 493 538551 527
rect 539778 524 539784 536
rect 539739 496 539784 524
rect 538493 487 538551 493
rect 539778 484 539784 496
rect 539836 484 539842 536
rect 543108 524 543136 552
rect 546466 524 546494 564
rect 560846 552 560852 564
rect 560904 552 560910 604
rect 562042 592 562048 604
rect 562003 564 562048 592
rect 562042 552 562048 564
rect 562100 552 562106 604
rect 563238 592 563244 604
rect 563199 564 563244 592
rect 563238 552 563244 564
rect 563296 552 563302 604
rect 573910 552 573916 604
rect 573968 552 573974 604
rect 575106 552 575112 604
rect 575164 552 575170 604
rect 549254 524 549260 536
rect 543108 496 546494 524
rect 549215 496 549260 524
rect 549254 484 549260 496
rect 549312 484 549318 536
rect 550082 484 550088 536
rect 550140 524 550146 536
rect 551557 527 551615 533
rect 551557 524 551569 527
rect 550140 496 551569 524
rect 550140 484 550146 496
rect 551557 493 551569 496
rect 551603 493 551615 527
rect 554590 524 554596 536
rect 554551 496 554596 524
rect 551557 487 551615 493
rect 554590 484 554596 496
rect 554648 484 554654 536
rect 555786 484 555792 536
rect 555844 524 555850 536
rect 573928 524 573956 552
rect 555844 496 573956 524
rect 555844 484 555850 496
rect 535822 456 535828 468
rect 528526 428 535828 456
rect 535822 416 535828 428
rect 535880 416 535886 468
rect 536466 416 536472 468
rect 536524 456 536530 468
rect 553486 456 553492 468
rect 536524 428 553492 456
rect 536524 416 536530 428
rect 553486 416 553492 428
rect 553544 416 553550 468
rect 556890 416 556896 468
rect 556948 456 556954 468
rect 575124 456 575152 552
rect 556948 428 575152 456
rect 556948 416 556954 428
rect 473262 388 473268 400
rect 457956 360 465672 388
rect 465736 360 473268 388
rect 457956 348 457962 360
rect 465350 320 465356 332
rect 451332 292 455414 320
rect 456766 292 465356 320
rect 451332 280 451338 292
rect 418798 252 418804 264
rect 415136 224 418804 252
rect 418798 212 418804 224
rect 418856 212 418862 264
rect 421742 212 421748 264
rect 421800 252 421806 264
rect 434070 252 434076 264
rect 421800 224 434076 252
rect 421800 212 421806 224
rect 434070 212 434076 224
rect 434128 212 434134 264
rect 434165 255 434223 261
rect 434165 221 434177 255
rect 434211 252 434223 255
rect 442629 255 442687 261
rect 442629 252 442641 255
rect 434211 224 442641 252
rect 434211 221 434223 224
rect 434165 215 434223 221
rect 442629 221 442641 224
rect 442675 221 442687 255
rect 442629 215 442687 221
rect 443270 212 443276 264
rect 443328 252 443334 264
rect 454773 255 454831 261
rect 454773 252 454785 255
rect 443328 224 454785 252
rect 443328 212 443334 224
rect 454773 221 454785 224
rect 454819 221 454831 255
rect 455386 252 455414 292
rect 465350 280 465356 292
rect 465408 280 465414 332
rect 465644 320 465672 360
rect 473262 348 473268 360
rect 473320 348 473326 400
rect 487617 391 487675 397
rect 487617 388 487629 391
rect 474706 360 487629 388
rect 472253 323 472311 329
rect 472253 320 472265 323
rect 465644 292 472265 320
rect 472253 289 472265 292
rect 472299 289 472311 323
rect 472253 283 472311 289
rect 472802 280 472808 332
rect 472860 320 472866 332
rect 474706 320 474734 360
rect 487617 357 487629 360
rect 487663 357 487675 391
rect 487617 351 487675 357
rect 487798 348 487804 400
rect 487856 388 487862 400
rect 492582 388 492588 400
rect 487856 360 492588 388
rect 487856 348 487862 360
rect 492582 348 492588 360
rect 492640 348 492646 400
rect 494422 348 494428 400
rect 494480 388 494486 400
rect 503809 391 503867 397
rect 503809 388 503821 391
rect 494480 360 503821 388
rect 494480 348 494486 360
rect 503809 357 503821 360
rect 503855 357 503867 391
rect 503990 388 503996 400
rect 503951 360 503996 388
rect 503809 351 503867 357
rect 503990 348 503996 360
rect 504048 348 504054 400
rect 509234 348 509240 400
rect 509292 388 509298 400
rect 525242 388 525248 400
rect 509292 360 525248 388
rect 509292 348 509298 360
rect 525242 348 525248 360
rect 525300 348 525306 400
rect 527174 348 527180 400
rect 527232 388 527238 400
rect 544381 391 544439 397
rect 544381 388 544393 391
rect 527232 360 544393 388
rect 527232 348 527238 360
rect 544381 357 544393 360
rect 544427 357 544439 391
rect 544381 351 544439 357
rect 547690 348 547696 400
rect 547748 388 547754 400
rect 552477 391 552535 397
rect 552477 388 552489 391
rect 547748 360 552489 388
rect 547748 348 547754 360
rect 552477 357 552489 360
rect 552523 357 552535 391
rect 552477 351 552535 357
rect 553302 348 553308 400
rect 553360 388 553366 400
rect 571150 388 571156 400
rect 553360 360 571156 388
rect 553360 348 553366 360
rect 571150 348 571156 360
rect 571208 348 571214 400
rect 472860 292 474734 320
rect 472860 280 472866 292
rect 483750 280 483756 332
rect 483808 320 483814 332
rect 495526 320 495532 332
rect 483808 292 495532 320
rect 483808 280 483814 292
rect 495526 280 495532 292
rect 495584 280 495590 332
rect 497826 280 497832 332
rect 497884 320 497890 332
rect 511169 323 511227 329
rect 511169 320 511181 323
rect 497884 292 511181 320
rect 497884 280 497890 292
rect 511169 289 511181 292
rect 511215 289 511227 323
rect 511169 283 511227 289
rect 520366 280 520372 332
rect 520424 320 520430 332
rect 536926 320 536932 332
rect 520424 292 536932 320
rect 520424 280 520430 292
rect 536926 280 536932 292
rect 536984 280 536990 332
rect 541710 280 541716 332
rect 541768 320 541774 332
rect 542357 323 542415 329
rect 542357 320 542369 323
rect 541768 292 542369 320
rect 541768 280 541774 292
rect 542357 289 542369 292
rect 542403 289 542415 323
rect 542357 283 542415 289
rect 542449 323 542507 329
rect 542449 289 542461 323
rect 542495 320 542507 323
rect 555878 320 555884 332
rect 542495 292 555884 320
rect 542495 289 542507 292
rect 542449 283 542507 289
rect 555878 280 555884 292
rect 555936 280 555942 332
rect 557994 320 558000 332
rect 557955 292 558000 320
rect 557994 280 558000 292
rect 558052 280 558058 332
rect 559006 280 559012 332
rect 559064 320 559070 332
rect 576762 320 576768 332
rect 559064 292 576768 320
rect 559064 280 559070 292
rect 576762 280 576768 292
rect 576820 280 576826 332
rect 463050 252 463056 264
rect 455386 224 463056 252
rect 454773 215 454831 221
rect 463050 212 463056 224
rect 463108 212 463114 264
rect 464890 212 464896 264
rect 464948 252 464954 264
rect 464948 224 470594 252
rect 464948 212 464954 224
rect 409414 184 409420 196
rect 403084 156 409420 184
rect 397733 147 397791 153
rect 409414 144 409420 156
rect 409472 144 409478 196
rect 411530 144 411536 196
rect 411588 184 411594 196
rect 420917 187 420975 193
rect 420917 184 420929 187
rect 411588 156 420929 184
rect 411588 144 411594 156
rect 420917 153 420929 156
rect 420963 153 420975 187
rect 420917 147 420975 153
rect 422386 144 422392 196
rect 422444 184 422450 196
rect 434714 184 434720 196
rect 422444 156 434720 184
rect 422444 144 422450 156
rect 434714 144 434720 156
rect 434772 144 434778 196
rect 435358 144 435364 196
rect 435416 184 435422 196
rect 448238 184 448244 196
rect 435416 156 448244 184
rect 435416 144 435422 156
rect 448238 144 448244 156
rect 448296 144 448302 196
rect 448974 144 448980 196
rect 449032 184 449038 196
rect 462406 184 462412 196
rect 449032 156 462412 184
rect 449032 144 449038 156
rect 462406 144 462412 156
rect 462464 144 462470 196
rect 467834 184 467840 196
rect 465736 156 467840 184
rect 364889 119 364947 125
rect 364889 116 364901 119
rect 360856 88 364901 116
rect 364889 85 364901 88
rect 364935 85 364947 119
rect 364889 79 364947 85
rect 367830 76 367836 128
rect 367888 116 367894 128
rect 378686 116 378692 128
rect 367888 88 378692 116
rect 367888 76 367894 88
rect 378686 76 378692 88
rect 378744 76 378750 128
rect 379514 76 379520 128
rect 379572 116 379578 128
rect 390278 116 390284 128
rect 379572 88 390284 116
rect 379572 76 379578 88
rect 390278 76 390284 88
rect 390336 76 390342 128
rect 394053 119 394111 125
rect 394053 85 394065 119
rect 394099 116 394111 119
rect 395522 116 395528 128
rect 394099 88 395528 116
rect 394099 85 394111 88
rect 394053 79 394111 85
rect 395522 76 395528 88
rect 395580 76 395586 128
rect 396258 76 396264 128
rect 396316 116 396322 128
rect 402149 119 402207 125
rect 402149 116 402161 119
rect 396316 88 402161 116
rect 396316 76 396322 88
rect 402149 85 402161 88
rect 402195 85 402207 119
rect 402149 79 402207 85
rect 402330 76 402336 128
rect 402388 116 402394 128
rect 414293 119 414351 125
rect 414293 116 414305 119
rect 402388 88 414305 116
rect 402388 76 402394 88
rect 414293 85 414305 88
rect 414339 85 414351 119
rect 414293 79 414351 85
rect 419442 76 419448 128
rect 419500 116 419506 128
rect 432049 119 432107 125
rect 432049 116 432061 119
rect 419500 88 432061 116
rect 419500 76 419506 88
rect 432049 85 432061 88
rect 432095 85 432107 119
rect 432049 79 432107 85
rect 434254 76 434260 128
rect 434312 116 434318 128
rect 447134 116 447140 128
rect 434312 88 447140 116
rect 434312 76 434318 88
rect 447134 76 447140 88
rect 447192 76 447198 128
rect 453482 116 453488 128
rect 453443 88 453488 116
rect 453482 76 453488 88
rect 453540 76 453546 128
rect 456518 76 456524 128
rect 456576 116 456582 128
rect 465736 116 465764 156
rect 467834 144 467840 156
rect 467892 144 467898 196
rect 470566 184 470594 224
rect 478506 212 478512 264
rect 478564 252 478570 264
rect 490282 252 490288 264
rect 478564 224 490288 252
rect 478564 212 478570 224
rect 490282 212 490288 224
rect 490340 212 490346 264
rect 492122 212 492128 264
rect 492180 252 492186 264
rect 502702 252 502708 264
rect 492180 224 502708 252
rect 492180 212 492186 224
rect 502702 212 502708 224
rect 502760 212 502766 264
rect 503530 212 503536 264
rect 503588 252 503594 264
rect 513653 255 513711 261
rect 513653 252 513665 255
rect 503588 224 513665 252
rect 503588 212 503594 224
rect 513653 221 513665 224
rect 513699 221 513711 255
rect 528830 252 528836 264
rect 513653 215 513711 221
rect 518866 224 528836 252
rect 479518 184 479524 196
rect 470566 156 479524 184
rect 479518 144 479524 156
rect 479576 144 479582 196
rect 480806 144 480812 196
rect 480864 184 480870 196
rect 485133 187 485191 193
rect 485133 184 485145 187
rect 480864 156 485145 184
rect 480864 144 480870 156
rect 485133 153 485145 156
rect 485179 153 485191 187
rect 485133 147 485191 153
rect 489730 144 489736 196
rect 489788 184 489794 196
rect 505186 184 505192 196
rect 489788 156 505192 184
rect 489788 144 489794 156
rect 505186 144 505192 156
rect 505244 144 505250 196
rect 506934 144 506940 196
rect 506992 184 506998 196
rect 510249 187 510307 193
rect 510249 184 510261 187
rect 506992 156 510261 184
rect 506992 144 506998 156
rect 510249 153 510261 156
rect 510295 153 510307 187
rect 510249 147 510307 153
rect 512178 144 512184 196
rect 512236 184 512242 196
rect 518866 184 518894 224
rect 528830 212 528836 224
rect 528888 212 528894 264
rect 529658 212 529664 264
rect 529716 252 529722 264
rect 546494 252 546500 264
rect 529716 224 546500 252
rect 529716 212 529722 224
rect 546494 212 546500 224
rect 546552 212 546558 264
rect 562594 212 562600 264
rect 562652 252 562658 264
rect 581822 252 581828 264
rect 562652 224 581828 252
rect 562652 212 562658 224
rect 581822 212 581828 224
rect 581880 212 581886 264
rect 512236 156 518894 184
rect 512236 144 512242 156
rect 521562 144 521568 196
rect 521620 184 521626 196
rect 538030 184 538036 196
rect 521620 156 538036 184
rect 521620 144 521626 156
rect 538030 144 538036 156
rect 538088 144 538094 196
rect 539870 144 539876 196
rect 539928 184 539934 196
rect 557166 184 557172 196
rect 539928 156 557172 184
rect 539928 144 539934 156
rect 557166 144 557172 156
rect 557224 144 557230 196
rect 560202 144 560208 196
rect 560260 184 560266 196
rect 578326 184 578332 196
rect 560260 156 578332 184
rect 560260 144 560266 156
rect 578326 144 578332 156
rect 578384 144 578390 196
rect 456576 88 465764 116
rect 456576 76 456582 88
rect 465994 76 466000 128
rect 466052 116 466058 128
rect 480714 116 480720 128
rect 466052 88 480720 116
rect 466052 76 466058 88
rect 480714 76 480720 88
rect 480772 76 480778 128
rect 481450 76 481456 128
rect 481508 116 481514 128
rect 496814 116 496820 128
rect 481508 88 496820 116
rect 481508 76 481514 88
rect 496814 76 496820 88
rect 496872 76 496878 128
rect 500126 76 500132 128
rect 500184 116 500190 128
rect 514481 119 514539 125
rect 514481 116 514493 119
rect 500184 88 514493 116
rect 500184 76 500190 88
rect 514481 85 514493 88
rect 514527 85 514539 119
rect 514481 79 514539 85
rect 515582 76 515588 128
rect 515640 116 515646 128
rect 532326 116 532332 128
rect 515640 88 532332 116
rect 515640 76 515646 88
rect 532326 76 532332 88
rect 532384 76 532390 128
rect 534534 116 534540 128
rect 534495 88 534540 116
rect 534534 76 534540 88
rect 534592 76 534598 128
rect 538493 119 538551 125
rect 538493 85 538505 119
rect 538539 116 538551 119
rect 550450 116 550456 128
rect 538539 88 550456 116
rect 538539 85 538551 88
rect 538493 79 538551 85
rect 550450 76 550456 88
rect 550508 76 550514 128
rect 564618 116 564624 128
rect 553366 88 564624 116
rect 44082 8 44088 60
rect 44140 48 44146 60
rect 46198 48 46204 60
rect 44140 20 46204 48
rect 44140 8 44146 20
rect 46198 8 46204 20
rect 46256 8 46262 60
rect 215018 8 215024 60
rect 215076 48 215082 60
rect 219434 48 219440 60
rect 215076 20 219440 48
rect 215076 8 215082 20
rect 219434 8 219440 20
rect 219492 8 219498 60
rect 289814 8 289820 60
rect 289872 48 289878 60
rect 296990 48 296996 60
rect 289872 20 296996 48
rect 289872 8 289878 20
rect 296990 8 296996 20
rect 297048 8 297054 60
rect 314746 8 314752 60
rect 314804 48 314810 60
rect 322842 48 322848 60
rect 314804 20 322848 48
rect 314804 8 314810 20
rect 322842 8 322848 20
rect 322900 8 322906 60
rect 330846 8 330852 60
rect 330904 48 330910 60
rect 338761 51 338819 57
rect 338761 48 338773 51
rect 330904 20 338773 48
rect 330904 8 330910 20
rect 338761 17 338773 20
rect 338807 17 338819 51
rect 338761 11 338819 17
rect 339494 8 339500 60
rect 339552 48 339558 60
rect 348234 48 348240 60
rect 339552 20 348240 48
rect 339552 8 339558 20
rect 348234 8 348240 20
rect 348292 8 348298 60
rect 353570 8 353576 60
rect 353628 48 353634 60
rect 363690 48 363696 60
rect 353628 20 363696 48
rect 353628 8 353634 20
rect 363690 8 363696 20
rect 363748 8 363754 60
rect 376294 8 376300 60
rect 376352 48 376358 60
rect 386782 48 386788 60
rect 376352 20 386788 48
rect 376352 8 376358 20
rect 386782 8 386788 20
rect 386840 8 386846 60
rect 387610 8 387616 60
rect 387668 48 387674 60
rect 399110 48 399116 60
rect 387668 20 399116 48
rect 387668 8 387674 20
rect 399110 8 399116 20
rect 399168 8 399174 60
rect 399849 51 399907 57
rect 399849 17 399861 51
rect 399895 48 399907 51
rect 407022 48 407028 60
rect 399895 20 407028 48
rect 399895 17 399907 20
rect 399849 11 399907 17
rect 407022 8 407028 20
rect 407080 8 407086 60
rect 414934 8 414940 60
rect 414992 48 414998 60
rect 423861 51 423919 57
rect 423861 48 423873 51
rect 414992 20 423873 48
rect 414992 8 414998 20
rect 423861 17 423873 20
rect 423907 17 423919 51
rect 423861 11 423919 17
rect 426986 8 426992 60
rect 427044 48 427050 60
rect 440142 48 440148 60
rect 427044 20 440148 48
rect 427044 8 427050 20
rect 440142 8 440148 20
rect 440200 8 440206 60
rect 441062 8 441068 60
rect 441120 48 441126 60
rect 454497 51 454555 57
rect 454497 48 454509 51
rect 441120 20 454509 48
rect 441120 8 441126 20
rect 454497 17 454509 20
rect 454543 17 454555 51
rect 454497 11 454555 17
rect 455322 8 455328 60
rect 455380 48 455386 60
rect 469582 48 469588 60
rect 455380 20 469588 48
rect 455380 8 455386 20
rect 469582 8 469588 20
rect 469640 8 469646 60
rect 476206 8 476212 60
rect 476264 48 476270 60
rect 491113 51 491171 57
rect 491113 48 491125 51
rect 476264 20 491125 48
rect 476264 8 476270 20
rect 491113 17 491125 20
rect 491159 17 491171 51
rect 491113 11 491171 17
rect 493318 8 493324 60
rect 493376 48 493382 60
rect 508590 48 508596 60
rect 493376 20 508596 48
rect 493376 8 493382 20
rect 508590 8 508596 20
rect 508648 8 508654 60
rect 521749 51 521807 57
rect 521749 17 521761 51
rect 521795 48 521807 51
rect 526254 48 526260 60
rect 521795 20 526260 48
rect 521795 17 521807 20
rect 521749 11 521807 17
rect 526254 8 526260 20
rect 526312 8 526318 60
rect 528462 8 528468 60
rect 528520 48 528526 60
rect 545485 51 545543 57
rect 545485 48 545497 51
rect 528520 20 545497 48
rect 528520 8 528526 20
rect 545485 17 545497 20
rect 545531 17 545543 51
rect 545485 11 545543 17
rect 546494 8 546500 60
rect 546552 48 546558 60
rect 553366 48 553394 88
rect 564618 76 564624 88
rect 564676 76 564682 128
rect 546552 20 553394 48
rect 546552 8 546558 20
rect 561398 8 561404 60
rect 561456 48 561462 60
rect 580718 48 580724 60
rect 561456 20 580724 48
rect 561456 8 561462 20
rect 580718 8 580724 20
rect 580776 8 580782 60
<< via1 >>
rect 271788 703808 271840 703860
rect 364708 703808 364760 703860
rect 257252 703740 257304 703792
rect 371608 703740 371660 703792
rect 276848 703672 276900 703724
rect 332324 703672 332376 703724
rect 235356 703536 235408 703588
rect 300860 703604 300912 703656
rect 242440 703536 242492 703588
rect 400864 703536 400916 703588
rect 170312 703400 170364 703452
rect 315488 703468 315540 703520
rect 227628 703400 227680 703452
rect 497464 703400 497516 703452
rect 1492 703332 1544 703384
rect 359740 703332 359792 703384
rect 213000 703264 213052 703316
rect 576400 703264 576452 703316
rect 1584 703196 1636 703248
rect 374460 703196 374512 703248
rect 198280 703128 198332 703180
rect 575112 703128 575164 703180
rect 1676 703060 1728 703112
rect 389180 703060 389232 703112
rect 183376 702992 183428 703044
rect 573732 702992 573784 703044
rect 1860 702924 1912 702976
rect 403900 702924 403952 702976
rect 158628 702856 158680 702908
rect 575020 702856 575072 702908
rect 756 702788 808 702840
rect 423680 702788 423732 702840
rect 2320 702720 2372 702772
rect 477592 702720 477644 702772
rect 388 702652 440 702704
rect 497280 702652 497332 702704
rect 296 702584 348 702636
rect 507124 702584 507176 702636
rect 112 702516 164 702568
rect 536840 702516 536892 702568
rect 35808 702448 35860 702500
rect 574744 702448 574796 702500
rect 154028 702380 154080 702432
rect 311164 702380 311216 702432
rect 75460 702312 75512 702364
rect 573456 702312 573508 702364
rect 237104 702244 237156 702296
rect 305828 702244 305880 702296
rect 311072 702176 311124 702228
rect 364616 702176 364668 702228
rect 178592 702108 178644 702160
rect 339316 702108 339368 702160
rect 163872 702040 163924 702092
rect 331312 702040 331364 702092
rect 335912 702040 335964 702092
rect 467840 702040 467892 702092
rect 188436 701972 188488 702024
rect 243360 701972 243412 702024
rect 262128 701972 262180 702024
rect 482560 701972 482612 702024
rect 266360 701904 266412 701956
rect 502340 701904 502392 701956
rect 70124 701836 70176 701888
rect 329380 701836 329432 701888
rect 350540 701836 350592 701888
rect 512000 701836 512052 701888
rect 1308 701768 1360 701820
rect 414204 701768 414256 701820
rect 148968 701700 149020 701752
rect 577504 701700 577556 701752
rect 4344 701632 4396 701684
rect 443276 701632 443328 701684
rect 444288 701632 444340 701684
rect 541532 701632 541584 701684
rect 129464 701564 129516 701616
rect 574928 701564 574980 701616
rect 2596 701496 2648 701548
rect 458180 701496 458232 701548
rect 119712 701428 119764 701480
rect 576308 701428 576360 701480
rect 104808 701360 104860 701412
rect 574836 701360 574888 701412
rect 100024 701292 100076 701344
rect 576216 701292 576268 701344
rect 90180 701224 90232 701276
rect 573548 701224 573600 701276
rect 85304 701156 85356 701208
rect 569316 701156 569368 701208
rect 572 701088 624 701140
rect 487436 701088 487488 701140
rect 55772 701020 55824 701072
rect 271512 701020 271564 701072
rect 282920 701020 282972 701072
rect 291200 701020 291252 701072
rect 291384 701020 291436 701072
rect 295892 701020 295944 701072
rect 331220 701020 331272 701072
rect 335360 701020 335412 701072
rect 339408 701020 339460 701072
rect 344928 701020 344980 701072
rect 8116 700952 8168 701004
rect 349896 701020 349948 701072
rect 400864 700952 400916 701004
rect 494796 700952 494848 701004
rect 497464 700952 497516 701004
rect 559656 700952 559708 701004
rect 40500 700884 40552 700936
rect 339408 700884 339460 700936
rect 371608 700884 371660 700936
rect 429844 700884 429896 700936
rect 72976 700816 73028 700868
rect 331220 700816 331272 700868
rect 202788 700748 202840 700800
rect 305736 700748 305788 700800
rect 305828 700748 305880 700800
rect 543464 700748 543516 700800
rect 137836 700680 137888 700732
rect 320456 700680 320508 700732
rect 339316 700680 339368 700732
rect 580724 700680 580776 700732
rect 105452 700612 105504 700664
rect 330300 700612 330352 700664
rect 331312 700612 331364 700664
rect 580632 700612 580684 700664
rect 89168 700544 89220 700596
rect 340052 700544 340104 700596
rect 3884 700476 3936 700528
rect 262128 700476 262180 700528
rect 281356 700476 281408 700528
rect 348792 700476 348844 700528
rect 3700 700408 3752 700460
rect 266360 700408 266412 700460
rect 267648 700408 267700 700460
rect 282920 700408 282972 700460
rect 284116 700408 284168 700460
rect 291384 700408 291436 700460
rect 291476 700408 291528 700460
rect 300124 700408 300176 700460
rect 311164 700408 311216 700460
rect 580540 700408 580592 700460
rect 232688 700340 232740 700392
rect 527180 700340 527232 700392
rect 24308 700272 24360 700324
rect 354956 700272 355008 700324
rect 252284 700204 252336 700256
rect 478512 700204 478564 700256
rect 247086 700136 247138 700188
rect 462320 700136 462372 700188
rect 154120 700068 154172 700120
rect 325654 700068 325706 700120
rect 329380 700068 329432 700120
rect 580356 700068 580408 700120
rect 267004 700000 267056 700052
rect 413652 700000 413704 700052
rect 262128 699932 262180 699984
rect 397460 699932 397512 699984
rect 218980 699864 219032 699916
rect 310612 699864 310664 699916
rect 217876 699796 217928 699848
rect 563520 699796 563572 699848
rect 3240 699728 3292 699780
rect 369768 699728 369820 699780
rect 3792 699660 3844 699712
rect 384304 699660 384356 699712
rect 3056 699592 3108 699644
rect 311072 699592 311124 699644
rect 271512 699524 271564 699576
rect 580264 699524 580316 699576
rect 3976 699456 4028 699508
rect 335912 699456 335964 699508
rect 50896 699431 50948 699440
rect 50896 699397 50905 699431
rect 50905 699397 50939 699431
rect 50939 699397 50948 699431
rect 50896 699388 50948 699397
rect 65616 699431 65668 699440
rect 65616 699397 65625 699431
rect 65625 699397 65659 699431
rect 65659 699397 65668 699431
rect 65616 699388 65668 699397
rect 80152 699431 80204 699440
rect 80152 699397 80161 699431
rect 80161 699397 80195 699431
rect 80195 699397 80204 699431
rect 80152 699388 80204 699397
rect 95148 699431 95200 699440
rect 95148 699397 95157 699431
rect 95157 699397 95191 699431
rect 95191 699397 95200 699431
rect 95148 699388 95200 699397
rect 109868 699431 109920 699440
rect 109868 699397 109877 699431
rect 109877 699397 109911 699431
rect 109911 699397 109920 699431
rect 109868 699388 109920 699397
rect 114560 699431 114612 699440
rect 114560 699397 114569 699431
rect 114569 699397 114603 699431
rect 114603 699397 114612 699431
rect 114560 699388 114612 699397
rect 124588 699431 124640 699440
rect 124588 699397 124597 699431
rect 124597 699397 124631 699431
rect 124631 699397 124640 699431
rect 124588 699388 124640 699397
rect 139308 699431 139360 699440
rect 139308 699397 139317 699431
rect 139317 699397 139351 699431
rect 139351 699397 139360 699431
rect 139308 699388 139360 699397
rect 144276 699431 144328 699440
rect 144276 699397 144285 699431
rect 144285 699397 144319 699431
rect 144319 699397 144328 699431
rect 144276 699388 144328 699397
rect 168840 699431 168892 699440
rect 168840 699397 168849 699431
rect 168849 699397 168883 699431
rect 168883 699397 168892 699431
rect 168840 699388 168892 699397
rect 173716 699431 173768 699440
rect 173716 699397 173725 699431
rect 173725 699397 173759 699431
rect 173759 699397 173768 699431
rect 173716 699388 173768 699397
rect 3516 699320 3568 699372
rect 193220 699320 193272 699372
rect 202972 699320 203024 699372
rect 208124 699388 208176 699440
rect 222844 699320 222896 699372
rect 243360 699388 243412 699440
rect 580816 699388 580868 699440
rect 350540 699320 350592 699372
rect 394148 699363 394200 699372
rect 394148 699329 394157 699363
rect 394157 699329 394191 699363
rect 394191 699329 394200 699363
rect 394148 699320 394200 699329
rect 462872 699363 462924 699372
rect 462872 699329 462881 699363
rect 462881 699329 462915 699363
rect 462915 699329 462924 699363
rect 462872 699320 462924 699329
rect 492588 699363 492640 699372
rect 492588 699329 492597 699363
rect 492597 699329 492631 699363
rect 492631 699329 492640 699363
rect 492588 699320 492640 699329
rect 521844 699363 521896 699372
rect 521844 699329 521853 699363
rect 521853 699329 521887 699363
rect 521887 699329 521896 699363
rect 521844 699320 521896 699329
rect 563704 699252 563756 699304
rect 567844 699184 567896 699236
rect 578976 699116 579028 699168
rect 572168 699048 572220 699100
rect 848 698980 900 699032
rect 566832 698912 566884 698964
rect 573640 698844 573692 698896
rect 570696 698776 570748 698828
rect 578884 698708 578936 698760
rect 572076 698640 572128 698692
rect 570604 698572 570656 698624
rect 569500 698504 569552 698556
rect 565360 698436 565412 698488
rect 566740 698368 566792 698420
rect 566556 698300 566608 698352
rect 563520 698232 563572 698284
rect 580172 698232 580224 698284
rect 2412 697756 2464 697808
rect 480 697688 532 697740
rect 204 697620 256 697672
rect 573364 697552 573416 697604
rect 563704 684428 563756 684480
rect 580172 684428 580224 684480
rect 576400 671984 576452 672036
rect 580172 671984 580224 672036
rect 3240 661036 3292 661088
rect 4344 661036 4396 661088
rect 567844 632000 567896 632052
rect 580172 632000 580224 632052
rect 1308 619556 1360 619608
rect 2780 619556 2832 619608
rect 575112 618196 575164 618248
rect 580172 618196 580224 618248
rect 572168 578144 572220 578196
rect 579804 578144 579856 578196
rect 3792 565836 3844 565888
rect 4252 565836 4304 565888
rect 573732 564340 573784 564392
rect 580172 564340 580224 564392
rect 573640 538160 573692 538212
rect 580172 538160 580224 538212
rect 566832 511912 566884 511964
rect 580172 511912 580224 511964
rect 575020 485732 575072 485784
rect 579620 485732 579672 485784
rect 3332 463632 3384 463684
rect 4436 463632 4488 463684
rect 577504 419432 577556 419484
rect 579620 419432 579672 419484
rect 570696 405628 570748 405680
rect 579804 405628 579856 405680
rect 574928 379448 574980 379500
rect 579804 379448 579856 379500
rect 572076 353200 572128 353252
rect 580172 353200 580224 353252
rect 570604 325592 570656 325644
rect 580172 325592 580224 325644
rect 576308 313216 576360 313268
rect 580172 313216 580224 313268
rect 569500 299412 569552 299464
rect 580172 299412 580224 299464
rect 576216 273164 576268 273216
rect 580172 273164 580224 273216
rect 574836 259360 574888 259412
rect 579620 259360 579672 259412
rect 565360 245556 565412 245608
rect 580172 245556 580224 245608
rect 569316 233180 569368 233232
rect 580172 233180 580224 233232
rect 573548 219376 573600 219428
rect 580172 219376 580224 219428
rect 566740 206932 566792 206984
rect 579896 206932 579948 206984
rect 573456 179324 573508 179376
rect 579988 179324 580040 179376
rect 566556 166948 566608 167000
rect 580172 166948 580224 167000
rect 565176 139340 565228 139392
rect 580172 139340 580224 139392
rect 573364 126896 573416 126948
rect 580172 126896 580224 126948
rect 566648 113092 566700 113144
rect 579804 113092 579856 113144
rect 571984 100648 572036 100700
rect 580172 100648 580224 100700
rect 574744 86912 574796 86964
rect 580172 86912 580224 86964
rect 565268 73108 565320 73160
rect 580172 73108 580224 73160
rect 569408 60664 569460 60716
rect 580172 60664 580224 60716
rect 576124 46860 576176 46912
rect 580172 46860 580224 46912
rect 569224 33056 569276 33108
rect 580172 33056 580224 33108
rect 566464 20612 566516 20664
rect 579988 20612 580040 20664
rect 565084 6808 565136 6860
rect 580172 6808 580224 6860
rect 563704 3000 563756 3052
rect 583392 3000 583444 3052
rect 563520 2864 563572 2916
rect 572720 2864 572772 2916
rect 569868 2796 569920 2848
rect 576308 2796 576360 2848
rect 563520 1028 563572 1080
rect 1676 620 1728 672
rect 5356 620 5408 672
rect 6460 620 6512 672
rect 10048 620 10100 672
rect 572 552 624 604
rect 4344 552 4396 604
rect 5264 552 5316 604
rect 8852 552 8904 604
rect 7472 527 7524 536
rect 7472 493 7481 527
rect 7481 493 7515 527
rect 7515 493 7524 527
rect 7472 484 7524 493
rect 8576 484 8628 536
rect 11152 552 11204 604
rect 11520 620 11572 672
rect 19432 620 19484 672
rect 22376 620 22428 672
rect 12348 552 12400 604
rect 15568 552 15620 604
rect 21824 552 21876 604
rect 24860 620 24912 672
rect 25320 620 25372 672
rect 28080 620 28132 672
rect 28724 620 28776 672
rect 29184 620 29236 672
rect 31300 620 31352 672
rect 33784 620 33836 672
rect 34796 620 34848 672
rect 37280 620 37332 672
rect 38384 620 38436 672
rect 23020 552 23072 604
rect 25780 552 25832 604
rect 28816 552 28868 604
rect 3240 416 3292 468
rect 6644 416 6696 468
rect 12624 484 12676 536
rect 13268 484 13320 536
rect 16672 484 16724 536
rect 17408 484 17460 536
rect 20076 484 20128 536
rect 30104 552 30156 604
rect 32588 552 32640 604
rect 33600 552 33652 604
rect 36084 552 36136 604
rect 37188 552 37240 604
rect 40684 620 40736 672
rect 42800 620 42852 672
rect 46664 620 46716 672
rect 48504 620 48556 672
rect 48964 620 49016 672
rect 50804 620 50856 672
rect 53748 620 53800 672
rect 55404 620 55456 672
rect 64328 620 64380 672
rect 65616 620 65668 672
rect 66720 620 66772 672
rect 68008 620 68060 672
rect 69112 620 69164 672
rect 70584 620 70636 672
rect 133236 620 133288 672
rect 134156 620 134208 672
rect 136180 620 136232 672
rect 137652 620 137704 672
rect 138756 620 138808 672
rect 140044 620 140096 672
rect 151360 620 151412 672
rect 153016 620 153068 672
rect 153660 620 153712 672
rect 155408 620 155460 672
rect 162768 620 162820 672
rect 164884 620 164936 672
rect 40776 552 40828 604
rect 41880 552 41932 604
rect 43996 552 44048 604
rect 47860 552 47912 604
rect 49608 552 49660 604
rect 50160 552 50212 604
rect 51356 552 51408 604
rect 53012 552 53064 604
rect 54944 552 54996 604
rect 56416 552 56468 604
rect 60832 552 60884 604
rect 62120 552 62172 604
rect 65524 552 65576 604
rect 66812 552 66864 604
rect 70308 552 70360 604
rect 71228 552 71280 604
rect 76196 552 76248 604
rect 76932 552 76984 604
rect 77392 552 77444 604
rect 78036 552 78088 604
rect 78588 552 78640 604
rect 79140 552 79192 604
rect 79692 552 79744 604
rect 80336 552 80388 604
rect 80888 552 80940 604
rect 81440 552 81492 604
rect 82084 552 82136 604
rect 82728 552 82780 604
rect 121828 552 121880 604
rect 122288 552 122340 604
rect 124128 552 124180 604
rect 124680 552 124732 604
rect 125232 552 125284 604
rect 125876 552 125928 604
rect 126428 552 126480 604
rect 126980 552 127032 604
rect 127532 552 127584 604
rect 128176 552 128228 604
rect 128636 552 128688 604
rect 129372 552 129424 604
rect 133880 552 133932 604
rect 135260 552 135312 604
rect 136456 552 136508 604
rect 137560 552 137612 604
rect 138848 552 138900 604
rect 139952 552 140004 604
rect 141240 552 141292 604
rect 144552 552 144604 604
rect 145932 552 145984 604
rect 146852 552 146904 604
rect 148324 552 148376 604
rect 152556 552 152608 604
rect 154212 552 154264 604
rect 154764 552 154816 604
rect 156604 552 156656 604
rect 157064 552 157116 604
rect 158904 552 158956 604
rect 161572 552 161624 604
rect 163688 552 163740 604
rect 31668 484 31720 536
rect 33232 484 33284 536
rect 34980 484 35032 536
rect 14464 416 14516 468
rect 24400 416 24452 468
rect 26884 416 26936 468
rect 51908 484 51960 536
rect 63500 484 63552 536
rect 64512 484 64564 536
rect 67732 484 67784 536
rect 69388 484 69440 536
rect 134984 484 135036 536
rect 141056 484 141108 536
rect 142068 484 142120 536
rect 158168 484 158220 536
rect 159732 484 159784 536
rect 39856 416 39908 468
rect 163412 416 163464 468
rect 166080 620 166132 672
rect 167092 620 167144 672
rect 169576 620 169628 672
rect 180892 620 180944 672
rect 183744 620 183796 672
rect 190000 620 190052 672
rect 193220 620 193272 672
rect 194324 620 194376 672
rect 197912 620 197964 672
rect 213828 620 213880 672
rect 165988 552 166040 604
rect 168380 552 168432 604
rect 170680 552 170732 604
rect 173164 552 173216 604
rect 179788 552 179840 604
rect 182548 552 182600 604
rect 183192 552 183244 604
rect 186136 552 186188 604
rect 188804 552 188856 604
rect 192300 552 192352 604
rect 195612 552 195664 604
rect 196900 552 196952 604
rect 205732 552 205784 604
rect 209780 552 209832 604
rect 210424 552 210476 604
rect 187700 484 187752 536
rect 191012 484 191064 536
rect 192208 484 192260 536
rect 192944 484 192996 536
rect 211620 552 211672 604
rect 215668 620 215720 672
rect 217968 620 218020 672
rect 218428 620 218480 672
rect 222752 620 222804 672
rect 214472 552 214524 604
rect 220176 552 220228 604
rect 220452 552 220504 604
rect 221832 552 221884 604
rect 226340 620 226392 672
rect 223948 552 224000 604
rect 226156 552 226208 604
rect 231032 620 231084 672
rect 219532 484 219584 536
rect 224776 484 224828 536
rect 229836 552 229888 604
rect 229652 484 229704 536
rect 234620 620 234672 672
rect 235448 620 235500 672
rect 237748 620 237800 672
rect 242900 620 242952 672
rect 247960 620 248012 672
rect 253480 620 253532 672
rect 257068 620 257120 672
rect 257252 620 257304 672
rect 258264 620 258316 672
rect 231860 552 231912 604
rect 237012 552 237064 604
rect 238116 552 238168 604
rect 233148 484 233200 536
rect 212724 416 212776 468
rect 216588 416 216640 468
rect 234344 416 234396 468
rect 239312 552 239364 604
rect 240508 595 240560 604
rect 240508 561 240517 595
rect 240517 561 240551 595
rect 240551 561 240560 595
rect 240508 552 240560 561
rect 241152 552 241204 604
rect 246028 552 246080 604
rect 249984 552 250036 604
rect 251180 552 251232 604
rect 252376 552 252428 604
rect 253388 552 253440 604
rect 254584 552 254636 604
rect 260656 620 260708 672
rect 262680 620 262732 672
rect 268844 620 268896 672
rect 272892 620 272944 672
rect 285404 620 285456 672
rect 244556 484 244608 536
rect 239956 416 240008 468
rect 244924 416 244976 468
rect 245660 416 245712 468
rect 14556 348 14608 400
rect 17868 348 17920 400
rect 39304 348 39356 400
rect 42156 348 42208 400
rect 42892 348 42944 400
rect 45100 348 45152 400
rect 71320 348 71372 400
rect 72332 348 72384 400
rect 72424 348 72476 400
rect 73528 348 73580 400
rect 73620 348 73672 400
rect 74632 348 74684 400
rect 130936 348 130988 400
rect 131948 348 132000 400
rect 132040 348 132092 400
rect 133144 348 133196 400
rect 160468 348 160520 400
rect 162676 348 162728 400
rect 220176 348 220228 400
rect 225328 348 225380 400
rect 246764 348 246816 400
rect 259460 552 259512 604
rect 260472 552 260524 604
rect 266544 552 266596 604
rect 270040 552 270092 604
rect 274088 552 274140 604
rect 263692 484 263744 536
rect 270500 484 270552 536
rect 276756 484 276808 536
rect 279516 552 279568 604
rect 284300 552 284352 604
rect 257988 416 258040 468
rect 259276 416 259328 468
rect 264980 416 265032 468
rect 268384 416 268436 468
rect 274548 416 274600 468
rect 277492 416 277544 468
rect 281540 484 281592 536
rect 288992 620 289044 672
rect 291108 620 291160 672
rect 293408 620 293460 672
rect 298468 620 298520 672
rect 300768 620 300820 672
rect 301320 620 301372 672
rect 288808 552 288860 604
rect 296076 552 296128 604
rect 303160 552 303212 604
rect 287612 484 287664 536
rect 293868 484 293920 536
rect 295616 484 295668 536
rect 304724 620 304776 672
rect 303620 552 303672 604
rect 307944 663 307996 672
rect 307944 629 307953 663
rect 307953 629 307987 663
rect 307987 629 307996 663
rect 307944 620 307996 629
rect 309968 620 310020 672
rect 309048 552 309100 604
rect 310244 552 310296 604
rect 311440 595 311492 604
rect 311440 561 311449 595
rect 311449 561 311483 595
rect 311483 561 311492 595
rect 311440 552 311492 561
rect 312636 595 312688 604
rect 312636 561 312645 595
rect 312645 561 312679 595
rect 312679 561 312688 595
rect 312636 552 312688 561
rect 318524 620 318576 672
rect 318708 620 318760 672
rect 319536 620 319588 672
rect 315948 552 316000 604
rect 280896 416 280948 468
rect 284116 416 284168 468
rect 291200 416 291252 468
rect 300216 416 300268 468
rect 263140 348 263192 400
rect 269488 348 269540 400
rect 276204 348 276256 400
rect 278596 348 278648 400
rect 294512 348 294564 400
rect 301780 348 301832 400
rect 302424 348 302476 400
rect 316040 484 316092 536
rect 317144 552 317196 604
rect 325608 552 325660 604
rect 326804 620 326856 672
rect 328460 620 328512 672
rect 331956 620 332008 672
rect 328000 552 328052 604
rect 330392 552 330444 604
rect 242256 280 242308 332
rect 247316 280 247368 332
rect 250904 280 250956 332
rect 256884 280 256936 332
rect 262772 280 262824 332
rect 271788 280 271840 332
rect 278504 280 278556 332
rect 297916 280 297968 332
rect 305736 280 305788 332
rect 308772 280 308824 332
rect 316592 416 316644 468
rect 318340 416 318392 468
rect 318708 416 318760 468
rect 321560 484 321612 536
rect 337476 620 337528 672
rect 342168 620 342220 672
rect 338672 595 338724 604
rect 338672 561 338681 595
rect 338681 561 338715 595
rect 338715 561 338724 595
rect 338672 552 338724 561
rect 339868 552 339920 604
rect 340972 552 341024 604
rect 342076 552 342128 604
rect 348240 620 348292 672
rect 349068 620 349120 672
rect 351644 620 351696 672
rect 352472 620 352524 672
rect 361948 620 362000 672
rect 369584 620 369636 672
rect 370412 663 370464 672
rect 370412 629 370421 663
rect 370421 629 370455 663
rect 370455 629 370464 663
rect 370412 620 370464 629
rect 370688 620 370740 672
rect 371608 620 371660 672
rect 375196 663 375248 672
rect 375196 629 375205 663
rect 375205 629 375239 663
rect 375239 629 375248 663
rect 375196 620 375248 629
rect 377404 620 377456 672
rect 344468 552 344520 604
rect 354036 552 354088 604
rect 343180 484 343232 536
rect 351828 484 351880 536
rect 324228 416 324280 468
rect 325148 416 325200 468
rect 333612 416 333664 468
rect 346768 416 346820 468
rect 356336 552 356388 604
rect 358728 595 358780 604
rect 358728 561 358737 595
rect 358737 561 358771 595
rect 358771 561 358780 595
rect 358728 552 358780 561
rect 354680 484 354732 536
rect 364800 552 364852 604
rect 368204 552 368256 604
rect 369308 552 369360 604
rect 379980 552 380032 604
rect 381176 552 381228 604
rect 382372 620 382424 672
rect 385960 620 386012 672
rect 388812 663 388864 672
rect 388812 629 388821 663
rect 388821 629 388855 663
rect 388855 629 388864 663
rect 388812 620 388864 629
rect 388260 552 388312 604
rect 359280 484 359332 536
rect 362684 484 362736 536
rect 373080 484 373132 536
rect 356980 416 357032 468
rect 311072 348 311124 400
rect 319904 348 319956 400
rect 327448 348 327500 400
rect 336464 348 336516 400
rect 349068 348 349120 400
rect 360384 416 360436 468
rect 366732 416 366784 468
rect 377404 484 377456 536
rect 385408 484 385460 536
rect 396540 620 396592 672
rect 391020 552 391072 604
rect 400036 663 400088 672
rect 400036 629 400045 663
rect 400045 629 400079 663
rect 400079 629 400088 663
rect 400036 620 400088 629
rect 402520 620 402572 672
rect 403440 620 403492 672
rect 409236 663 409288 672
rect 397736 595 397788 604
rect 397736 561 397745 595
rect 397745 561 397779 595
rect 397779 561 397788 595
rect 397736 552 397788 561
rect 398840 552 398892 604
rect 400220 595 400272 604
rect 400220 561 400229 595
rect 400229 561 400263 595
rect 400263 561 400272 595
rect 400220 552 400272 561
rect 400312 552 400364 604
rect 403532 552 403584 604
rect 389824 484 389876 536
rect 409236 629 409245 663
rect 409245 629 409279 663
rect 409279 629 409288 663
rect 409236 620 409288 629
rect 410800 620 410852 672
rect 404728 595 404780 604
rect 404728 561 404737 595
rect 404737 561 404771 595
rect 404771 561 404780 595
rect 404728 552 404780 561
rect 404820 595 404872 604
rect 404820 561 404829 595
rect 404829 561 404863 595
rect 404863 561 404872 595
rect 404820 552 404872 561
rect 405648 552 405700 604
rect 412640 595 412692 604
rect 412640 561 412649 595
rect 412649 561 412683 595
rect 412683 561 412692 595
rect 412640 552 412692 561
rect 413744 595 413796 604
rect 413744 561 413753 595
rect 413753 561 413787 595
rect 413787 561 413796 595
rect 413744 552 413796 561
rect 414296 595 414348 604
rect 414296 561 414305 595
rect 414305 561 414339 595
rect 414339 561 414348 595
rect 414296 552 414348 561
rect 415492 595 415544 604
rect 415492 561 415501 595
rect 415501 561 415535 595
rect 415535 561 415544 595
rect 415492 552 415544 561
rect 416688 620 416740 672
rect 418344 663 418396 672
rect 418344 629 418353 663
rect 418353 629 418387 663
rect 418387 629 418396 663
rect 418344 620 418396 629
rect 421012 663 421064 672
rect 421012 629 421021 663
rect 421021 629 421055 663
rect 421055 629 421064 663
rect 421012 620 421064 629
rect 421104 620 421156 672
rect 423496 620 423548 672
rect 425520 663 425572 672
rect 425520 629 425529 663
rect 425529 629 425563 663
rect 425563 629 425572 663
rect 425520 620 425572 629
rect 425612 620 425664 672
rect 430856 620 430908 672
rect 431868 663 431920 672
rect 431868 629 431877 663
rect 431877 629 431911 663
rect 431911 629 431920 663
rect 431868 620 431920 629
rect 432052 663 432104 672
rect 432052 629 432061 663
rect 432061 629 432095 663
rect 432095 629 432104 663
rect 432052 620 432104 629
rect 417884 552 417936 604
rect 423772 552 423824 604
rect 427268 552 427320 604
rect 428372 595 428424 604
rect 428372 561 428381 595
rect 428381 561 428415 595
rect 428415 561 428424 595
rect 428372 552 428424 561
rect 429476 552 429528 604
rect 433248 552 433300 604
rect 434720 552 434772 604
rect 435548 552 435600 604
rect 436468 663 436520 672
rect 436468 629 436477 663
rect 436477 629 436511 663
rect 436511 629 436520 663
rect 436468 620 436520 629
rect 436744 620 436796 672
rect 437480 620 437532 672
rect 439872 663 439924 672
rect 439136 552 439188 604
rect 439872 629 439881 663
rect 439881 629 439915 663
rect 439915 629 439924 663
rect 439872 620 439924 629
rect 449992 620 450044 672
rect 453580 663 453632 672
rect 453580 629 453589 663
rect 453589 629 453623 663
rect 453623 629 453632 663
rect 453580 620 453632 629
rect 454224 663 454276 672
rect 454224 629 454233 663
rect 454233 629 454267 663
rect 454267 629 454276 663
rect 454224 620 454276 629
rect 454500 663 454552 672
rect 454500 629 454509 663
rect 454509 629 454543 663
rect 454543 629 454552 663
rect 454500 620 454552 629
rect 456892 620 456944 672
rect 460388 620 460440 672
rect 460664 620 460716 672
rect 462136 663 462188 672
rect 462136 629 462145 663
rect 462145 629 462179 663
rect 462179 629 462188 663
rect 462136 620 462188 629
rect 466368 663 466420 672
rect 466368 629 466377 663
rect 466377 629 466411 663
rect 466411 629 466420 663
rect 466368 620 466420 629
rect 467196 663 467248 672
rect 467196 629 467205 663
rect 467205 629 467239 663
rect 467239 629 467248 663
rect 467196 620 467248 629
rect 468300 663 468352 672
rect 468300 629 468309 663
rect 468309 629 468343 663
rect 468343 629 468352 663
rect 468300 620 468352 629
rect 468668 620 468720 672
rect 441528 552 441580 604
rect 442632 595 442684 604
rect 442632 561 442641 595
rect 442641 561 442675 595
rect 442675 561 442684 595
rect 442632 552 442684 561
rect 444472 595 444524 604
rect 444472 561 444481 595
rect 444481 561 444515 595
rect 444515 561 444524 595
rect 444472 552 444524 561
rect 445024 595 445076 604
rect 445024 561 445033 595
rect 445033 561 445067 595
rect 445067 561 445076 595
rect 445024 552 445076 561
rect 373908 416 373960 468
rect 384580 416 384632 468
rect 393320 459 393372 468
rect 393320 425 393329 459
rect 393329 425 393363 459
rect 393363 425 393372 459
rect 393320 416 393372 425
rect 395620 416 395672 468
rect 408224 484 408276 536
rect 410340 484 410392 536
rect 422760 484 422812 536
rect 405740 416 405792 468
rect 408132 416 408184 468
rect 419908 416 419960 468
rect 420552 416 420604 468
rect 438768 484 438820 536
rect 430672 416 430724 468
rect 367284 348 367336 400
rect 372436 348 372488 400
rect 312452 280 312504 332
rect 320732 280 320784 332
rect 333152 280 333204 332
rect 340604 280 340656 332
rect 347780 280 347832 332
rect 351276 280 351328 332
rect 360844 280 360896 332
rect 363788 280 363840 332
rect 374276 280 374328 332
rect 378600 348 378652 400
rect 389180 348 389232 400
rect 389916 348 389968 400
rect 393780 348 393832 400
rect 383292 280 383344 332
rect 386972 280 387024 332
rect 394424 280 394476 332
rect 233240 212 233292 264
rect 236552 212 236604 264
rect 241428 212 241480 264
rect 255688 212 255740 264
rect 261484 212 261536 264
rect 261576 212 261628 264
rect 267556 212 267608 264
rect 280436 212 280488 264
rect 287060 212 287112 264
rect 296812 212 296864 264
rect 303988 212 304040 264
rect 307668 212 307720 264
rect 313648 212 313700 264
rect 321836 212 321888 264
rect 322848 212 322900 264
rect 331220 212 331272 264
rect 337200 212 337252 264
rect 16304 76 16356 128
rect 18972 76 19024 128
rect 45744 76 45796 128
rect 47400 76 47452 128
rect 129832 76 129884 128
rect 130292 76 130344 128
rect 155960 76 156012 128
rect 157524 76 157576 128
rect 159364 76 159416 128
rect 161480 76 161532 128
rect 184296 76 184348 128
rect 186964 144 187016 196
rect 228548 144 228600 196
rect 264888 144 264940 196
rect 271052 144 271104 196
rect 282920 144 282972 196
rect 290004 144 290056 196
rect 292212 144 292264 196
rect 299388 144 299440 196
rect 324044 144 324096 196
rect 332508 144 332560 196
rect 338304 144 338356 196
rect 345572 212 345624 264
rect 354956 212 355008 264
rect 355876 212 355928 264
rect 365996 212 366048 264
rect 382004 212 382056 264
rect 393228 212 393280 264
rect 393964 212 394016 264
rect 401140 348 401192 400
rect 397460 212 397512 264
rect 411720 348 411772 400
rect 424692 348 424744 400
rect 433064 416 433116 468
rect 446220 552 446272 604
rect 446680 595 446732 604
rect 446680 561 446689 595
rect 446689 561 446723 595
rect 446723 561 446732 595
rect 446680 552 446732 561
rect 447876 552 447928 604
rect 458088 595 458140 604
rect 458088 561 458097 595
rect 458097 561 458131 595
rect 458131 561 458140 595
rect 458088 552 458140 561
rect 461492 595 461544 604
rect 461492 561 461501 595
rect 461501 561 461535 595
rect 461535 561 461544 595
rect 461492 552 461544 561
rect 463608 552 463660 604
rect 477868 620 477920 672
rect 482928 620 482980 672
rect 483020 663 483072 672
rect 483020 629 483029 663
rect 483029 629 483063 663
rect 483063 629 483072 663
rect 484032 663 484084 672
rect 483020 620 483072 629
rect 484032 629 484041 663
rect 484041 629 484075 663
rect 484075 629 484084 663
rect 484032 620 484084 629
rect 486608 663 486660 672
rect 486608 629 486617 663
rect 486617 629 486651 663
rect 486651 629 486660 663
rect 486608 620 486660 629
rect 487436 663 487488 672
rect 487436 629 487445 663
rect 487445 629 487479 663
rect 487479 629 487488 663
rect 487436 620 487488 629
rect 487620 663 487672 672
rect 487620 629 487629 663
rect 487629 629 487663 663
rect 487663 629 487672 663
rect 487620 620 487672 629
rect 488264 663 488316 672
rect 488264 629 488273 663
rect 488273 629 488307 663
rect 488307 629 488316 663
rect 488264 620 488316 629
rect 492680 620 492732 672
rect 496820 663 496872 672
rect 496820 629 496829 663
rect 496829 629 496863 663
rect 496863 629 496872 663
rect 496820 620 496872 629
rect 498200 620 498252 672
rect 498936 663 498988 672
rect 498936 629 498945 663
rect 498945 629 498979 663
rect 498979 629 498988 663
rect 498936 620 498988 629
rect 502340 663 502392 672
rect 502340 629 502349 663
rect 502349 629 502383 663
rect 502383 629 502392 663
rect 502340 620 502392 629
rect 502984 663 503036 672
rect 502984 629 502993 663
rect 502993 629 503027 663
rect 503027 629 503036 663
rect 502984 620 503036 629
rect 505744 663 505796 672
rect 505744 629 505753 663
rect 505753 629 505787 663
rect 505787 629 505796 663
rect 505744 620 505796 629
rect 507860 663 507912 672
rect 507860 629 507869 663
rect 507869 629 507903 663
rect 507903 629 507912 663
rect 509884 663 509936 672
rect 507860 620 507912 629
rect 509884 629 509893 663
rect 509893 629 509927 663
rect 509927 629 509936 663
rect 509884 620 509936 629
rect 510988 620 511040 672
rect 470600 595 470652 604
rect 470600 561 470609 595
rect 470609 561 470643 595
rect 470643 561 470652 595
rect 470600 552 470652 561
rect 471704 595 471756 604
rect 471704 561 471713 595
rect 471713 561 471747 595
rect 471747 561 471756 595
rect 471704 552 471756 561
rect 472256 595 472308 604
rect 472256 561 472265 595
rect 472265 561 472299 595
rect 472299 561 472308 595
rect 472256 552 472308 561
rect 474556 595 474608 604
rect 474556 561 474565 595
rect 474565 561 474599 595
rect 474599 561 474608 595
rect 474556 552 474608 561
rect 475752 595 475804 604
rect 475752 561 475761 595
rect 475761 561 475795 595
rect 475795 561 475804 595
rect 475752 552 475804 561
rect 476948 595 477000 604
rect 476948 561 476957 595
rect 476957 561 476991 595
rect 476991 561 477000 595
rect 476948 552 477000 561
rect 481732 595 481784 604
rect 481732 561 481741 595
rect 481741 561 481775 595
rect 481775 561 481784 595
rect 481732 552 481784 561
rect 485136 552 485188 604
rect 485412 552 485464 604
rect 486332 552 486384 604
rect 490932 595 490984 604
rect 406936 280 406988 332
rect 185492 76 185544 128
rect 188252 76 188304 128
rect 227352 76 227404 128
rect 232044 76 232096 128
rect 252008 76 252060 128
rect 257252 76 257304 128
rect 266084 76 266136 128
rect 272156 76 272208 128
rect 286416 76 286468 128
rect 291568 76 291620 128
rect 299020 76 299072 128
rect 306932 76 306984 128
rect 320640 76 320692 128
rect 329012 76 329064 128
rect 329748 76 329800 128
rect 345940 144 345992 196
rect 347412 144 347464 196
rect 357348 144 357400 196
rect 358084 144 358136 196
rect 347688 76 347740 128
rect 350172 76 350224 128
rect 359740 76 359792 128
rect 361488 144 361540 196
rect 371976 144 372028 196
rect 380808 144 380860 196
rect 385776 144 385828 196
rect 386512 144 386564 196
rect 412916 212 412968 264
rect 416044 280 416096 332
rect 428648 280 428700 332
rect 443644 348 443696 400
rect 437572 280 437624 332
rect 442172 280 442224 332
rect 455880 484 455932 536
rect 459008 484 459060 536
rect 450636 416 450688 468
rect 459560 416 459612 468
rect 460204 416 460256 468
rect 449624 348 449676 400
rect 452292 391 452344 400
rect 452292 357 452301 391
rect 452301 357 452335 391
rect 452335 357 452344 391
rect 452292 348 452344 357
rect 452384 348 452436 400
rect 451280 280 451332 332
rect 457904 348 457956 400
rect 477408 484 477460 536
rect 489276 484 489328 536
rect 490932 561 490941 595
rect 490941 561 490975 595
rect 490975 561 490984 595
rect 490932 552 490984 561
rect 491116 595 491168 604
rect 491116 561 491125 595
rect 491125 561 491159 595
rect 491159 561 491168 595
rect 491116 552 491168 561
rect 501788 552 501840 604
rect 510252 552 510304 604
rect 496728 484 496780 536
rect 512460 620 512512 672
rect 514392 663 514444 672
rect 514392 629 514401 663
rect 514401 629 514435 663
rect 514435 629 514444 663
rect 514392 620 514444 629
rect 515956 620 516008 672
rect 516968 663 517020 672
rect 516968 629 516977 663
rect 516977 629 517011 663
rect 517011 629 517020 663
rect 516968 620 517020 629
rect 518256 663 518308 672
rect 518256 629 518265 663
rect 518265 629 518299 663
rect 518299 629 518308 663
rect 518256 620 518308 629
rect 518348 663 518400 672
rect 518348 629 518357 663
rect 518357 629 518391 663
rect 518391 629 518400 663
rect 518348 620 518400 629
rect 519452 620 519504 672
rect 520740 663 520792 672
rect 513564 552 513616 604
rect 519544 552 519596 604
rect 520740 629 520749 663
rect 520749 629 520783 663
rect 520783 629 520792 663
rect 520740 620 520792 629
rect 521936 663 521988 672
rect 521936 629 521945 663
rect 521945 629 521979 663
rect 521979 629 521988 663
rect 521936 620 521988 629
rect 522856 620 522908 672
rect 569868 960 569920 1012
rect 569132 892 569184 944
rect 523500 620 523552 672
rect 523040 595 523092 604
rect 523040 561 523049 595
rect 523049 561 523083 595
rect 523083 561 523092 595
rect 523040 552 523092 561
rect 530124 620 530176 672
rect 531136 663 531188 672
rect 531136 629 531145 663
rect 531145 629 531179 663
rect 531179 629 531188 663
rect 531136 620 531188 629
rect 531320 663 531372 672
rect 531320 629 531329 663
rect 531329 629 531363 663
rect 531363 629 531372 663
rect 531320 620 531372 629
rect 531872 620 531924 672
rect 548340 620 548392 672
rect 548984 620 549036 672
rect 566832 824 566884 876
rect 568028 756 568080 808
rect 570328 688 570380 740
rect 551100 663 551152 672
rect 551100 629 551109 663
rect 551109 629 551143 663
rect 551143 629 551152 663
rect 551100 620 551152 629
rect 524236 595 524288 604
rect 524236 561 524245 595
rect 524245 561 524279 595
rect 524279 561 524288 595
rect 524236 552 524288 561
rect 525064 552 525116 604
rect 526260 552 526312 604
rect 538772 595 538824 604
rect 538772 561 538781 595
rect 538781 561 538815 595
rect 538815 561 538824 595
rect 538772 552 538824 561
rect 540796 595 540848 604
rect 540796 561 540805 595
rect 540805 561 540839 595
rect 540839 561 540848 595
rect 540796 552 540848 561
rect 541992 595 542044 604
rect 541992 561 542001 595
rect 542001 561 542035 595
rect 542035 561 542044 595
rect 541992 552 542044 561
rect 543096 552 543148 604
rect 543372 595 543424 604
rect 543372 561 543381 595
rect 543381 561 543415 595
rect 543415 561 543424 595
rect 544200 595 544252 604
rect 543372 552 543424 561
rect 544200 561 544209 595
rect 544209 561 544243 595
rect 544243 561 544252 595
rect 544200 552 544252 561
rect 544384 595 544436 604
rect 544384 561 544393 595
rect 544393 561 544427 595
rect 544427 561 544436 595
rect 544384 552 544436 561
rect 545120 595 545172 604
rect 545120 561 545129 595
rect 545129 561 545163 595
rect 545163 561 545172 595
rect 545120 552 545172 561
rect 545488 595 545540 604
rect 545488 561 545497 595
rect 545497 561 545531 595
rect 545531 561 545540 595
rect 545488 552 545540 561
rect 552388 620 552440 672
rect 565636 620 565688 672
rect 469220 416 469272 468
rect 495348 416 495400 468
rect 504640 459 504692 468
rect 504640 425 504649 459
rect 504649 425 504683 459
rect 504683 425 504692 459
rect 504640 416 504692 425
rect 506204 459 506256 468
rect 506204 425 506213 459
rect 506213 425 506247 459
rect 506247 425 506256 459
rect 506204 416 506256 425
rect 506940 416 506992 468
rect 509700 416 509752 468
rect 511448 416 511500 468
rect 513288 416 513340 468
rect 514944 459 514996 468
rect 514944 425 514953 459
rect 514953 425 514987 459
rect 514987 425 514996 459
rect 514944 416 514996 425
rect 527548 416 527600 468
rect 533068 484 533120 536
rect 539784 527 539836 536
rect 539784 493 539793 527
rect 539793 493 539827 527
rect 539827 493 539836 527
rect 539784 484 539836 493
rect 560852 552 560904 604
rect 562048 595 562100 604
rect 562048 561 562057 595
rect 562057 561 562091 595
rect 562091 561 562100 595
rect 562048 552 562100 561
rect 563244 595 563296 604
rect 563244 561 563253 595
rect 563253 561 563287 595
rect 563287 561 563296 595
rect 563244 552 563296 561
rect 573916 552 573968 604
rect 575112 552 575164 604
rect 549260 527 549312 536
rect 549260 493 549269 527
rect 549269 493 549303 527
rect 549303 493 549312 527
rect 549260 484 549312 493
rect 550088 484 550140 536
rect 554596 527 554648 536
rect 554596 493 554605 527
rect 554605 493 554639 527
rect 554639 493 554648 527
rect 554596 484 554648 493
rect 555792 484 555844 536
rect 535828 416 535880 468
rect 536472 416 536524 468
rect 553492 416 553544 468
rect 556896 416 556948 468
rect 418804 212 418856 264
rect 421748 212 421800 264
rect 434076 212 434128 264
rect 443276 212 443328 264
rect 465356 280 465408 332
rect 473268 348 473320 400
rect 472808 280 472860 332
rect 487804 348 487856 400
rect 492588 348 492640 400
rect 494428 348 494480 400
rect 503996 391 504048 400
rect 503996 357 504005 391
rect 504005 357 504039 391
rect 504039 357 504048 391
rect 503996 348 504048 357
rect 509240 348 509292 400
rect 525248 348 525300 400
rect 527180 348 527232 400
rect 547696 348 547748 400
rect 553308 348 553360 400
rect 571156 348 571208 400
rect 483756 280 483808 332
rect 495532 280 495584 332
rect 497832 280 497884 332
rect 520372 280 520424 332
rect 536932 280 536984 332
rect 541716 280 541768 332
rect 555884 280 555936 332
rect 558000 323 558052 332
rect 558000 289 558009 323
rect 558009 289 558043 323
rect 558043 289 558052 323
rect 558000 280 558052 289
rect 559012 280 559064 332
rect 576768 280 576820 332
rect 463056 212 463108 264
rect 464896 212 464948 264
rect 409420 144 409472 196
rect 411536 144 411588 196
rect 422392 144 422444 196
rect 434720 144 434772 196
rect 435364 144 435416 196
rect 448244 144 448296 196
rect 448980 144 449032 196
rect 462412 144 462464 196
rect 367836 76 367888 128
rect 378692 76 378744 128
rect 379520 76 379572 128
rect 390284 76 390336 128
rect 395528 76 395580 128
rect 396264 76 396316 128
rect 402336 76 402388 128
rect 419448 76 419500 128
rect 434260 76 434312 128
rect 447140 76 447192 128
rect 453488 119 453540 128
rect 453488 85 453497 119
rect 453497 85 453531 119
rect 453531 85 453540 119
rect 453488 76 453540 85
rect 456524 76 456576 128
rect 467840 144 467892 196
rect 478512 212 478564 264
rect 490288 212 490340 264
rect 492128 212 492180 264
rect 502708 212 502760 264
rect 503536 212 503588 264
rect 479524 144 479576 196
rect 480812 144 480864 196
rect 489736 144 489788 196
rect 505192 144 505244 196
rect 506940 144 506992 196
rect 512184 144 512236 196
rect 528836 212 528888 264
rect 529664 212 529716 264
rect 546500 212 546552 264
rect 562600 212 562652 264
rect 581828 212 581880 264
rect 521568 144 521620 196
rect 538036 144 538088 196
rect 539876 144 539928 196
rect 557172 144 557224 196
rect 560208 144 560260 196
rect 578332 144 578384 196
rect 466000 76 466052 128
rect 480720 76 480772 128
rect 481456 76 481508 128
rect 496820 76 496872 128
rect 500132 76 500184 128
rect 515588 76 515640 128
rect 532332 76 532384 128
rect 534540 119 534592 128
rect 534540 85 534549 119
rect 534549 85 534583 119
rect 534583 85 534592 119
rect 534540 76 534592 85
rect 550456 76 550508 128
rect 44088 8 44140 60
rect 46204 8 46256 60
rect 215024 8 215076 60
rect 219440 8 219492 60
rect 289820 8 289872 60
rect 296996 8 297048 60
rect 314752 8 314804 60
rect 322848 8 322900 60
rect 330852 8 330904 60
rect 339500 8 339552 60
rect 348240 8 348292 60
rect 353576 8 353628 60
rect 363696 8 363748 60
rect 376300 8 376352 60
rect 386788 8 386840 60
rect 387616 8 387668 60
rect 399116 8 399168 60
rect 407028 8 407080 60
rect 414940 8 414992 60
rect 426992 8 427044 60
rect 440148 8 440200 60
rect 441068 8 441120 60
rect 455328 8 455380 60
rect 469588 8 469640 60
rect 476212 8 476264 60
rect 493324 8 493376 60
rect 508596 8 508648 60
rect 526260 8 526312 60
rect 528468 8 528520 60
rect 546500 8 546552 60
rect 564624 76 564676 128
rect 561404 8 561456 60
rect 580724 8 580776 60
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 235356 703588 235408 703594
rect 235356 703530 235408 703536
rect 242440 703588 242492 703594
rect 242440 703530 242492 703536
rect 1492 703384 1544 703390
rect 1492 703326 1544 703332
rect 756 702840 808 702846
rect 756 702782 808 702788
rect 388 702704 440 702710
rect 388 702646 440 702652
rect 296 702636 348 702642
rect 296 702578 348 702584
rect 112 702568 164 702574
rect 112 702510 164 702516
rect 18 702128 74 702137
rect 18 702063 74 702072
rect 32 19961 60 702063
rect 124 71913 152 702510
rect 204 697672 256 697678
rect 204 697614 256 697620
rect 216 111217 244 697614
rect 308 171134 336 702578
rect 400 209774 428 702646
rect 572 701140 624 701146
rect 572 701082 624 701088
rect 480 697740 532 697746
rect 480 697682 532 697688
rect 492 214962 520 697682
rect 584 254153 612 701082
rect 662 700224 718 700233
rect 662 700159 718 700168
rect 676 397497 704 700159
rect 768 449585 796 702782
rect 1308 701820 1360 701826
rect 1308 701762 1360 701768
rect 938 700632 994 700641
rect 938 700567 994 700576
rect 848 699032 900 699038
rect 848 698974 900 698980
rect 860 553897 888 698974
rect 952 606121 980 700567
rect 1320 619614 1348 701762
rect 1504 684321 1532 703326
rect 1584 703248 1636 703254
rect 1584 703190 1636 703196
rect 1490 684312 1546 684321
rect 1490 684247 1546 684256
rect 1596 632097 1624 703190
rect 1676 703112 1728 703118
rect 1676 703054 1728 703060
rect 1582 632088 1638 632097
rect 1582 632023 1638 632032
rect 1308 619608 1360 619614
rect 1308 619550 1360 619556
rect 938 606112 994 606121
rect 938 606047 994 606056
rect 1688 580009 1716 703054
rect 1860 702976 1912 702982
rect 1860 702918 1912 702924
rect 1766 698184 1822 698193
rect 1766 698119 1822 698128
rect 1674 580000 1730 580009
rect 1674 579935 1730 579944
rect 846 553888 902 553897
rect 846 553823 902 553832
rect 1780 475697 1808 698119
rect 1872 527921 1900 702918
rect 2320 702772 2372 702778
rect 2320 702714 2372 702720
rect 2226 701448 2282 701457
rect 2226 701383 2282 701392
rect 2042 701312 2098 701321
rect 2042 701247 2098 701256
rect 1950 697912 2006 697921
rect 1950 697847 2006 697856
rect 1858 527912 1914 527921
rect 1858 527847 1914 527856
rect 1766 475688 1822 475697
rect 1766 475623 1822 475632
rect 754 449576 810 449585
rect 754 449511 810 449520
rect 1964 423609 1992 697847
rect 1950 423600 2006 423609
rect 1950 423535 2006 423544
rect 662 397488 718 397497
rect 662 397423 718 397432
rect 570 254144 626 254153
rect 570 254079 626 254088
rect 570 214976 626 214985
rect 492 214934 570 214962
rect 570 214911 626 214920
rect 400 209746 612 209774
rect 584 188873 612 209746
rect 570 188864 626 188873
rect 570 188799 626 188808
rect 308 171106 612 171134
rect 584 162897 612 171106
rect 570 162888 626 162897
rect 570 162823 626 162832
rect 202 111208 258 111217
rect 202 111143 258 111152
rect 110 71904 166 71913
rect 110 71839 166 71848
rect 18 19952 74 19961
rect 18 19887 74 19896
rect 2056 6497 2084 701247
rect 2134 699816 2190 699825
rect 2134 699751 2190 699760
rect 2148 32473 2176 699751
rect 2240 58585 2268 701383
rect 2332 267209 2360 702714
rect 4250 701856 4306 701865
rect 4250 701791 4306 701800
rect 2596 701548 2648 701554
rect 2596 701490 2648 701496
rect 2412 697808 2464 697814
rect 2412 697750 2464 697756
rect 2424 319297 2452 697750
rect 2502 697640 2558 697649
rect 2502 697575 2558 697584
rect 2516 345409 2544 697575
rect 2608 358465 2636 701490
rect 3884 700528 3936 700534
rect 2962 700496 3018 700505
rect 3884 700470 3936 700476
rect 2962 700431 3018 700440
rect 3700 700460 3752 700466
rect 2686 697776 2742 697785
rect 2686 697711 2742 697720
rect 2700 371385 2728 697711
rect 2780 619608 2832 619614
rect 2780 619550 2832 619556
rect 2792 514865 2820 619550
rect 2976 566953 3004 700431
rect 3700 700402 3752 700408
rect 3146 700360 3202 700369
rect 3146 700295 3202 700304
rect 3056 699644 3108 699650
rect 3056 699586 3108 699592
rect 3068 658209 3096 699586
rect 3054 658200 3110 658209
rect 3054 658135 3110 658144
rect 2962 566944 3018 566953
rect 2962 566879 3018 566888
rect 2778 514856 2834 514865
rect 2778 514791 2834 514800
rect 3160 462641 3188 700295
rect 3606 699952 3662 699961
rect 3606 699887 3662 699896
rect 3240 699780 3292 699786
rect 3240 699722 3292 699728
rect 3252 671265 3280 699722
rect 3516 699372 3568 699378
rect 3516 699314 3568 699320
rect 3422 699136 3478 699145
rect 3422 699071 3478 699080
rect 3330 698048 3386 698057
rect 3330 697983 3386 697992
rect 3238 671256 3294 671265
rect 3238 671191 3294 671200
rect 3240 661088 3292 661094
rect 3240 661030 3292 661036
rect 3146 462632 3202 462641
rect 3146 462567 3202 462576
rect 3252 410553 3280 661030
rect 3344 501809 3372 697983
rect 3330 501800 3386 501809
rect 3330 501735 3386 501744
rect 3332 463684 3384 463690
rect 3332 463626 3384 463632
rect 3238 410544 3294 410553
rect 3238 410479 3294 410488
rect 2686 371376 2742 371385
rect 2686 371311 2742 371320
rect 2594 358456 2650 358465
rect 2594 358391 2650 358400
rect 2502 345400 2558 345409
rect 2502 345335 2558 345344
rect 2410 319288 2466 319297
rect 2410 319223 2466 319232
rect 2318 267200 2374 267209
rect 2318 267135 2374 267144
rect 3344 97617 3372 463626
rect 3330 97608 3386 97617
rect 3330 97543 3386 97552
rect 2226 58576 2282 58585
rect 2226 58511 2282 58520
rect 3436 45529 3464 699071
rect 3528 136785 3556 699314
rect 3620 149841 3648 699887
rect 3712 201929 3740 700402
rect 3792 699712 3844 699718
rect 3792 699654 3844 699660
rect 3804 619177 3832 699654
rect 3790 619168 3846 619177
rect 3790 619103 3846 619112
rect 3792 565888 3844 565894
rect 3792 565830 3844 565836
rect 3698 201920 3754 201929
rect 3698 201855 3754 201864
rect 3606 149832 3662 149841
rect 3606 149767 3662 149776
rect 3514 136776 3570 136785
rect 3514 136711 3570 136720
rect 3804 84697 3832 565830
rect 3896 241097 3924 700470
rect 4066 700088 4122 700097
rect 4066 700023 4122 700032
rect 3976 699508 4028 699514
rect 3976 699450 4028 699456
rect 3988 293185 4016 699450
rect 4080 306241 4108 700023
rect 4264 565894 4292 701791
rect 4344 701684 4396 701690
rect 4344 701626 4396 701632
rect 4356 661094 4384 701626
rect 4434 701584 4490 701593
rect 4434 701519 4490 701528
rect 4344 661088 4396 661094
rect 4344 661030 4396 661036
rect 4252 565888 4304 565894
rect 4252 565830 4304 565836
rect 4448 463690 4476 701519
rect 8128 701010 8156 703520
rect 21454 702536 21510 702545
rect 21454 702471 21510 702480
rect 8116 701004 8168 701010
rect 8116 700946 8168 700952
rect 21468 699938 21496 702471
rect 24320 700330 24348 703520
rect 35808 702500 35860 702506
rect 35808 702442 35860 702448
rect 24308 700324 24360 700330
rect 24308 700266 24360 700272
rect 35820 700210 35848 702442
rect 40512 700942 40540 703520
rect 60646 701992 60702 702001
rect 60646 701927 60702 701936
rect 46018 701720 46074 701729
rect 46018 701655 46074 701664
rect 40500 700936 40552 700942
rect 40500 700878 40552 700884
rect 35820 700182 35894 700210
rect 21160 699910 21496 699938
rect 35866 699924 35894 700182
rect 46032 699938 46060 701655
rect 55772 701072 55824 701078
rect 55772 701014 55824 701020
rect 55784 699938 55812 701014
rect 60660 699938 60688 701927
rect 70124 701888 70176 701894
rect 70124 701830 70176 701836
rect 45724 699910 46060 699938
rect 55476 699910 55812 699938
rect 60444 699910 60688 699938
rect 70136 699666 70164 701830
rect 72988 700874 73016 703520
rect 75460 702364 75512 702370
rect 75460 702306 75512 702312
rect 72976 700868 73028 700874
rect 72976 700810 73028 700816
rect 75472 699938 75500 702306
rect 85304 701208 85356 701214
rect 85304 701150 85356 701156
rect 85316 699938 85344 701150
rect 89180 700602 89208 703520
rect 104808 701412 104860 701418
rect 104808 701354 104860 701360
rect 100024 701344 100076 701350
rect 100024 701286 100076 701292
rect 90180 701276 90232 701282
rect 90180 701218 90232 701224
rect 89168 700596 89220 700602
rect 89168 700538 89220 700544
rect 90192 699938 90220 701218
rect 100036 699938 100064 701286
rect 104820 699938 104848 701354
rect 105464 700670 105492 703520
rect 129464 701616 129516 701622
rect 129464 701558 129516 701564
rect 119712 701480 119764 701486
rect 119712 701422 119764 701428
rect 105452 700664 105504 700670
rect 105452 700606 105504 700612
rect 119724 699938 119752 701422
rect 129476 699938 129504 701558
rect 134430 701176 134486 701185
rect 134430 701111 134486 701120
rect 134444 699938 134472 701111
rect 137848 700738 137876 703520
rect 154028 702432 154080 702438
rect 154028 702374 154080 702380
rect 148968 701752 149020 701758
rect 148968 701694 149020 701700
rect 137836 700732 137888 700738
rect 137836 700674 137888 700680
rect 148980 699938 149008 701694
rect 154040 699938 154068 702374
rect 154132 700126 154160 703520
rect 170324 703458 170352 703520
rect 170312 703452 170364 703458
rect 170312 703394 170364 703400
rect 198280 703180 198332 703186
rect 198280 703122 198332 703128
rect 183376 703044 183428 703050
rect 183376 702986 183428 702992
rect 158628 702908 158680 702914
rect 158628 702850 158680 702856
rect 158640 700210 158668 702850
rect 178592 702160 178644 702166
rect 178592 702102 178644 702108
rect 163872 702092 163924 702098
rect 163872 702034 163924 702040
rect 158640 700182 158714 700210
rect 154120 700120 154172 700126
rect 154120 700062 154172 700068
rect 75164 699910 75500 699938
rect 85008 699910 85344 699938
rect 89884 699910 90220 699938
rect 99728 699910 100064 699938
rect 104604 699910 104848 699938
rect 119416 699910 119752 699938
rect 129168 699910 129504 699938
rect 134136 699910 134472 699938
rect 148856 699910 149008 699938
rect 153732 699910 154068 699938
rect 158686 699924 158714 700182
rect 163884 699938 163912 702034
rect 178604 699938 178632 702102
rect 183388 699938 183416 702986
rect 188436 702024 188488 702030
rect 188436 701966 188488 701972
rect 188448 699938 188476 701966
rect 198292 699938 198320 703122
rect 202800 700806 202828 703520
rect 213000 703316 213052 703322
rect 213000 703258 213052 703264
rect 202788 700800 202840 700806
rect 202788 700742 202840 700748
rect 213012 699938 213040 703258
rect 163576 699910 163912 699938
rect 178296 699910 178632 699938
rect 183264 699910 183416 699938
rect 188140 699910 188476 699938
rect 197984 699910 198320 699938
rect 212704 699910 213040 699938
rect 218992 699922 219020 703520
rect 235184 703474 235212 703520
rect 235368 703474 235396 703530
rect 227628 703452 227680 703458
rect 235184 703446 235396 703474
rect 227628 703394 227680 703400
rect 227640 699938 227668 703394
rect 237104 702296 237156 702302
rect 237104 702238 237156 702244
rect 232688 700392 232740 700398
rect 232688 700334 232740 700340
rect 232700 699938 232728 700334
rect 218980 699916 219032 699922
rect 227424 699910 227668 699938
rect 232392 699910 232728 699938
rect 218980 699858 219032 699864
rect 217876 699848 217928 699854
rect 217580 699796 217876 699802
rect 217580 699790 217928 699796
rect 217580 699774 217916 699790
rect 237116 699666 237144 702238
rect 242452 699938 242480 703530
rect 251426 703520 251538 704960
rect 257252 703792 257304 703798
rect 257252 703734 257304 703740
rect 243360 702024 243412 702030
rect 243360 701966 243412 701972
rect 242144 699910 242480 699938
rect 70136 699638 70288 699666
rect 237116 699638 237268 699666
rect 243372 699446 243400 701966
rect 252284 700256 252336 700262
rect 252284 700198 252336 700204
rect 247086 700188 247138 700194
rect 247086 700130 247138 700136
rect 247098 699924 247126 700130
rect 252296 699938 252324 700198
rect 257264 699938 257292 703734
rect 267618 703520 267730 704960
rect 271788 703860 271840 703866
rect 271788 703802 271840 703808
rect 262128 702024 262180 702030
rect 262128 701966 262180 701972
rect 262140 700534 262168 701966
rect 266360 701956 266412 701962
rect 266360 701898 266412 701904
rect 262128 700528 262180 700534
rect 262128 700470 262180 700476
rect 266372 700466 266400 701898
rect 267660 700466 267688 703520
rect 271512 701072 271564 701078
rect 271512 701014 271564 701020
rect 266360 700460 266412 700466
rect 266360 700402 266412 700408
rect 267648 700460 267700 700466
rect 267648 700402 267700 700408
rect 267004 700052 267056 700058
rect 267004 699994 267056 700000
rect 262128 699984 262180 699990
rect 251988 699910 252324 699938
rect 256956 699910 257292 699938
rect 261832 699932 262128 699938
rect 267016 699938 267044 699994
rect 261832 699926 262180 699932
rect 261832 699910 262168 699926
rect 266708 699910 267044 699938
rect 271524 699582 271552 701014
rect 271800 699938 271828 703802
rect 276848 703724 276900 703730
rect 276848 703666 276900 703672
rect 276860 699938 276888 703666
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 300860 703656 300912 703662
rect 300860 703598 300912 703604
rect 283852 702434 283880 703520
rect 283852 702406 284156 702434
rect 282920 701072 282972 701078
rect 282920 701014 282972 701020
rect 281356 700528 281408 700534
rect 281356 700470 281408 700476
rect 271676 699910 271828 699938
rect 276552 699910 276888 699938
rect 281368 699802 281396 700470
rect 282932 700466 282960 701014
rect 284128 700466 284156 702406
rect 286690 701176 286746 701185
rect 286690 701111 286746 701120
rect 291474 701176 291530 701185
rect 291474 701111 291530 701120
rect 282920 700460 282972 700466
rect 282920 700402 282972 700408
rect 284116 700460 284168 700466
rect 284116 700402 284168 700408
rect 286704 699938 286732 701111
rect 291200 701072 291252 701078
rect 291200 701014 291252 701020
rect 291384 701072 291436 701078
rect 291384 701014 291436 701020
rect 291212 700074 291240 701014
rect 291396 700466 291424 701014
rect 291488 700466 291516 701111
rect 295892 701072 295944 701078
rect 295892 701014 295944 701020
rect 291384 700460 291436 700466
rect 291384 700402 291436 700408
rect 291476 700460 291528 700466
rect 291476 700402 291528 700408
rect 291212 700046 291286 700074
rect 286396 699910 286732 699938
rect 291258 699924 291286 700046
rect 295904 699938 295932 701014
rect 300136 700466 300164 703520
rect 300124 700460 300176 700466
rect 300124 700402 300176 700408
rect 300872 699938 300900 703598
rect 315488 703520 315540 703526
rect 316286 703520 316398 704960
rect 332324 703724 332376 703730
rect 332324 703666 332376 703672
rect 315488 703462 315540 703468
rect 332336 703474 332364 703666
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364708 703860 364760 703866
rect 364708 703802 364760 703808
rect 364720 703610 364748 703802
rect 364720 703582 364840 703610
rect 332520 703474 332548 703520
rect 311164 702432 311216 702438
rect 311164 702374 311216 702380
rect 305828 702296 305880 702302
rect 305828 702238 305880 702244
rect 305840 700806 305868 702238
rect 311072 702228 311124 702234
rect 311072 702170 311124 702176
rect 305736 700800 305788 700806
rect 305736 700742 305788 700748
rect 305828 700800 305880 700806
rect 305828 700742 305880 700748
rect 305748 699938 305776 700742
rect 295904 699910 296240 699938
rect 300872 699910 301116 699938
rect 305748 699910 306084 699938
rect 310624 699922 310960 699938
rect 310612 699916 310960 699922
rect 310664 699910 310960 699916
rect 310612 699858 310664 699864
rect 281368 699774 281520 699802
rect 311084 699650 311112 702170
rect 311176 700466 311204 702374
rect 311164 700460 311216 700466
rect 311164 700402 311216 700408
rect 315500 699938 315528 703462
rect 332336 703446 332548 703474
rect 339316 702160 339368 702166
rect 339316 702102 339368 702108
rect 331312 702092 331364 702098
rect 331312 702034 331364 702040
rect 335912 702092 335964 702098
rect 335912 702034 335964 702040
rect 329380 701888 329432 701894
rect 329380 701830 329432 701836
rect 320456 700732 320508 700738
rect 320456 700674 320508 700680
rect 320468 699938 320496 700674
rect 329392 700126 329420 701830
rect 331220 701072 331272 701078
rect 331220 701014 331272 701020
rect 331232 700874 331260 701014
rect 331220 700868 331272 700874
rect 331220 700810 331272 700816
rect 331324 700670 331352 702034
rect 335360 701072 335412 701078
rect 335360 701014 335412 701020
rect 330300 700664 330352 700670
rect 330300 700606 330352 700612
rect 331312 700664 331364 700670
rect 331312 700606 331364 700612
rect 325654 700120 325706 700126
rect 325654 700062 325706 700068
rect 329380 700120 329432 700126
rect 329380 700062 329432 700068
rect 315500 699910 315836 699938
rect 320468 699910 320804 699938
rect 325666 699924 325694 700062
rect 330312 699938 330340 700606
rect 330312 699910 330648 699938
rect 335372 699802 335400 701014
rect 335372 699774 335524 699802
rect 311072 699644 311124 699650
rect 311072 699586 311124 699592
rect 271512 699576 271564 699582
rect 271512 699518 271564 699524
rect 335924 699514 335952 702034
rect 339328 700738 339356 702102
rect 339408 701072 339460 701078
rect 339408 701014 339460 701020
rect 344928 701072 344980 701078
rect 344980 701020 345060 701026
rect 344928 701014 345060 701020
rect 339420 700942 339448 701014
rect 344940 700998 345060 701014
rect 339408 700936 339460 700942
rect 339408 700878 339460 700884
rect 339316 700732 339368 700738
rect 339316 700674 339368 700680
rect 340052 700596 340104 700602
rect 340052 700538 340104 700544
rect 340064 699938 340092 700538
rect 345032 699938 345060 700998
rect 348804 700534 348832 703520
rect 364812 703474 364840 703582
rect 364954 703520 365066 704960
rect 371608 703792 371660 703798
rect 371608 703734 371660 703740
rect 364996 703474 365024 703520
rect 364812 703446 365024 703474
rect 359740 703384 359792 703390
rect 359740 703326 359792 703332
rect 350540 701888 350592 701894
rect 350540 701830 350592 701836
rect 349896 701072 349948 701078
rect 349896 701014 349948 701020
rect 348792 700528 348844 700534
rect 348792 700470 348844 700476
rect 349908 699938 349936 701014
rect 340064 699910 340400 699938
rect 345032 699910 345368 699938
rect 349908 699910 350244 699938
rect 335912 699508 335964 699514
rect 335912 699450 335964 699456
rect 50896 699440 50948 699446
rect 6642 699408 6698 699417
rect 6440 699366 6642 699394
rect 11610 699408 11666 699417
rect 11316 699366 11610 699394
rect 6642 699343 6698 699352
rect 16394 699408 16450 699417
rect 16192 699366 16394 699394
rect 11610 699343 11666 699352
rect 26146 699408 26202 699417
rect 26036 699366 26146 699394
rect 16394 699343 16450 699352
rect 31206 699408 31262 699417
rect 30912 699366 31206 699394
rect 26146 699343 26202 699352
rect 41050 699408 41106 699417
rect 40756 699366 41050 699394
rect 31206 699343 31262 699352
rect 50600 699388 50896 699394
rect 65616 699440 65668 699446
rect 50600 699382 50948 699388
rect 65320 699388 65616 699394
rect 80152 699440 80204 699446
rect 65320 699382 65668 699388
rect 80040 699388 80152 699394
rect 95148 699440 95200 699446
rect 80040 699382 80204 699388
rect 94852 699388 95148 699394
rect 109868 699440 109920 699446
rect 94852 699382 95200 699388
rect 109572 699388 109868 699394
rect 114560 699440 114612 699446
rect 109572 699382 109920 699388
rect 114448 699388 114560 699394
rect 124588 699440 124640 699446
rect 114448 699382 114612 699388
rect 124292 699388 124588 699394
rect 139308 699440 139360 699446
rect 124292 699382 124640 699388
rect 139012 699388 139308 699394
rect 144276 699440 144328 699446
rect 139012 699382 139360 699388
rect 143980 699388 144276 699394
rect 168840 699440 168892 699446
rect 143980 699382 144328 699388
rect 168544 699388 168840 699394
rect 173716 699440 173768 699446
rect 168544 699382 168892 699388
rect 173420 699388 173716 699394
rect 208124 699440 208176 699446
rect 173420 699382 173768 699388
rect 50600 699366 50936 699382
rect 65320 699366 65656 699382
rect 80040 699366 80192 699382
rect 94852 699366 95188 699382
rect 109572 699366 109908 699382
rect 114448 699366 114600 699382
rect 124292 699366 124628 699382
rect 139012 699366 139348 699382
rect 143980 699366 144316 699382
rect 168544 699366 168880 699382
rect 173420 699366 173756 699382
rect 193108 699378 193260 699394
rect 202860 699378 203012 699394
rect 207828 699388 208124 699394
rect 243360 699440 243412 699446
rect 207828 699382 208176 699388
rect 193108 699372 193272 699378
rect 193108 699366 193220 699372
rect 41050 699343 41106 699352
rect 202860 699372 203024 699378
rect 202860 699366 202972 699372
rect 193220 699314 193272 699320
rect 207828 699366 208164 699382
rect 222548 699378 222884 699394
rect 243360 699382 243412 699388
rect 350552 699378 350580 701830
rect 354956 700324 355008 700330
rect 354956 700266 355008 700272
rect 354968 699938 354996 700266
rect 359752 699938 359780 703326
rect 364616 702228 364668 702234
rect 364616 702170 364668 702176
rect 364628 699938 364656 702170
rect 371620 700942 371648 703734
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 400864 703588 400916 703594
rect 400864 703530 400916 703536
rect 374460 703248 374512 703254
rect 374460 703190 374512 703196
rect 371608 700936 371660 700942
rect 371608 700878 371660 700884
rect 374472 699938 374500 703190
rect 389180 703112 389232 703118
rect 389180 703054 389232 703060
rect 379518 700632 379574 700641
rect 379518 700567 379574 700576
rect 379532 699938 379560 700567
rect 389192 699938 389220 703054
rect 397472 699990 397500 703520
rect 400876 701010 400904 703530
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 403900 702976 403952 702982
rect 403900 702918 403952 702924
rect 400864 701004 400916 701010
rect 400864 700946 400916 700952
rect 399022 700496 399078 700505
rect 399022 700431 399078 700440
rect 397460 699984 397512 699990
rect 354968 699910 355212 699938
rect 359752 699910 360088 699938
rect 364628 699910 364964 699938
rect 374472 699910 374808 699938
rect 379532 699910 379776 699938
rect 389192 699910 389528 699938
rect 397460 699926 397512 699932
rect 399036 699938 399064 700431
rect 403912 699938 403940 702918
rect 413664 700058 413692 703520
rect 423680 702840 423732 702846
rect 423680 702782 423732 702788
rect 414204 701820 414256 701826
rect 414204 701762 414256 701768
rect 413652 700052 413704 700058
rect 413652 699994 413704 700000
rect 399036 699910 399372 699938
rect 403912 699910 404248 699938
rect 369780 699786 369932 699802
rect 369768 699780 369932 699786
rect 369820 699774 369932 699780
rect 369768 699722 369820 699728
rect 384304 699712 384356 699718
rect 414216 699666 414244 701762
rect 423692 699938 423720 702782
rect 429856 700942 429884 703520
rect 443276 701684 443328 701690
rect 443276 701626 443328 701632
rect 444288 701684 444340 701690
rect 444288 701626 444340 701632
rect 429844 700936 429896 700942
rect 429844 700878 429896 700884
rect 428462 700360 428518 700369
rect 428462 700295 428518 700304
rect 428476 699938 428504 700295
rect 438628 700224 438684 700233
rect 438628 700159 438684 700168
rect 423692 699910 423936 699938
rect 428476 699910 428812 699938
rect 438642 699924 438670 700159
rect 443288 699938 443316 701626
rect 443288 699910 443624 699938
rect 384356 699660 384652 699666
rect 384304 699654 384652 699660
rect 384316 699638 384652 699654
rect 414092 699638 414244 699666
rect 433430 699544 433486 699553
rect 433486 699502 433780 699530
rect 433430 699479 433486 699488
rect 444300 699417 444328 701626
rect 458180 701548 458232 701554
rect 458180 701490 458232 701496
rect 458192 699938 458220 701490
rect 462332 700194 462360 703520
rect 477592 702772 477644 702778
rect 477592 702714 477644 702720
rect 467840 702092 467892 702098
rect 467840 702034 467892 702040
rect 462320 700188 462372 700194
rect 462320 700130 462372 700136
rect 467852 699938 467880 702034
rect 472714 700088 472770 700097
rect 472714 700023 472770 700032
rect 472728 699938 472756 700023
rect 477604 699938 477632 702714
rect 478524 700262 478552 703520
rect 482560 702024 482612 702030
rect 482560 701966 482612 701972
rect 478512 700256 478564 700262
rect 478512 700198 478564 700204
rect 482572 699938 482600 701966
rect 487436 701140 487488 701146
rect 487436 701082 487488 701088
rect 487448 699938 487476 701082
rect 494808 701010 494836 703520
rect 497464 703452 497516 703458
rect 497464 703394 497516 703400
rect 497280 702704 497332 702710
rect 497280 702646 497332 702652
rect 494796 701004 494848 701010
rect 494796 700946 494848 700952
rect 497292 699938 497320 702646
rect 497476 701010 497504 703394
rect 507124 702636 507176 702642
rect 507124 702578 507176 702584
rect 502340 701956 502392 701962
rect 502340 701898 502392 701904
rect 497464 701004 497516 701010
rect 497464 700946 497516 700952
rect 502352 699938 502380 701898
rect 507136 699938 507164 702578
rect 512000 701888 512052 701894
rect 512000 701830 512052 701836
rect 526718 701856 526774 701865
rect 512012 699938 512040 701830
rect 526718 701791 526774 701800
rect 516966 699952 517022 699961
rect 458192 699910 458344 699938
rect 467852 699910 468188 699938
rect 472728 699910 473064 699938
rect 477604 699910 477940 699938
rect 482572 699910 482908 699938
rect 487448 699910 487784 699938
rect 497292 699910 497628 699938
rect 502352 699910 502504 699938
rect 507136 699910 507472 699938
rect 512012 699910 512348 699938
rect 526732 699938 526760 701791
rect 527192 700398 527220 703520
rect 536840 702568 536892 702574
rect 536840 702510 536892 702516
rect 531686 701584 531742 701593
rect 531686 701519 531742 701528
rect 527180 700392 527232 700398
rect 527180 700334 527232 700340
rect 531700 699938 531728 701519
rect 536852 700210 536880 702510
rect 541532 701684 541584 701690
rect 541532 701626 541584 701632
rect 536852 700182 536926 700210
rect 517022 699910 517316 699938
rect 526732 699910 527068 699938
rect 531700 699910 532036 699938
rect 536898 699924 536926 700182
rect 541544 699938 541572 701626
rect 543476 700806 543504 703520
rect 546498 701448 546554 701457
rect 546498 701383 546554 701392
rect 543464 700800 543516 700806
rect 543464 700742 543516 700748
rect 546512 699938 546540 701383
rect 556250 701312 556306 701321
rect 556250 701247 556306 701256
rect 556264 699938 556292 701247
rect 559668 701010 559696 703520
rect 576400 703316 576452 703322
rect 576400 703258 576452 703264
rect 575112 703180 575164 703186
rect 575112 703122 575164 703128
rect 573732 703044 573784 703050
rect 573732 702986 573784 702992
rect 573456 702364 573508 702370
rect 573456 702306 573508 702312
rect 561126 702128 561182 702137
rect 561126 702063 561182 702072
rect 559656 701004 559708 701010
rect 559656 700946 559708 700952
rect 561140 699938 561168 702063
rect 565174 701992 565230 702001
rect 565174 701927 565230 701936
rect 541544 699910 541880 699938
rect 546512 699910 546756 699938
rect 556264 699910 556600 699938
rect 561140 699910 561476 699938
rect 516966 699887 517022 699896
rect 563520 699848 563572 699854
rect 551282 699816 551338 699825
rect 551338 699774 551632 699802
rect 563520 699790 563572 699796
rect 551282 699751 551338 699760
rect 408958 699408 409014 699417
rect 394160 699378 394496 699394
rect 222548 699372 222896 699378
rect 222548 699366 222844 699372
rect 202972 699314 203024 699320
rect 222844 699314 222896 699320
rect 350540 699372 350592 699378
rect 350540 699314 350592 699320
rect 394148 699372 394496 699378
rect 394200 699366 394496 699372
rect 418710 699408 418766 699417
rect 409014 699366 409216 699394
rect 408958 699343 409014 699352
rect 444286 699408 444342 699417
rect 418766 699366 419060 699394
rect 418710 699343 418766 699352
rect 444286 699343 444342 699352
rect 448150 699408 448206 699417
rect 453118 699408 453174 699417
rect 448206 699366 448500 699394
rect 448150 699343 448206 699352
rect 453174 699366 453376 699394
rect 462884 699378 463220 699394
rect 492600 699378 492752 699394
rect 521856 699378 522192 699394
rect 462872 699372 463220 699378
rect 453118 699343 453174 699352
rect 394148 699314 394200 699320
rect 462924 699366 463220 699372
rect 492588 699372 492752 699378
rect 462872 699314 462924 699320
rect 492640 699366 492752 699372
rect 521844 699372 522192 699378
rect 492588 699314 492640 699320
rect 521896 699366 522192 699372
rect 521844 699314 521896 699320
rect 563532 698290 563560 699790
rect 563704 699304 563756 699310
rect 563704 699246 563756 699252
rect 563520 698284 563572 698290
rect 563520 698226 563572 698232
rect 563716 684486 563744 699246
rect 565082 698320 565138 698329
rect 565082 698255 565138 698264
rect 563704 684480 563756 684486
rect 563704 684422 563756 684428
rect 4436 463684 4488 463690
rect 4436 463626 4488 463632
rect 4066 306232 4122 306241
rect 4066 306167 4122 306176
rect 3974 293176 4030 293185
rect 3974 293111 4030 293120
rect 3882 241088 3938 241097
rect 3882 241023 3938 241032
rect 3790 84688 3846 84697
rect 3790 84623 3846 84632
rect 3422 45520 3478 45529
rect 3422 45455 3478 45464
rect 2134 32464 2190 32473
rect 2134 32399 2190 32408
rect 565096 6866 565124 698255
rect 565188 139398 565216 701927
rect 571982 701720 572038 701729
rect 571982 701655 572038 701664
rect 569316 701208 569368 701214
rect 569316 701150 569368 701156
rect 567844 699236 567896 699242
rect 567844 699178 567896 699184
rect 566646 699000 566702 699009
rect 566646 698935 566702 698944
rect 566832 698964 566884 698970
rect 565266 698728 565322 698737
rect 565266 698663 565322 698672
rect 565176 139392 565228 139398
rect 565176 139334 565228 139340
rect 565280 73166 565308 698663
rect 566462 698592 566518 698601
rect 566462 698527 566518 698536
rect 565360 698488 565412 698494
rect 565360 698430 565412 698436
rect 565372 245614 565400 698430
rect 565360 245608 565412 245614
rect 565360 245550 565412 245556
rect 565268 73160 565320 73166
rect 565268 73102 565320 73108
rect 566476 20670 566504 698527
rect 566556 698352 566608 698358
rect 566556 698294 566608 698300
rect 566568 167006 566596 698294
rect 566556 167000 566608 167006
rect 566556 166942 566608 166948
rect 566660 113150 566688 698935
rect 566832 698906 566884 698912
rect 566740 698420 566792 698426
rect 566740 698362 566792 698368
rect 566752 206990 566780 698362
rect 566844 511970 566872 698906
rect 567856 632058 567884 699178
rect 569222 698456 569278 698465
rect 569222 698391 569278 698400
rect 567844 632052 567896 632058
rect 567844 631994 567896 632000
rect 566832 511964 566884 511970
rect 566832 511906 566884 511912
rect 566740 206984 566792 206990
rect 566740 206926 566792 206932
rect 566648 113144 566700 113150
rect 566648 113086 566700 113092
rect 569236 33114 569264 698391
rect 569328 233238 569356 701150
rect 569406 698864 569462 698873
rect 569406 698799 569462 698808
rect 570696 698828 570748 698834
rect 569316 233232 569368 233238
rect 569316 233174 569368 233180
rect 569420 60722 569448 698799
rect 570696 698770 570748 698776
rect 570604 698624 570656 698630
rect 570604 698566 570656 698572
rect 569500 698556 569552 698562
rect 569500 698498 569552 698504
rect 569512 299470 569540 698498
rect 570616 325650 570644 698566
rect 570708 405686 570736 698770
rect 570696 405680 570748 405686
rect 570696 405622 570748 405628
rect 570604 325644 570656 325650
rect 570604 325586 570656 325592
rect 569500 299464 569552 299470
rect 569500 299406 569552 299412
rect 571996 100706 572024 701655
rect 572168 699100 572220 699106
rect 572168 699042 572220 699048
rect 572076 698692 572128 698698
rect 572076 698634 572128 698640
rect 572088 353258 572116 698634
rect 572180 578202 572208 699042
rect 573364 697604 573416 697610
rect 573364 697546 573416 697552
rect 572168 578196 572220 578202
rect 572168 578138 572220 578144
rect 572076 353252 572128 353258
rect 572076 353194 572128 353200
rect 573376 126954 573404 697546
rect 573468 179382 573496 702306
rect 573548 701276 573600 701282
rect 573548 701218 573600 701224
rect 573560 219434 573588 701218
rect 573640 698896 573692 698902
rect 573640 698838 573692 698844
rect 573652 538218 573680 698838
rect 573744 564398 573772 702986
rect 575020 702908 575072 702914
rect 575020 702850 575072 702856
rect 574744 702500 574796 702506
rect 574744 702442 574796 702448
rect 573732 564392 573784 564398
rect 573732 564334 573784 564340
rect 573640 538212 573692 538218
rect 573640 538154 573692 538160
rect 573548 219428 573600 219434
rect 573548 219370 573600 219376
rect 573456 179376 573508 179382
rect 573456 179318 573508 179324
rect 573364 126948 573416 126954
rect 573364 126890 573416 126896
rect 571984 100700 572036 100706
rect 571984 100642 572036 100648
rect 574756 86970 574784 702442
rect 574928 701616 574980 701622
rect 574928 701558 574980 701564
rect 574836 701412 574888 701418
rect 574836 701354 574888 701360
rect 574848 259418 574876 701354
rect 574940 379506 574968 701558
rect 575032 485790 575060 702850
rect 575124 618254 575152 703122
rect 576122 702536 576178 702545
rect 576122 702471 576178 702480
rect 575112 618248 575164 618254
rect 575112 618190 575164 618196
rect 575020 485784 575072 485790
rect 575020 485726 575072 485732
rect 574928 379500 574980 379506
rect 574928 379442 574980 379448
rect 574836 259412 574888 259418
rect 574836 259354 574888 259360
rect 574744 86964 574796 86970
rect 574744 86906 574796 86912
rect 569408 60716 569460 60722
rect 569408 60658 569460 60664
rect 576136 46918 576164 702471
rect 576308 701480 576360 701486
rect 576308 701422 576360 701428
rect 576216 701344 576268 701350
rect 576216 701286 576268 701292
rect 576228 273222 576256 701286
rect 576320 313274 576348 701422
rect 576412 672042 576440 703258
rect 577504 701752 577556 701758
rect 577504 701694 577556 701700
rect 576400 672036 576452 672042
rect 576400 671978 576452 671984
rect 577516 419490 577544 701694
rect 580724 700732 580776 700738
rect 580724 700674 580776 700680
rect 580632 700664 580684 700670
rect 580632 700606 580684 700612
rect 580540 700460 580592 700466
rect 580540 700402 580592 700408
rect 580356 700120 580408 700126
rect 580356 700062 580408 700068
rect 580264 699576 580316 699582
rect 580264 699518 580316 699524
rect 578976 699168 579028 699174
rect 578976 699110 579028 699116
rect 578884 698760 578936 698766
rect 578884 698702 578936 698708
rect 578896 431633 578924 698702
rect 578988 644065 579016 699110
rect 580172 698284 580224 698290
rect 580172 698226 580224 698232
rect 580184 697241 580212 698226
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580172 684480 580224 684486
rect 580172 684422 580224 684428
rect 580184 683913 580212 684422
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580172 672036 580224 672042
rect 580172 671978 580224 671984
rect 580184 670721 580212 671978
rect 580170 670712 580226 670721
rect 580170 670647 580226 670656
rect 578974 644056 579030 644065
rect 578974 643991 579030 644000
rect 580172 632052 580224 632058
rect 580172 631994 580224 632000
rect 580184 630873 580212 631994
rect 580170 630864 580226 630873
rect 580170 630799 580226 630808
rect 580172 618248 580224 618254
rect 580172 618190 580224 618196
rect 580184 617545 580212 618190
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 579804 578196 579856 578202
rect 579804 578138 579856 578144
rect 579816 577697 579844 578138
rect 579802 577688 579858 577697
rect 579802 577623 579858 577632
rect 580172 564392 580224 564398
rect 580170 564360 580172 564369
rect 580224 564360 580226 564369
rect 580170 564295 580226 564304
rect 580172 538212 580224 538218
rect 580172 538154 580224 538160
rect 580184 537849 580212 538154
rect 580170 537840 580226 537849
rect 580170 537775 580226 537784
rect 580172 511964 580224 511970
rect 580172 511906 580224 511912
rect 580184 511329 580212 511906
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 579620 485784 579672 485790
rect 579620 485726 579672 485732
rect 579632 484673 579660 485726
rect 579618 484664 579674 484673
rect 579618 484599 579674 484608
rect 578882 431624 578938 431633
rect 578882 431559 578938 431568
rect 577504 419484 577556 419490
rect 577504 419426 577556 419432
rect 579620 419484 579672 419490
rect 579620 419426 579672 419432
rect 579632 418305 579660 419426
rect 579618 418296 579674 418305
rect 579618 418231 579674 418240
rect 579804 405680 579856 405686
rect 579804 405622 579856 405628
rect 579816 404977 579844 405622
rect 579802 404968 579858 404977
rect 579802 404903 579858 404912
rect 579804 379500 579856 379506
rect 579804 379442 579856 379448
rect 579816 378457 579844 379442
rect 579802 378448 579858 378457
rect 579802 378383 579858 378392
rect 580172 353252 580224 353258
rect 580172 353194 580224 353200
rect 580184 351937 580212 353194
rect 580170 351928 580226 351937
rect 580170 351863 580226 351872
rect 580172 325644 580224 325650
rect 580172 325586 580224 325592
rect 580184 325281 580212 325586
rect 580170 325272 580226 325281
rect 580170 325207 580226 325216
rect 576308 313268 576360 313274
rect 576308 313210 576360 313216
rect 580172 313268 580224 313274
rect 580172 313210 580224 313216
rect 580184 312089 580212 313210
rect 580170 312080 580226 312089
rect 580170 312015 580226 312024
rect 580172 299464 580224 299470
rect 580172 299406 580224 299412
rect 580184 298761 580212 299406
rect 580170 298752 580226 298761
rect 580170 298687 580226 298696
rect 576216 273216 576268 273222
rect 576216 273158 576268 273164
rect 580172 273216 580224 273222
rect 580172 273158 580224 273164
rect 580184 272241 580212 273158
rect 580170 272232 580226 272241
rect 580170 272167 580226 272176
rect 579620 259412 579672 259418
rect 579620 259354 579672 259360
rect 579632 258913 579660 259354
rect 579618 258904 579674 258913
rect 579618 258839 579674 258848
rect 580172 245608 580224 245614
rect 580170 245576 580172 245585
rect 580224 245576 580226 245585
rect 580170 245511 580226 245520
rect 580172 233232 580224 233238
rect 580172 233174 580224 233180
rect 580184 232393 580212 233174
rect 580170 232384 580226 232393
rect 580170 232319 580226 232328
rect 580172 219428 580224 219434
rect 580172 219370 580224 219376
rect 580184 219065 580212 219370
rect 580170 219056 580226 219065
rect 580170 218991 580226 219000
rect 579896 206984 579948 206990
rect 579896 206926 579948 206932
rect 579908 205737 579936 206926
rect 579894 205728 579950 205737
rect 579894 205663 579950 205672
rect 579988 179376 580040 179382
rect 579988 179318 580040 179324
rect 580000 179217 580028 179318
rect 579986 179208 580042 179217
rect 579986 179143 580042 179152
rect 580172 167000 580224 167006
rect 580172 166942 580224 166948
rect 580184 165889 580212 166942
rect 580170 165880 580226 165889
rect 580170 165815 580226 165824
rect 580276 152697 580304 699518
rect 580368 192545 580396 700062
rect 580446 698048 580502 698057
rect 580446 697983 580502 697992
rect 580460 365129 580488 697983
rect 580552 458153 580580 700402
rect 580644 471481 580672 700606
rect 580736 524521 580764 700674
rect 580816 699440 580868 699446
rect 580816 699382 580868 699388
rect 580828 591025 580856 699382
rect 580814 591016 580870 591025
rect 580814 590951 580870 590960
rect 580722 524512 580778 524521
rect 580722 524447 580778 524456
rect 580630 471472 580686 471481
rect 580630 471407 580686 471416
rect 580538 458144 580594 458153
rect 580538 458079 580594 458088
rect 580446 365120 580502 365129
rect 580446 365055 580502 365064
rect 580354 192536 580410 192545
rect 580354 192471 580410 192480
rect 580262 152688 580318 152697
rect 580262 152623 580318 152632
rect 580172 139392 580224 139398
rect 580170 139360 580172 139369
rect 580224 139360 580226 139369
rect 580170 139295 580226 139304
rect 580172 126948 580224 126954
rect 580172 126890 580224 126896
rect 580184 126041 580212 126890
rect 580170 126032 580226 126041
rect 580170 125967 580226 125976
rect 579804 113144 579856 113150
rect 579804 113086 579856 113092
rect 579816 112849 579844 113086
rect 579802 112840 579858 112849
rect 579802 112775 579858 112784
rect 580172 100700 580224 100706
rect 580172 100642 580224 100648
rect 580184 99521 580212 100642
rect 580170 99512 580226 99521
rect 580170 99447 580226 99456
rect 580172 86964 580224 86970
rect 580172 86906 580224 86912
rect 580184 86193 580212 86906
rect 580170 86184 580226 86193
rect 580170 86119 580226 86128
rect 580172 73160 580224 73166
rect 580172 73102 580224 73108
rect 580184 73001 580212 73102
rect 580170 72992 580226 73001
rect 580170 72927 580226 72936
rect 580172 60716 580224 60722
rect 580172 60658 580224 60664
rect 580184 59673 580212 60658
rect 580170 59664 580226 59673
rect 580170 59599 580226 59608
rect 576124 46912 576176 46918
rect 576124 46854 576176 46860
rect 580172 46912 580224 46918
rect 580172 46854 580224 46860
rect 580184 46345 580212 46854
rect 580170 46336 580226 46345
rect 580170 46271 580226 46280
rect 580170 33144 580226 33153
rect 569224 33108 569276 33114
rect 580170 33079 580172 33088
rect 569224 33050 569276 33056
rect 580224 33079 580226 33088
rect 580172 33050 580224 33056
rect 566464 20664 566516 20670
rect 566464 20606 566516 20612
rect 579988 20664 580040 20670
rect 579988 20606 580040 20612
rect 580000 19825 580028 20606
rect 579986 19816 580042 19825
rect 579986 19751 580042 19760
rect 565084 6860 565136 6866
rect 565084 6802 565136 6808
rect 580172 6860 580224 6866
rect 580172 6802 580224 6808
rect 580184 6633 580212 6802
rect 580170 6624 580226 6633
rect 580170 6559 580226 6568
rect 2042 6488 2098 6497
rect 2042 6423 2098 6432
rect 563704 3052 563756 3058
rect 563704 2994 563756 3000
rect 583392 3052 583444 3058
rect 583392 2994 583444 3000
rect 563520 2916 563572 2922
rect 563520 2858 563572 2864
rect 563532 1086 563560 2858
rect 563520 1080 563572 1086
rect 563520 1022 563572 1028
rect 563716 762 563744 2994
rect 572720 2916 572772 2922
rect 572720 2858 572772 2864
rect 569868 2848 569920 2854
rect 569868 2790 569920 2796
rect 569880 1018 569908 2790
rect 569868 1012 569920 1018
rect 569868 954 569920 960
rect 569132 944 569184 950
rect 569132 886 569184 892
rect 566832 876 566884 882
rect 566832 818 566884 824
rect 1676 672 1728 678
rect 5356 672 5408 678
rect 1676 614 1728 620
rect 4066 640 4122 649
rect 572 604 624 610
rect 572 546 624 552
rect 584 480 612 546
rect 1688 480 1716 614
rect 2884 564 3096 592
rect 4356 610 4600 626
rect 6460 672 6512 678
rect 5408 620 5704 626
rect 5356 614 5704 620
rect 10048 672 10100 678
rect 7838 640 7894 649
rect 6460 614 6512 620
rect 4066 575 4122 584
rect 4344 604 4600 610
rect 2884 480 2912 564
rect 3068 490 3096 564
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 3068 474 3280 490
rect 4080 480 4108 575
rect 4396 598 4600 604
rect 5264 604 5316 610
rect 4344 546 4396 552
rect 5368 598 5704 614
rect 5264 546 5316 552
rect 5276 480 5304 546
rect 6472 480 6500 614
rect 7484 598 7696 626
rect 7484 542 7512 598
rect 7472 536 7524 542
rect 3068 468 3292 474
rect 3068 462 3240 468
rect 3240 410 3292 416
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 6656 474 6808 490
rect 7472 478 7524 484
rect 7668 480 7696 598
rect 9954 640 10010 649
rect 7894 598 8004 626
rect 8588 598 8800 626
rect 8864 610 9108 626
rect 7838 575 7894 584
rect 8588 542 8616 598
rect 8576 536 8628 542
rect 6644 468 6808 474
rect 6696 462 6808 468
rect 6644 410 6696 416
rect 7626 -960 7738 480
rect 8576 478 8628 484
rect 8772 480 8800 598
rect 8852 604 9108 610
rect 8904 598 9108 604
rect 11520 672 11572 678
rect 10100 620 10212 626
rect 10048 614 10212 620
rect 10060 598 10212 614
rect 11408 620 11520 626
rect 19432 672 19484 678
rect 11408 614 11572 620
rect 13266 640 13322 649
rect 11152 604 11204 610
rect 9954 575 10010 584
rect 8852 546 8904 552
rect 9968 480 9996 575
rect 11408 598 11560 614
rect 12348 604 12400 610
rect 11152 546 11204 552
rect 13322 598 13616 626
rect 14476 598 14812 626
rect 15580 610 15916 626
rect 15568 604 15916 610
rect 13266 575 13322 584
rect 12348 546 12400 552
rect 11164 480 11192 546
rect 12360 480 12388 546
rect 12624 536 12676 542
rect 12512 484 12624 490
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 12512 478 12676 484
rect 13268 536 13320 542
rect 13268 478 13320 484
rect 12512 462 12664 478
rect 13280 218 13308 478
rect 13514 218 13626 480
rect 14476 474 14504 598
rect 15620 598 15916 604
rect 16684 598 17020 626
rect 17880 598 18216 626
rect 22376 672 22428 678
rect 19432 614 19484 620
rect 20626 640 20682 649
rect 15568 546 15620 552
rect 16684 542 16712 598
rect 16672 536 16724 542
rect 14464 468 14516 474
rect 14464 410 14516 416
rect 14556 400 14608 406
rect 14710 354 14822 480
rect 14608 348 14822 354
rect 14556 342 14822 348
rect 14568 326 14822 342
rect 13280 190 13626 218
rect 13514 -960 13626 190
rect 14710 -960 14822 326
rect 15906 82 16018 480
rect 16672 478 16724 484
rect 17408 536 17460 542
rect 17010 354 17122 480
rect 17408 478 17460 484
rect 17420 354 17448 478
rect 17880 406 17908 598
rect 18510 504 18566 513
rect 17010 326 17448 354
rect 17868 400 17920 406
rect 17868 342 17920 348
rect 16304 128 16356 134
rect 15906 76 16304 82
rect 15906 70 16356 76
rect 15906 54 16344 70
rect 15906 -960 16018 54
rect 17010 -960 17122 326
rect 18206 218 18318 480
rect 19444 480 19472 614
rect 24860 672 24912 678
rect 23478 640 23534 649
rect 22428 620 22724 626
rect 22376 614 22724 620
rect 20626 575 20682 584
rect 21824 604 21876 610
rect 20076 536 20128 542
rect 20128 484 20424 490
rect 18510 439 18566 448
rect 18524 218 18552 439
rect 18206 190 18552 218
rect 18206 -960 18318 190
rect 18972 128 19024 134
rect 19024 76 19320 82
rect 18972 70 19320 76
rect 18984 54 19320 70
rect 19402 -960 19514 480
rect 20076 478 20424 484
rect 20640 480 20668 575
rect 22388 598 22724 614
rect 23020 604 23072 610
rect 21824 546 21876 552
rect 23534 598 23828 626
rect 25320 672 25372 678
rect 24912 620 25024 626
rect 24860 614 25024 620
rect 28080 672 28132 678
rect 26514 640 26570 649
rect 25320 614 25372 620
rect 24872 598 25024 614
rect 23478 575 23534 584
rect 23020 546 23072 552
rect 24228 564 24440 592
rect 21270 504 21326 513
rect 20088 462 20424 478
rect 20598 -960 20710 480
rect 21326 462 21620 490
rect 21836 480 21864 546
rect 23032 480 23060 546
rect 24228 480 24256 564
rect 21270 439 21326 448
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 24412 474 24440 564
rect 25332 480 25360 614
rect 25792 610 26128 626
rect 25780 604 26128 610
rect 25832 598 26128 604
rect 28724 672 28776 678
rect 28722 640 28724 649
rect 29184 672 29236 678
rect 28776 640 28778 649
rect 28132 620 28428 626
rect 28080 614 28428 620
rect 28092 598 28428 614
rect 26514 575 26570 584
rect 25780 546 25832 552
rect 26528 480 26556 575
rect 27724 564 27936 592
rect 31300 672 31352 678
rect 30286 640 30342 649
rect 29236 620 29532 626
rect 29184 614 29532 620
rect 28722 575 28778 584
rect 28816 604 28868 610
rect 24400 468 24452 474
rect 24400 410 24452 416
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 26896 474 27232 490
rect 27724 480 27752 564
rect 27908 513 27936 564
rect 29196 598 29532 614
rect 30104 604 30156 610
rect 28868 564 28948 592
rect 28816 546 28868 552
rect 27894 504 27950 513
rect 26884 468 27232 474
rect 26936 462 27232 468
rect 26884 410 26936 416
rect 27682 -960 27794 480
rect 28920 480 28948 564
rect 30342 598 30636 626
rect 33784 672 33836 678
rect 31300 614 31352 620
rect 32402 640 32458 649
rect 30286 575 30342 584
rect 30104 546 30156 552
rect 30116 480 30144 546
rect 31312 480 31340 614
rect 33230 640 33286 649
rect 32600 610 32936 626
rect 32402 575 32458 584
rect 32588 604 32936 610
rect 31668 536 31720 542
rect 31720 484 31832 490
rect 27894 439 27950 448
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 31668 478 31832 484
rect 32416 480 32444 575
rect 32640 598 32936 604
rect 34796 672 34848 678
rect 33836 620 34132 626
rect 33784 614 34132 620
rect 37280 672 37332 678
rect 34796 614 34848 620
rect 35990 640 36046 649
rect 33230 575 33286 584
rect 33600 604 33652 610
rect 32588 546 32640 552
rect 33244 542 33272 575
rect 33796 598 34132 614
rect 33600 546 33652 552
rect 33232 536 33284 542
rect 31680 462 31832 478
rect 32374 -960 32486 480
rect 33232 478 33284 484
rect 33612 480 33640 546
rect 34808 480 34836 614
rect 36096 610 36340 626
rect 38384 672 38436 678
rect 37332 620 37536 626
rect 37280 614 37536 620
rect 40684 672 40736 678
rect 38384 614 38436 620
rect 38474 640 38530 649
rect 35990 575 36046 584
rect 36084 604 36340 610
rect 34980 536 35032 542
rect 35032 484 35236 490
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 34980 478 35236 484
rect 36004 480 36032 575
rect 36136 598 36340 604
rect 37188 604 37240 610
rect 36084 546 36136 552
rect 37292 598 37536 614
rect 37188 546 37240 552
rect 37200 480 37228 546
rect 38396 480 38424 614
rect 38530 598 38640 626
rect 39316 598 39620 626
rect 42800 672 42852 678
rect 40684 614 40736 620
rect 38474 575 38530 584
rect 34992 462 35236 478
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39316 406 39344 598
rect 39592 480 39620 598
rect 39304 400 39356 406
rect 39304 342 39356 348
rect 39550 -960 39662 480
rect 39744 474 39896 490
rect 40696 480 40724 614
rect 40788 610 40940 626
rect 46664 672 46716 678
rect 42852 620 43148 626
rect 42800 614 43148 620
rect 40776 604 40940 610
rect 40828 598 40940 604
rect 41880 604 41932 610
rect 40776 546 40828 552
rect 42812 598 43148 614
rect 44008 610 44344 626
rect 43996 604 44344 610
rect 41880 546 41932 552
rect 44048 598 44344 604
rect 45112 598 45448 626
rect 46664 614 46716 620
rect 48504 672 48556 678
rect 48964 672 49016 678
rect 48556 620 48852 626
rect 48504 614 48852 620
rect 50804 672 50856 678
rect 48964 614 49016 620
rect 43996 546 44048 552
rect 41892 480 41920 546
rect 39744 468 39908 474
rect 39744 462 39856 468
rect 39856 410 39908 416
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 42156 400 42208 406
rect 42044 348 42156 354
rect 42044 342 42208 348
rect 42892 400 42944 406
rect 43046 354 43158 480
rect 42944 348 43158 354
rect 42892 342 43158 348
rect 42044 326 42196 342
rect 42904 326 43158 342
rect 43046 -960 43158 326
rect 44242 82 44354 480
rect 45112 406 45140 598
rect 46676 480 46704 614
rect 47860 604 47912 610
rect 48516 598 48852 614
rect 47860 546 47912 552
rect 47872 480 47900 546
rect 48976 480 49004 614
rect 49620 610 49956 626
rect 53748 672 53800 678
rect 52550 640 52606 649
rect 50856 620 51152 626
rect 50804 614 51152 620
rect 49608 604 49956 610
rect 49660 598 49956 604
rect 50160 604 50212 610
rect 49608 546 49660 552
rect 50816 598 51152 614
rect 51356 604 51408 610
rect 50160 546 50212 552
rect 53024 610 53360 626
rect 53748 614 53800 620
rect 55404 672 55456 678
rect 64328 672 64380 678
rect 56046 640 56102 649
rect 55456 620 55660 626
rect 55404 614 55660 620
rect 52550 575 52606 584
rect 53012 604 53360 610
rect 51356 546 51408 552
rect 50172 480 50200 546
rect 51368 480 51396 546
rect 51908 536 51960 542
rect 51960 484 52256 490
rect 45100 400 45152 406
rect 45100 342 45152 348
rect 44100 66 44354 82
rect 44088 60 44354 66
rect 44140 54 44354 60
rect 44088 2 44140 8
rect 44242 -960 44354 54
rect 45438 82 45550 480
rect 45744 128 45796 134
rect 45438 76 45744 82
rect 45438 70 45796 76
rect 45438 54 45784 70
rect 46216 66 46552 82
rect 46204 60 46552 66
rect 45438 -960 45550 54
rect 46256 54 46552 60
rect 46204 2 46256 8
rect 46634 -960 46746 480
rect 47400 128 47452 134
rect 47452 76 47748 82
rect 47400 70 47748 76
rect 47412 54 47748 70
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 51908 478 52256 484
rect 52564 480 52592 575
rect 53064 598 53360 604
rect 53012 546 53064 552
rect 53760 480 53788 614
rect 54944 604 54996 610
rect 55416 598 55660 614
rect 57610 640 57666 649
rect 56428 610 56764 626
rect 56046 575 56102 584
rect 56416 604 56764 610
rect 54944 546 54996 552
rect 54206 504 54262 513
rect 51920 462 52256 478
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54262 462 54556 490
rect 54956 480 54984 546
rect 56060 480 56088 575
rect 56468 598 56764 604
rect 56416 546 56468 552
rect 57256 564 57468 592
rect 58438 640 58494 649
rect 57666 598 57960 626
rect 57610 575 57666 584
rect 59818 640 59874 649
rect 58438 575 58494 584
rect 57256 480 57284 564
rect 57440 513 57468 564
rect 57426 504 57482 513
rect 54206 439 54262 448
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58452 480 58480 575
rect 59464 564 59676 592
rect 62026 640 62082 649
rect 59874 598 60168 626
rect 60832 604 60884 610
rect 59818 575 59874 584
rect 59464 513 59492 564
rect 58806 504 58862 513
rect 57426 439 57482 448
rect 58410 -960 58522 480
rect 59450 504 59506 513
rect 58862 462 59064 490
rect 58806 439 58862 448
rect 59648 480 59676 564
rect 63498 640 63554 649
rect 62132 610 62468 626
rect 62026 575 62082 584
rect 62120 604 62468 610
rect 60832 546 60884 552
rect 60844 480 60872 546
rect 61106 504 61162 513
rect 59450 439 59506 448
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61162 462 61364 490
rect 62040 480 62068 575
rect 62172 598 62468 604
rect 62120 546 62172 552
rect 63236 564 63448 592
rect 63554 598 63664 626
rect 64328 614 64380 620
rect 65616 672 65668 678
rect 66720 672 66772 678
rect 65668 620 65872 626
rect 65616 614 65872 620
rect 68008 672 68060 678
rect 66720 614 66772 620
rect 63498 575 63554 584
rect 63236 480 63264 564
rect 63420 490 63448 564
rect 63500 536 63552 542
rect 63420 484 63500 490
rect 61106 439 61162 448
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 63420 478 63552 484
rect 64340 480 64368 614
rect 65524 604 65576 610
rect 65628 598 65872 614
rect 65524 546 65576 552
rect 64512 536 64564 542
rect 64564 484 64768 490
rect 63420 462 63540 478
rect 64298 -960 64410 480
rect 64512 478 64768 484
rect 65536 480 65564 546
rect 66732 480 66760 614
rect 66824 610 67068 626
rect 66812 604 67068 610
rect 66864 598 67068 604
rect 67744 598 67956 626
rect 69112 672 69164 678
rect 68060 620 68172 626
rect 68008 614 68172 620
rect 70584 672 70636 678
rect 69112 614 69164 620
rect 70472 620 70584 626
rect 133236 672 133288 678
rect 70472 614 70636 620
rect 68020 598 68172 614
rect 66812 546 66864 552
rect 67744 542 67772 598
rect 67732 536 67784 542
rect 64524 462 64768 478
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67732 478 67784 484
rect 67928 480 67956 598
rect 69124 480 69152 614
rect 70308 604 70360 610
rect 70472 598 70624 614
rect 71240 610 71576 626
rect 71228 604 71576 610
rect 70308 546 70360 552
rect 71280 598 71576 604
rect 72344 598 72680 626
rect 73540 598 73876 626
rect 74644 598 74980 626
rect 76944 610 77280 626
rect 78048 610 78384 626
rect 79152 610 79488 626
rect 80348 610 80684 626
rect 81452 610 81788 626
rect 82740 610 82892 626
rect 76196 604 76248 610
rect 71228 546 71280 552
rect 69388 536 69440 542
rect 69276 484 69388 490
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 69276 478 69440 484
rect 70320 480 70348 546
rect 69276 462 69428 478
rect 70278 -960 70390 480
rect 71320 400 71372 406
rect 71474 354 71586 480
rect 72344 406 72372 598
rect 71372 348 71586 354
rect 71320 342 71586 348
rect 72332 400 72384 406
rect 72332 342 72384 348
rect 72424 400 72476 406
rect 72578 354 72690 480
rect 73540 406 73568 598
rect 72476 348 72690 354
rect 72424 342 72690 348
rect 73528 400 73580 406
rect 73528 342 73580 348
rect 73620 400 73672 406
rect 73774 354 73886 480
rect 74644 406 74672 598
rect 76196 546 76248 552
rect 76932 604 77280 610
rect 76984 598 77280 604
rect 77392 604 77444 610
rect 76932 546 76984 552
rect 77392 546 77444 552
rect 78036 604 78384 610
rect 78088 598 78384 604
rect 78588 604 78640 610
rect 78036 546 78088 552
rect 78588 546 78640 552
rect 79140 604 79488 610
rect 79192 598 79488 604
rect 79692 604 79744 610
rect 79140 546 79192 552
rect 79692 546 79744 552
rect 80336 604 80684 610
rect 80388 598 80684 604
rect 80888 604 80940 610
rect 80336 546 80388 552
rect 80888 546 80940 552
rect 81440 604 81788 610
rect 81492 598 81788 604
rect 82084 604 82136 610
rect 81440 546 81492 552
rect 82084 546 82136 552
rect 82728 604 82892 610
rect 82780 598 82892 604
rect 83292 598 83504 626
rect 82728 546 82780 552
rect 76208 480 76236 546
rect 77404 480 77432 546
rect 78600 480 78628 546
rect 79704 480 79732 546
rect 80900 480 80928 546
rect 82096 480 82124 546
rect 83292 480 83320 598
rect 83476 490 83504 598
rect 84488 598 85192 626
rect 85684 598 85896 626
rect 73672 348 73886 354
rect 73620 342 73886 348
rect 74632 400 74684 406
rect 74632 342 74684 348
rect 71332 326 71586 342
rect 72436 326 72690 342
rect 73632 326 73886 342
rect 71474 -960 71586 326
rect 72578 -960 72690 326
rect 73774 -960 73886 326
rect 74970 82 75082 480
rect 74970 54 76084 82
rect 74970 -960 75082 54
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 83476 462 84088 490
rect 84488 480 84516 598
rect 85684 480 85712 598
rect 85868 490 85896 598
rect 86880 598 87492 626
rect 87984 598 88596 626
rect 89180 598 89392 626
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 85868 462 86296 490
rect 86880 480 86908 598
rect 87984 480 88012 598
rect 89180 480 89208 598
rect 89364 490 89392 598
rect 90376 598 90896 626
rect 91572 598 92000 626
rect 92768 598 93196 626
rect 93964 598 94300 626
rect 95160 598 95404 626
rect 96264 598 96600 626
rect 97460 598 97704 626
rect 98656 598 98808 626
rect 99852 598 100004 626
rect 105616 598 105768 626
rect 106812 598 106964 626
rect 107916 598 108160 626
rect 109020 598 109356 626
rect 110216 598 110552 626
rect 111320 598 111656 626
rect 112424 598 112852 626
rect 113620 598 114048 626
rect 114724 598 115244 626
rect 115828 598 116440 626
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 89364 462 89792 490
rect 90376 480 90404 598
rect 91572 480 91600 598
rect 92768 480 92796 598
rect 93964 480 93992 598
rect 95160 480 95188 598
rect 96264 480 96292 598
rect 97460 480 97488 598
rect 98656 480 98684 598
rect 99852 480 99880 598
rect 105740 480 105768 598
rect 106936 480 106964 598
rect 108132 480 108160 598
rect 109328 480 109356 598
rect 110524 480 110552 598
rect 111628 480 111656 598
rect 112824 480 112852 598
rect 114020 480 114048 598
rect 115216 480 115244 598
rect 116412 480 116440 598
rect 117424 598 117636 626
rect 118128 598 118832 626
rect 119324 598 119936 626
rect 117424 490 117452 598
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117024 462 117452 490
rect 117608 480 117636 598
rect 118804 480 118832 598
rect 119908 480 119936 598
rect 120920 598 121132 626
rect 121532 610 121868 626
rect 121532 604 121880 610
rect 121532 598 121828 604
rect 120920 490 120948 598
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 120428 462 120948 490
rect 121104 480 121132 598
rect 121828 546 121880 552
rect 122288 604 122340 610
rect 122288 546 122340 552
rect 123312 598 123524 626
rect 123832 610 124168 626
rect 124936 610 125272 626
rect 126132 610 126468 626
rect 127236 610 127572 626
rect 128340 610 128676 626
rect 123832 604 124180 610
rect 123832 598 124128 604
rect 122300 480 122328 546
rect 123312 490 123340 598
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 122728 462 123340 490
rect 123496 480 123524 598
rect 124128 546 124180 552
rect 124680 604 124732 610
rect 124936 604 125284 610
rect 124936 598 125232 604
rect 124680 546 124732 552
rect 125232 546 125284 552
rect 125876 604 125928 610
rect 126132 604 126480 610
rect 126132 598 126428 604
rect 125876 546 125928 552
rect 126428 546 126480 552
rect 126980 604 127032 610
rect 127236 604 127584 610
rect 127236 598 127532 604
rect 126980 546 127032 552
rect 127532 546 127584 552
rect 128176 604 128228 610
rect 128340 604 128688 610
rect 128340 598 128636 604
rect 128176 546 128228 552
rect 128636 546 128688 552
rect 129372 604 129424 610
rect 130640 598 130976 626
rect 131744 598 132080 626
rect 132940 620 133236 626
rect 134156 672 134208 678
rect 132940 614 133288 620
rect 132940 598 133276 614
rect 133892 610 134044 626
rect 134156 614 134208 620
rect 136180 672 136232 678
rect 137652 672 137704 678
rect 136232 620 136344 626
rect 136180 614 136344 620
rect 133880 604 134044 610
rect 129372 546 129424 552
rect 124692 480 124720 546
rect 125888 480 125916 546
rect 126992 480 127020 546
rect 128188 480 128216 546
rect 129384 480 129412 546
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 129832 128 129884 134
rect 129536 76 129832 82
rect 129536 70 129884 76
rect 130292 128 130344 134
rect 130538 82 130650 480
rect 130948 406 130976 598
rect 130936 400 130988 406
rect 130936 342 130988 348
rect 131734 354 131846 480
rect 132052 406 132080 598
rect 133932 598 134044 604
rect 133880 546 133932 552
rect 134168 480 134196 614
rect 135260 604 135312 610
rect 136192 598 136344 614
rect 137448 610 137600 626
rect 138756 672 138808 678
rect 137652 614 137704 620
rect 138552 620 138756 626
rect 140044 672 140096 678
rect 138552 614 138808 620
rect 136456 604 136508 610
rect 135260 546 135312 552
rect 137448 604 137612 610
rect 137448 598 137560 604
rect 136456 546 136508 552
rect 137560 546 137612 552
rect 134984 536 135036 542
rect 135036 484 135148 490
rect 131948 400 132000 406
rect 131734 348 131948 354
rect 131734 342 132000 348
rect 132040 400 132092 406
rect 132040 342 132092 348
rect 132930 354 133042 480
rect 133144 400 133196 406
rect 132930 348 133144 354
rect 132930 342 133196 348
rect 130344 76 130650 82
rect 130292 70 130650 76
rect 129536 54 129872 70
rect 130304 54 130650 70
rect 130538 -960 130650 54
rect 131734 326 131988 342
rect 132930 326 133184 342
rect 131734 -960 131846 326
rect 132930 -960 133042 326
rect 134126 -960 134238 480
rect 134984 478 135148 484
rect 135272 480 135300 546
rect 136468 480 136496 546
rect 137664 480 137692 614
rect 138552 598 138796 614
rect 139748 610 139992 626
rect 151360 672 151412 678
rect 142066 640 142122 649
rect 140044 614 140096 620
rect 138848 604 138900 610
rect 139748 604 140004 610
rect 139748 598 139952 604
rect 138848 546 138900 552
rect 139952 546 140004 552
rect 138860 480 138888 546
rect 140056 480 140084 614
rect 141240 604 141292 610
rect 141956 598 142066 626
rect 143446 640 143502 649
rect 142066 575 142122 584
rect 142264 598 142476 626
rect 143152 598 143446 626
rect 141240 546 141292 552
rect 141056 536 141108 542
rect 140852 484 141056 490
rect 134996 462 135148 478
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 140852 478 141108 484
rect 141252 480 141280 546
rect 142068 536 142120 542
rect 142264 490 142292 598
rect 142120 484 142292 490
rect 140852 462 141096 478
rect 141210 -960 141322 480
rect 142068 478 142292 484
rect 142448 480 142476 598
rect 144734 640 144790 649
rect 143446 575 143502 584
rect 143552 598 143764 626
rect 144256 610 144592 626
rect 144256 604 144604 610
rect 144256 598 144552 604
rect 143552 480 143580 598
rect 143736 513 143764 598
rect 145746 640 145802 649
rect 145452 598 145746 626
rect 144734 575 144790 584
rect 147126 640 147182 649
rect 146556 610 146892 626
rect 145746 575 145802 584
rect 145932 604 145984 610
rect 144552 546 144604 552
rect 143722 504 143778 513
rect 142080 462 142292 478
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144748 480 144776 575
rect 146556 604 146904 610
rect 146556 598 146852 604
rect 145932 546 145984 552
rect 148966 640 149022 649
rect 147126 575 147182 584
rect 148324 604 148376 610
rect 146852 546 146904 552
rect 145944 480 145972 546
rect 147140 480 147168 575
rect 148856 598 148966 626
rect 150622 640 150678 649
rect 148966 575 149022 584
rect 149348 598 149560 626
rect 148324 546 148376 552
rect 147770 504 147826 513
rect 143722 439 143778 448
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 147660 462 147770 490
rect 148336 480 148364 546
rect 149348 513 149376 598
rect 149334 504 149390 513
rect 147770 439 147826 448
rect 148294 -960 148406 480
rect 149532 480 149560 598
rect 151064 620 151360 626
rect 153016 672 153068 678
rect 151064 614 151412 620
rect 151818 640 151874 649
rect 151064 598 151400 614
rect 150622 575 150678 584
rect 152260 610 152596 626
rect 153660 672 153712 678
rect 153016 614 153068 620
rect 153364 620 153660 626
rect 155408 672 155460 678
rect 153364 614 153712 620
rect 152260 604 152608 610
rect 152260 598 152556 604
rect 151818 575 151874 584
rect 150254 504 150310 513
rect 149334 439 149390 448
rect 149490 -960 149602 480
rect 149960 462 150254 490
rect 150636 480 150664 575
rect 151832 480 151860 575
rect 152556 546 152608 552
rect 153028 480 153056 614
rect 153364 598 153700 614
rect 154468 610 154804 626
rect 162768 672 162820 678
rect 155408 614 155460 620
rect 154212 604 154264 610
rect 154468 604 154816 610
rect 154468 598 154764 604
rect 154212 546 154264 552
rect 154764 546 154816 552
rect 154224 480 154252 546
rect 155420 480 155448 614
rect 156768 610 157104 626
rect 156604 604 156656 610
rect 156768 604 157116 610
rect 156768 598 157064 604
rect 156604 546 156656 552
rect 157872 598 158208 626
rect 157064 546 157116 552
rect 156616 480 156644 546
rect 158180 542 158208 598
rect 158904 604 158956 610
rect 160172 598 160508 626
rect 161276 610 161612 626
rect 162472 620 162768 626
rect 164884 672 164936 678
rect 164790 640 164846 649
rect 162472 614 162820 620
rect 161276 604 161624 610
rect 161276 598 161572 604
rect 158904 546 158956 552
rect 158168 536 158220 542
rect 150254 439 150310 448
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 155960 128 156012 134
rect 155664 76 155960 82
rect 155664 70 156012 76
rect 155664 54 156000 70
rect 156574 -960 156686 480
rect 157524 128 157576 134
rect 157770 82 157882 480
rect 158168 478 158220 484
rect 158916 480 158944 546
rect 159732 536 159784 542
rect 157576 76 157882 82
rect 157524 70 157882 76
rect 157536 54 157882 70
rect 157770 -960 157882 54
rect 158874 -960 158986 480
rect 159732 478 159784 484
rect 159744 354 159772 478
rect 160070 354 160182 480
rect 160480 406 160508 598
rect 162472 598 162808 614
rect 163688 604 163740 610
rect 161572 546 161624 552
rect 164680 598 164790 626
rect 166080 672 166132 678
rect 164884 614 164936 620
rect 164790 575 164846 584
rect 163688 546 163740 552
rect 159744 326 160182 354
rect 160468 400 160520 406
rect 160468 342 160520 348
rect 159364 128 159416 134
rect 159068 76 159364 82
rect 159068 70 159416 76
rect 159068 54 159404 70
rect 160070 -960 160182 326
rect 161266 82 161378 480
rect 162462 354 162574 480
rect 163424 474 163576 490
rect 163700 480 163728 546
rect 164896 480 164924 614
rect 165876 610 166028 626
rect 167092 672 167144 678
rect 166080 614 166132 620
rect 166980 620 167092 626
rect 169576 672 169628 678
rect 167366 640 167422 649
rect 166980 614 167144 620
rect 165876 604 166040 610
rect 165876 598 165988 604
rect 165988 546 166040 552
rect 166092 480 166120 614
rect 166980 598 167132 614
rect 167196 598 167366 626
rect 167196 480 167224 598
rect 169482 640 169538 649
rect 167366 575 167422 584
rect 168380 604 168432 610
rect 169280 598 169482 626
rect 180892 672 180944 678
rect 171966 640 172022 649
rect 169576 614 169628 620
rect 169482 575 169538 584
rect 168380 546 168432 552
rect 168392 480 168420 546
rect 169588 480 169616 614
rect 170384 610 170720 626
rect 170384 604 170732 610
rect 170384 598 170680 604
rect 170680 546 170732 552
rect 170784 598 170996 626
rect 170784 480 170812 598
rect 163412 468 163576 474
rect 163464 462 163576 468
rect 163412 410 163464 416
rect 162676 400 162728 406
rect 162462 348 162676 354
rect 162462 342 162728 348
rect 162462 326 162716 342
rect 161480 128 161532 134
rect 161266 76 161480 82
rect 161266 70 161532 76
rect 161266 54 161520 70
rect 161266 -960 161378 54
rect 162462 -960 162574 326
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168194 368 168250 377
rect 168084 326 168194 354
rect 168194 303 168250 312
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 170968 377 170996 598
rect 172978 640 173034 649
rect 172684 598 172978 626
rect 171966 575 172022 584
rect 175462 640 175518 649
rect 172978 575 173034 584
rect 173164 604 173216 610
rect 171980 480 172008 575
rect 173164 546 173216 552
rect 174096 598 174308 626
rect 173176 480 173204 546
rect 173898 504 173954 513
rect 170954 368 171010 377
rect 171690 368 171746 377
rect 171488 326 171690 354
rect 170954 303 171010 312
rect 171690 303 171746 312
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 173788 462 173898 490
rect 174096 490 174124 598
rect 173898 439 173954 448
rect 174004 462 174124 490
rect 174280 480 174308 598
rect 176382 640 176438 649
rect 176088 598 176382 626
rect 175462 575 175518 584
rect 179050 640 179106 649
rect 176382 575 176438 584
rect 176672 598 176884 626
rect 175476 480 175504 575
rect 176672 480 176700 598
rect 176856 513 176884 598
rect 177684 598 177896 626
rect 176842 504 176898 513
rect 174004 377 174032 462
rect 173990 368 174046 377
rect 173990 303 174046 312
rect 174238 -960 174350 480
rect 175186 368 175242 377
rect 174984 326 175186 354
rect 175186 303 175242 312
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177486 504 177542 513
rect 177192 462 177486 490
rect 176842 439 176898 448
rect 177486 439 177542 448
rect 177684 377 177712 598
rect 177868 480 177896 598
rect 180246 640 180302 649
rect 179492 610 179828 626
rect 179492 604 179840 610
rect 179492 598 179788 604
rect 179050 575 179106 584
rect 179064 480 179092 575
rect 180596 620 180892 626
rect 183744 672 183796 678
rect 182086 640 182142 649
rect 180596 614 180944 620
rect 180596 598 180932 614
rect 181272 598 181484 626
rect 181792 598 182086 626
rect 180246 575 180302 584
rect 179788 546 179840 552
rect 180260 480 180288 575
rect 177670 368 177726 377
rect 177670 303 177726 312
rect 177826 -960 177938 480
rect 178682 368 178738 377
rect 178388 326 178682 354
rect 178682 303 178738 312
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181272 377 181300 598
rect 181456 480 181484 598
rect 182896 610 183232 626
rect 190000 672 190052 678
rect 183744 614 183796 620
rect 184938 640 184994 649
rect 182086 575 182142 584
rect 182548 604 182600 610
rect 182896 604 183244 610
rect 182896 598 183192 604
rect 182548 546 182600 552
rect 183192 546 183244 552
rect 182560 480 182588 546
rect 183756 480 183784 614
rect 184938 575 184994 584
rect 186136 604 186188 610
rect 184952 480 184980 575
rect 187404 598 187740 626
rect 188600 610 188844 626
rect 189704 620 190000 626
rect 193220 672 193272 678
rect 191102 640 191158 649
rect 189704 614 190052 620
rect 188600 604 188856 610
rect 188600 598 188804 604
rect 186136 546 186188 552
rect 186148 480 186176 546
rect 187712 542 187740 598
rect 189704 598 190040 614
rect 190808 598 191102 626
rect 192004 610 192340 626
rect 194324 672 194376 678
rect 193220 614 193272 620
rect 194212 620 194324 626
rect 197912 672 197964 678
rect 194212 614 194376 620
rect 194414 640 194470 649
rect 192004 604 192352 610
rect 192004 598 192300 604
rect 191102 575 191158 584
rect 188804 546 188856 552
rect 192300 546 192352 552
rect 187700 536 187752 542
rect 186594 504 186650 513
rect 181258 368 181314 377
rect 181258 303 181314 312
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184296 128 184348 134
rect 184000 76 184296 82
rect 184000 70 184348 76
rect 184000 54 184336 70
rect 184910 -960 185022 480
rect 185492 128 185544 134
rect 185196 76 185492 82
rect 185196 70 185544 76
rect 185196 54 185532 70
rect 186106 -960 186218 480
rect 186300 462 186594 490
rect 191012 536 191064 542
rect 186594 439 186650 448
rect 187302 218 187414 480
rect 187700 478 187752 484
rect 189906 504 189962 513
rect 186976 202 187414 218
rect 186964 196 187414 202
rect 187016 190 187414 196
rect 186964 138 187016 144
rect 187302 -960 187414 190
rect 188252 128 188304 134
rect 188498 82 188610 480
rect 188304 76 188610 82
rect 188252 70 188610 76
rect 188264 54 188610 70
rect 188498 -960 188610 54
rect 189694 218 189806 480
rect 189906 439 189962 448
rect 189920 218 189948 439
rect 189694 190 189948 218
rect 190798 354 190910 480
rect 191012 478 191064 484
rect 192208 536 192260 542
rect 191024 354 191052 478
rect 190798 326 191052 354
rect 191994 354 192106 480
rect 192208 478 192260 484
rect 192944 536 192996 542
rect 192996 484 193108 490
rect 192944 478 193108 484
rect 193232 480 193260 614
rect 194212 598 194364 614
rect 196714 640 196770 649
rect 194414 575 194470 584
rect 195612 604 195664 610
rect 194428 480 194456 575
rect 196512 598 196714 626
rect 196714 575 196770 584
rect 196820 610 196940 626
rect 213828 672 213880 678
rect 200302 640 200358 649
rect 197912 614 197964 620
rect 196820 604 196952 610
rect 196820 598 196900 604
rect 195612 546 195664 552
rect 195624 480 195652 546
rect 196820 480 196848 598
rect 196900 546 196952 552
rect 197924 480 197952 614
rect 198936 598 199148 626
rect 192220 354 192248 478
rect 192956 462 193108 478
rect 191994 326 192248 354
rect 189694 -960 189806 190
rect 190798 -960 190910 326
rect 191994 -960 192106 326
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195242 232 195298 241
rect 195298 190 195408 218
rect 195242 167 195298 176
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197726 368 197782 377
rect 197616 326 197726 354
rect 197726 303 197782 312
rect 197882 -960 197994 480
rect 198936 241 198964 598
rect 199120 480 199148 598
rect 200302 575 200358 584
rect 201498 640 201554 649
rect 203614 640 203670 649
rect 203320 598 203614 626
rect 201498 575 201554 584
rect 200316 480 200344 575
rect 201512 480 201540 575
rect 202524 564 202736 592
rect 207386 640 207442 649
rect 205620 610 205772 626
rect 205620 604 205784 610
rect 205620 598 205732 604
rect 203614 575 203670 584
rect 201866 504 201922 513
rect 198922 232 198978 241
rect 198922 167 198978 176
rect 198922 96 198978 105
rect 198812 54 198922 82
rect 198922 31 198978 40
rect 199078 -960 199190 480
rect 200026 368 200082 377
rect 199916 326 200026 354
rect 200026 303 200082 312
rect 200274 -960 200386 480
rect 201314 368 201370 377
rect 201112 326 201314 354
rect 201314 303 201370 312
rect 201470 -960 201582 480
rect 201866 439 201922 448
rect 201880 241 201908 439
rect 201866 232 201922 241
rect 202418 232 202474 241
rect 202216 190 202418 218
rect 201866 167 201922 176
rect 202418 167 202474 176
rect 202524 105 202552 564
rect 202708 480 202736 564
rect 203720 564 203932 592
rect 203720 513 203748 564
rect 203706 504 203762 513
rect 202510 96 202566 105
rect 202510 31 202566 40
rect 202666 -960 202778 480
rect 203904 480 203932 564
rect 204916 564 205128 592
rect 204810 504 204866 513
rect 203706 439 203762 448
rect 203862 -960 203974 480
rect 204516 462 204810 490
rect 204810 439 204866 448
rect 204916 377 204944 564
rect 205100 480 205128 564
rect 205732 546 205784 552
rect 206020 564 206232 592
rect 207386 575 207442 584
rect 208582 640 208638 649
rect 209318 640 209374 649
rect 209024 598 209318 626
rect 208582 575 208638 584
rect 213366 640 213422 649
rect 210128 610 210464 626
rect 209318 575 209374 584
rect 209780 604 209832 610
rect 204902 368 204958 377
rect 204902 303 204958 312
rect 205058 -960 205170 480
rect 206020 241 206048 564
rect 206204 480 206232 564
rect 207400 480 207428 575
rect 208214 504 208270 513
rect 206006 232 206062 241
rect 206006 167 206062 176
rect 206162 -960 206274 480
rect 206926 368 206982 377
rect 206724 326 206926 354
rect 206926 303 206982 312
rect 207358 -960 207470 480
rect 207920 462 208214 490
rect 208596 480 208624 575
rect 210128 604 210476 610
rect 210128 598 210424 604
rect 209780 546 209832 552
rect 210424 546 210476 552
rect 210804 598 211016 626
rect 211324 610 211660 626
rect 211324 604 211672 610
rect 211324 598 211620 604
rect 209792 480 209820 546
rect 208214 439 208270 448
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210804 377 210832 598
rect 210988 480 211016 598
rect 211620 546 211672 552
rect 212000 598 212212 626
rect 212000 513 212028 598
rect 211986 504 212042 513
rect 210790 368 210846 377
rect 210790 303 210846 312
rect 210946 -960 211058 480
rect 212184 480 212212 598
rect 213532 620 213828 626
rect 213532 614 213880 620
rect 215668 672 215720 678
rect 217968 672 218020 678
rect 215668 614 215720 620
rect 213532 598 213868 614
rect 214472 604 214524 610
rect 213366 575 213422 584
rect 211986 439 212042 448
rect 212142 -960 212254 480
rect 212428 474 212764 490
rect 213380 480 213408 575
rect 214472 546 214524 552
rect 214484 480 214512 546
rect 215680 480 215708 614
rect 216936 598 217272 626
rect 218428 672 218480 678
rect 218020 620 218054 626
rect 217968 614 218054 620
rect 217980 598 218054 614
rect 218132 620 218428 626
rect 222752 672 222804 678
rect 222474 640 222530 649
rect 218132 614 218480 620
rect 218132 598 218468 614
rect 219236 598 219572 626
rect 221536 610 221872 626
rect 216126 504 216182 513
rect 212428 468 212776 474
rect 212428 462 212724 468
rect 212724 410 212776 416
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 214728 66 215064 82
rect 214728 60 215076 66
rect 214728 54 215024 60
rect 215024 2 215076 8
rect 215638 -960 215750 480
rect 215832 462 216126 490
rect 216126 439 216182 448
rect 216588 468 216640 474
rect 216588 410 216640 416
rect 216600 354 216628 410
rect 216834 354 216946 480
rect 217244 377 217272 598
rect 218026 480 218054 598
rect 219544 542 219572 598
rect 220176 604 220228 610
rect 220176 546 220228 552
rect 220452 604 220504 610
rect 221536 604 221884 610
rect 221536 598 221832 604
rect 220452 546 220504 552
rect 222530 598 222640 626
rect 226340 672 226392 678
rect 222752 614 222804 620
rect 222474 575 222530 584
rect 221832 546 221884 552
rect 219532 536 219584 542
rect 220188 513 220216 546
rect 216600 326 216946 354
rect 216834 -960 216946 326
rect 217230 368 217286 377
rect 218026 326 218142 480
rect 217230 303 217286 312
rect 218030 -960 218142 326
rect 219226 82 219338 480
rect 219532 478 219584 484
rect 220174 504 220230 513
rect 220464 480 220492 546
rect 222764 480 222792 614
rect 223948 604 224000 610
rect 223948 546 224000 552
rect 225156 598 225368 626
rect 226044 610 226196 626
rect 231032 672 231084 678
rect 226340 614 226392 620
rect 227534 640 227590 649
rect 226044 604 226208 610
rect 226044 598 226156 604
rect 223578 504 223634 513
rect 220174 439 220230 448
rect 220176 400 220228 406
rect 220228 348 220340 354
rect 220176 342 220340 348
rect 220188 326 220340 342
rect 219226 66 219480 82
rect 219226 60 219492 66
rect 219226 54 219440 60
rect 219226 -960 219338 54
rect 219440 2 219492 8
rect 220422 -960 220534 480
rect 221526 354 221638 480
rect 221738 368 221794 377
rect 221526 326 221738 354
rect 221526 -960 221638 326
rect 221738 303 221794 312
rect 222722 -960 222834 480
rect 223634 462 223744 490
rect 223960 480 223988 546
rect 224776 536 224828 542
rect 224828 484 224940 490
rect 223578 439 223634 448
rect 223918 -960 224030 480
rect 224776 478 224940 484
rect 225156 480 225184 598
rect 224788 462 224940 478
rect 225114 -960 225226 480
rect 225340 406 225368 598
rect 226156 546 226208 552
rect 226352 480 226380 614
rect 227534 575 227590 584
rect 228730 640 228786 649
rect 230938 640 230994 649
rect 228730 575 228786 584
rect 229836 604 229888 610
rect 227548 480 227576 575
rect 228744 480 228772 575
rect 230644 598 230938 626
rect 234620 672 234672 678
rect 231032 614 231084 620
rect 230938 575 230994 584
rect 229836 546 229888 552
rect 229652 536 229704 542
rect 229448 484 229652 490
rect 225328 400 225380 406
rect 225328 342 225380 348
rect 226310 -960 226422 480
rect 227352 128 227404 134
rect 227148 76 227352 82
rect 227148 70 227404 76
rect 227148 54 227392 70
rect 227506 -960 227618 480
rect 228344 202 228588 218
rect 228344 196 228600 202
rect 228344 190 228548 196
rect 228548 138 228600 144
rect 228702 -960 228814 480
rect 229448 478 229704 484
rect 229848 480 229876 546
rect 231044 480 231072 614
rect 231748 610 231900 626
rect 231748 604 231912 610
rect 231748 598 231860 604
rect 231860 546 231912 552
rect 232056 598 232268 626
rect 229448 462 229692 478
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232056 134 232084 598
rect 232240 480 232268 598
rect 233252 598 233464 626
rect 235448 672 235500 678
rect 234620 614 234672 620
rect 235152 620 235448 626
rect 237748 672 237800 678
rect 235152 614 235500 620
rect 235814 640 235870 649
rect 233148 536 233200 542
rect 232852 484 233148 490
rect 232044 128 232096 134
rect 232044 70 232096 76
rect 232198 -960 232310 480
rect 232852 478 233200 484
rect 232852 462 233188 478
rect 233252 270 233280 598
rect 233436 480 233464 598
rect 233240 264 233292 270
rect 233240 206 233292 212
rect 233394 -960 233506 480
rect 234048 474 234384 490
rect 234632 480 234660 614
rect 235152 598 235488 614
rect 237452 620 237748 626
rect 242900 672 242952 678
rect 238850 640 238906 649
rect 237452 614 237800 620
rect 235814 575 235870 584
rect 237012 604 237064 610
rect 235828 480 235856 575
rect 237452 598 237788 614
rect 238116 604 238168 610
rect 237012 546 237064 552
rect 238556 598 238850 626
rect 240856 610 241192 626
rect 247960 672 248012 678
rect 242900 614 242952 620
rect 244094 640 244150 649
rect 238850 575 238906 584
rect 239312 604 239364 610
rect 238116 546 238168 552
rect 239312 546 239364 552
rect 240508 604 240560 610
rect 240856 604 241204 610
rect 240856 598 241152 604
rect 240508 546 240560 552
rect 241152 546 241204 552
rect 241532 564 241744 592
rect 237024 480 237052 546
rect 238128 480 238156 546
rect 239324 480 239352 546
rect 234048 468 234396 474
rect 234048 462 234344 468
rect 234344 410 234396 416
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236552 264 236604 270
rect 236256 212 236552 218
rect 236256 206 236604 212
rect 236256 190 236592 206
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 239660 474 239996 490
rect 240520 480 240548 546
rect 241532 490 241560 564
rect 239660 468 240008 474
rect 239660 462 239956 468
rect 239956 410 240008 416
rect 240478 -960 240590 480
rect 241440 462 241560 490
rect 241716 480 241744 564
rect 242912 480 242940 614
rect 246028 604 246080 610
rect 244094 575 244150 584
rect 243358 504 243414 513
rect 241440 270 241468 462
rect 241428 264 241480 270
rect 241428 206 241480 212
rect 241674 -960 241786 480
rect 241960 338 242296 354
rect 241960 332 242308 338
rect 241960 326 242256 332
rect 242256 274 242308 280
rect 242870 -960 242982 480
rect 243064 462 243358 490
rect 244108 480 244136 575
rect 244936 564 245240 592
rect 244556 536 244608 542
rect 244260 484 244556 490
rect 243358 439 243414 448
rect 244066 -960 244178 480
rect 244260 478 244608 484
rect 244260 462 244596 478
rect 244936 474 244964 564
rect 245212 480 245240 564
rect 246468 598 246804 626
rect 247664 620 247960 626
rect 253480 672 253532 678
rect 249062 640 249118 649
rect 247664 614 248012 620
rect 247664 598 248000 614
rect 248768 598 249062 626
rect 246028 546 246080 552
rect 244924 468 244976 474
rect 244924 410 244976 416
rect 245170 -960 245282 480
rect 245364 474 245700 490
rect 245364 468 245712 474
rect 245364 462 245660 468
rect 245660 410 245712 416
rect 246040 354 246068 546
rect 246366 354 246478 480
rect 246776 406 246804 598
rect 253276 610 253428 626
rect 257068 672 257120 678
rect 254674 640 254730 649
rect 253480 614 253532 620
rect 249062 575 249118 584
rect 249984 604 250036 610
rect 249984 546 250036 552
rect 251180 604 251232 610
rect 251180 546 251232 552
rect 252376 604 252428 610
rect 253276 604 253440 610
rect 253276 598 253388 604
rect 252376 546 252428 552
rect 253388 546 253440 552
rect 248970 504 249026 513
rect 246040 326 246478 354
rect 246764 400 246816 406
rect 247562 354 247674 480
rect 246764 342 246816 348
rect 247328 338 247674 354
rect 246366 -960 246478 326
rect 247316 332 247674 338
rect 247368 326 247674 332
rect 247316 274 247368 280
rect 247562 -960 247674 326
rect 248758 218 248870 480
rect 248970 439 249026 448
rect 249706 504 249762 513
rect 249762 462 249872 490
rect 249996 480 250024 546
rect 251192 480 251220 546
rect 252388 480 252416 546
rect 253492 480 253520 614
rect 254472 610 254624 626
rect 254472 604 254636 610
rect 254472 598 254584 604
rect 254674 575 254730 584
rect 255870 640 255926 649
rect 257068 614 257120 620
rect 257252 672 257304 678
rect 257252 614 257304 620
rect 258264 672 258316 678
rect 260656 672 260708 678
rect 258264 614 258316 620
rect 255870 575 255926 584
rect 254584 546 254636 552
rect 254688 480 254716 575
rect 255884 480 255912 575
rect 257080 480 257108 614
rect 249706 439 249762 448
rect 248984 218 249012 439
rect 248758 190 249012 218
rect 248758 -960 248870 190
rect 249954 -960 250066 480
rect 250916 338 251068 354
rect 250904 332 251068 338
rect 250956 326 251068 332
rect 250904 274 250956 280
rect 251150 -960 251262 480
rect 252008 128 252060 134
rect 252060 76 252172 82
rect 252008 70 252172 76
rect 252020 54 252172 70
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255688 264 255740 270
rect 255576 212 255688 218
rect 255576 206 255740 212
rect 255576 190 255728 206
rect 255842 -960 255954 480
rect 256772 338 256924 354
rect 256772 332 256936 338
rect 256772 326 256884 332
rect 256884 274 256936 280
rect 257038 -960 257150 480
rect 257264 134 257292 614
rect 257876 474 258028 490
rect 258276 480 258304 614
rect 260176 610 260512 626
rect 262680 672 262732 678
rect 260656 614 260708 620
rect 262384 620 262680 626
rect 268844 672 268896 678
rect 262384 614 262732 620
rect 263138 640 263194 649
rect 259460 604 259512 610
rect 260176 604 260524 610
rect 260176 598 260472 604
rect 259460 546 259512 552
rect 260472 546 260524 552
rect 257876 468 258040 474
rect 257876 462 257988 468
rect 257988 410 258040 416
rect 257252 128 257304 134
rect 257252 70 257304 76
rect 258234 -960 258346 480
rect 258980 474 259316 490
rect 259472 480 259500 546
rect 260668 480 260696 614
rect 262384 598 262720 614
rect 261588 564 261800 592
rect 261588 490 261616 564
rect 258980 468 259328 474
rect 258980 462 259276 468
rect 259276 410 259328 416
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261496 462 261616 490
rect 261772 480 261800 564
rect 262784 564 262996 592
rect 263138 575 263194 584
rect 264150 640 264206 649
rect 267278 640 267334 649
rect 266544 604 266596 610
rect 264150 575 264206 584
rect 261496 270 261524 462
rect 261484 264 261536 270
rect 261484 206 261536 212
rect 261576 264 261628 270
rect 261576 206 261628 212
rect 261588 82 261616 206
rect 261280 54 261616 82
rect 261730 -960 261842 480
rect 262784 338 262812 564
rect 262968 480 262996 564
rect 262772 332 262824 338
rect 262772 274 262824 280
rect 262926 -960 263038 480
rect 263152 406 263180 575
rect 263692 536 263744 542
rect 263580 484 263692 490
rect 263580 478 263744 484
rect 264164 480 264192 575
rect 265176 564 265388 592
rect 265176 490 265204 564
rect 263580 462 263732 478
rect 263140 400 263192 406
rect 263140 342 263192 348
rect 264122 -960 264234 480
rect 264992 474 265204 490
rect 265360 480 265388 564
rect 266984 598 267278 626
rect 267278 575 267334 584
rect 267568 598 267780 626
rect 272892 672 272944 678
rect 268844 614 268896 620
rect 266544 546 266596 552
rect 266556 480 266584 546
rect 264980 468 265204 474
rect 265032 462 265204 468
rect 264980 410 265032 416
rect 264684 202 264928 218
rect 264684 196 264940 202
rect 264684 190 264888 196
rect 264888 138 264940 144
rect 265318 -960 265430 480
rect 266084 128 266136 134
rect 265788 76 266084 82
rect 265788 70 266136 76
rect 265788 54 266124 70
rect 266514 -960 266626 480
rect 267568 270 267596 598
rect 267752 480 267780 598
rect 267556 264 267608 270
rect 267556 206 267608 212
rect 267710 -960 267822 480
rect 268088 474 268424 490
rect 268856 480 268884 614
rect 270040 604 270092 610
rect 270040 546 270092 552
rect 271064 598 271276 626
rect 270052 480 270080 546
rect 270500 536 270552 542
rect 270388 484 270500 490
rect 268088 468 268436 474
rect 268088 462 268384 468
rect 268384 410 268436 416
rect 268814 -960 268926 480
rect 269488 400 269540 406
rect 269192 348 269488 354
rect 269192 342 269540 348
rect 269192 326 269528 342
rect 270010 -960 270122 480
rect 270388 478 270552 484
rect 270388 462 270540 478
rect 271064 202 271092 598
rect 271248 480 271276 598
rect 272260 598 272472 626
rect 272596 620 272892 626
rect 285404 672 285456 678
rect 272596 614 272944 620
rect 273626 640 273682 649
rect 272596 598 272932 614
rect 271052 196 271104 202
rect 271052 138 271104 144
rect 271206 -960 271318 480
rect 272260 354 272288 598
rect 272444 480 272472 598
rect 275834 640 275890 649
rect 273792 610 274128 626
rect 273792 604 274140 610
rect 273792 598 274088 604
rect 273626 575 273682 584
rect 273640 480 273668 575
rect 274896 598 275232 626
rect 274088 546 274140 552
rect 275204 513 275232 598
rect 283102 640 283158 649
rect 275890 598 276000 626
rect 277196 598 277532 626
rect 278300 598 278636 626
rect 275834 575 275890 584
rect 276756 536 276808 542
rect 275190 504 275246 513
rect 271492 338 271828 354
rect 271492 332 271840 338
rect 271492 326 271788 332
rect 271788 274 271840 280
rect 272168 326 272288 354
rect 272168 134 272196 326
rect 272156 128 272208 134
rect 272156 70 272208 76
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274548 468 274600 474
rect 274548 410 274600 416
rect 274560 354 274588 410
rect 274794 354 274906 480
rect 275190 439 275246 448
rect 274560 326 274906 354
rect 274794 -960 274906 326
rect 275990 354 276102 480
rect 276756 478 276808 484
rect 276204 400 276256 406
rect 275990 348 276204 354
rect 275990 342 276256 348
rect 276768 354 276796 478
rect 277094 354 277206 480
rect 277504 474 277532 598
rect 277492 468 277544 474
rect 277492 410 277544 416
rect 275990 326 276244 342
rect 276768 326 277206 354
rect 275990 -960 276102 326
rect 277094 -960 277206 326
rect 278290 354 278402 480
rect 278608 406 278636 598
rect 279516 604 279568 610
rect 279516 546 279568 552
rect 280724 598 280936 626
rect 279528 480 279556 546
rect 280724 480 280752 598
rect 278596 400 278648 406
rect 278290 338 278544 354
rect 278596 342 278648 348
rect 279238 368 279294 377
rect 278290 332 278556 338
rect 278290 326 278504 332
rect 278290 -960 278402 326
rect 279294 326 279404 354
rect 279238 303 279294 312
rect 278504 274 278556 280
rect 279486 -960 279598 480
rect 280436 264 280488 270
rect 280488 212 280600 218
rect 280436 206 280600 212
rect 280448 190 280600 206
rect 280682 -960 280794 480
rect 280908 474 280936 598
rect 281920 598 282224 626
rect 281540 536 281592 542
rect 281592 484 281704 490
rect 281540 478 281704 484
rect 281920 480 281948 598
rect 282196 513 282224 598
rect 288992 672 289044 678
rect 285404 614 285456 620
rect 286598 640 286654 649
rect 283102 575 283158 584
rect 284300 604 284352 610
rect 282182 504 282238 513
rect 280896 468 280948 474
rect 281552 462 281704 478
rect 280896 410 280948 416
rect 281878 -960 281990 480
rect 283116 480 283144 575
rect 284300 546 284352 552
rect 282182 439 282238 448
rect 282808 202 282960 218
rect 282808 196 282972 202
rect 282808 190 282920 196
rect 282920 138 282972 144
rect 283074 -960 283186 480
rect 284004 474 284156 490
rect 284312 480 284340 546
rect 285218 504 285274 513
rect 284004 468 284168 474
rect 284004 462 284116 468
rect 284116 410 284168 416
rect 284270 -960 284382 480
rect 285108 462 285218 490
rect 285416 480 285444 614
rect 286598 575 286654 584
rect 287058 640 287114 649
rect 287058 575 287114 584
rect 287794 640 287850 649
rect 288512 610 288848 626
rect 291108 672 291160 678
rect 288992 614 289044 620
rect 288512 604 288860 610
rect 288512 598 288808 604
rect 287794 575 287850 584
rect 286612 480 286640 575
rect 285218 439 285274 448
rect 285374 -960 285486 480
rect 286416 128 286468 134
rect 286304 76 286416 82
rect 286304 70 286468 76
rect 286304 54 286456 70
rect 286570 -960 286682 480
rect 287072 270 287100 575
rect 287612 536 287664 542
rect 287408 484 287612 490
rect 287408 478 287664 484
rect 287808 480 287836 575
rect 288808 546 288860 552
rect 289004 480 289032 614
rect 290016 598 290228 626
rect 290812 620 291108 626
rect 293408 672 293460 678
rect 291566 640 291622 649
rect 290812 614 291160 620
rect 290812 598 291148 614
rect 291212 598 291424 626
rect 287408 462 287652 478
rect 287060 264 287112 270
rect 287060 206 287112 212
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290016 202 290044 598
rect 290200 480 290228 598
rect 290004 196 290056 202
rect 290004 138 290056 144
rect 289708 66 289860 82
rect 289708 60 289872 66
rect 289708 54 289820 60
rect 289820 2 289872 8
rect 290158 -960 290270 480
rect 291212 474 291240 598
rect 291396 480 291424 598
rect 291566 575 291622 584
rect 292592 598 292804 626
rect 293112 620 293408 626
rect 298468 672 298520 678
rect 293112 614 293460 620
rect 293682 640 293738 649
rect 293112 598 293448 614
rect 291200 468 291252 474
rect 291200 410 291252 416
rect 291354 -960 291466 480
rect 291580 134 291608 575
rect 292592 480 292620 598
rect 292776 513 292804 598
rect 293682 575 293738 584
rect 293866 640 293922 649
rect 293866 575 293922 584
rect 294878 640 294934 649
rect 294878 575 294934 584
rect 296076 604 296128 610
rect 292762 504 292818 513
rect 291916 202 292252 218
rect 291916 196 292264 202
rect 291916 190 292212 196
rect 292212 138 292264 144
rect 291568 128 291620 134
rect 291568 70 291620 76
rect 292550 -960 292662 480
rect 293696 480 293724 575
rect 293880 542 293908 575
rect 293868 536 293920 542
rect 292762 439 292818 448
rect 293654 -960 293766 480
rect 293868 478 293920 484
rect 294892 480 294920 575
rect 296076 546 296128 552
rect 297100 598 297312 626
rect 300768 672 300820 678
rect 298468 614 298520 620
rect 295616 536 295668 542
rect 295320 484 295616 490
rect 294512 400 294564 406
rect 294216 348 294512 354
rect 294216 342 294564 348
rect 294216 326 294552 342
rect 294850 -960 294962 480
rect 295320 478 295668 484
rect 296088 480 296116 546
rect 295320 462 295656 478
rect 296046 -960 296158 480
rect 297100 354 297128 598
rect 297284 480 297312 598
rect 298480 480 298508 614
rect 299492 598 299704 626
rect 301320 672 301372 678
rect 300768 614 300820 620
rect 301024 620 301320 626
rect 304724 672 304776 678
rect 301024 614 301372 620
rect 299492 490 299520 598
rect 297008 326 297128 354
rect 296812 264 296864 270
rect 296516 212 296812 218
rect 296516 206 296864 212
rect 296516 190 296852 206
rect 297008 66 297036 326
rect 296996 60 297048 66
rect 296996 2 297048 8
rect 297242 -960 297354 480
rect 297620 338 297956 354
rect 297620 332 297968 338
rect 297620 326 297916 332
rect 297916 274 297968 280
rect 298438 -960 298550 480
rect 299400 462 299520 490
rect 299676 480 299704 598
rect 299400 202 299428 462
rect 299388 196 299440 202
rect 299388 138 299440 144
rect 299020 128 299072 134
rect 298724 76 299020 82
rect 298724 70 299072 76
rect 298724 54 299060 70
rect 299634 -960 299746 480
rect 299920 474 300256 490
rect 300780 480 300808 614
rect 301024 598 301360 614
rect 303324 610 303660 626
rect 304428 620 304724 626
rect 307944 672 307996 678
rect 305826 640 305882 649
rect 304428 614 304776 620
rect 303160 604 303212 610
rect 301792 564 302004 592
rect 299920 468 300268 474
rect 299920 462 300216 468
rect 300216 410 300268 416
rect 300738 -960 300850 480
rect 301792 406 301820 564
rect 301976 480 302004 564
rect 303324 604 303672 610
rect 303324 598 303620 604
rect 303160 546 303212 552
rect 304428 598 304764 614
rect 305532 598 305826 626
rect 306728 598 307064 626
rect 307944 614 307996 620
rect 309968 672 310020 678
rect 318524 672 318576 678
rect 313830 640 313886 649
rect 310020 620 310132 626
rect 309968 614 310132 620
rect 305826 575 305882 584
rect 303620 546 303672 552
rect 303172 480 303200 546
rect 307036 513 307064 598
rect 307022 504 307078 513
rect 301780 400 301832 406
rect 301780 342 301832 348
rect 301934 -960 302046 480
rect 302424 400 302476 406
rect 302128 348 302424 354
rect 302128 342 302476 348
rect 302128 326 302464 342
rect 303130 -960 303242 480
rect 303988 264 304040 270
rect 304326 218 304438 480
rect 304040 212 304438 218
rect 303988 206 304438 212
rect 304000 190 304438 206
rect 304326 -960 304438 190
rect 305522 354 305634 480
rect 305522 338 305776 354
rect 305522 332 305788 338
rect 305522 326 305736 332
rect 305522 -960 305634 326
rect 305736 274 305788 280
rect 306718 82 306830 480
rect 307956 480 307984 614
rect 309048 604 309100 610
rect 309980 598 310132 614
rect 310244 604 310296 610
rect 309048 546 309100 552
rect 310244 546 310296 552
rect 311440 604 311492 610
rect 311440 546 311492 552
rect 312636 604 312688 610
rect 313830 575 313886 584
rect 315026 640 315082 649
rect 316590 640 316646 649
rect 315836 610 315988 626
rect 315836 604 316000 610
rect 315836 598 315948 604
rect 315026 575 315082 584
rect 312636 546 312688 552
rect 309060 480 309088 546
rect 310256 480 310284 546
rect 311452 480 311480 546
rect 312648 480 312676 546
rect 313844 480 313872 575
rect 315040 480 315068 575
rect 315948 546 316000 552
rect 316052 598 316264 626
rect 316052 542 316080 598
rect 316040 536 316092 542
rect 307022 439 307078 448
rect 307668 264 307720 270
rect 307720 212 307832 218
rect 307668 206 307832 212
rect 307680 190 307832 206
rect 306932 128 306984 134
rect 306718 76 306932 82
rect 306718 70 306984 76
rect 306718 54 306972 70
rect 306718 -960 306830 54
rect 307914 -960 308026 480
rect 308784 338 308936 354
rect 308772 332 308936 338
rect 308824 326 308936 332
rect 308772 274 308824 280
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311072 400 311124 406
rect 311124 348 311236 354
rect 311072 342 311236 348
rect 311084 326 311236 342
rect 311410 -960 311522 480
rect 312340 338 312492 354
rect 312340 332 312504 338
rect 312340 326 312452 332
rect 312452 274 312504 280
rect 312606 -960 312718 480
rect 313648 264 313700 270
rect 313536 212 313648 218
rect 313536 206 313700 212
rect 313536 190 313688 206
rect 313802 -960 313914 480
rect 314640 66 314792 82
rect 314640 60 314804 66
rect 314640 54 314752 60
rect 314752 2 314804 8
rect 314998 -960 315110 480
rect 316040 478 316092 484
rect 316236 480 316264 598
rect 317326 640 317382 649
rect 316940 610 317184 626
rect 316940 604 317196 610
rect 316940 598 317144 604
rect 316590 575 316646 584
rect 316194 -960 316306 480
rect 316604 474 316632 575
rect 318524 614 318576 620
rect 318708 672 318760 678
rect 319536 672 319588 678
rect 318708 614 318760 620
rect 319240 620 319536 626
rect 319240 614 319588 620
rect 326804 672 326856 678
rect 328460 672 328512 678
rect 326804 614 326856 620
rect 328256 620 328460 626
rect 331956 672 332008 678
rect 328256 614 328512 620
rect 331660 620 331956 626
rect 337476 672 337528 678
rect 334254 640 334310 649
rect 331660 614 332008 620
rect 317326 575 317382 584
rect 317144 546 317196 552
rect 317340 480 317368 575
rect 316592 468 316644 474
rect 316592 410 316644 416
rect 317298 -960 317410 480
rect 318044 474 318380 490
rect 318536 480 318564 614
rect 318044 468 318392 474
rect 318044 462 318340 468
rect 318340 410 318392 416
rect 318494 -960 318606 480
rect 318720 474 318748 614
rect 319240 598 319576 614
rect 325608 604 325660 610
rect 319732 564 319944 592
rect 319732 480 319760 564
rect 318708 468 318760 474
rect 318708 410 318760 416
rect 319690 -960 319802 480
rect 319916 406 319944 564
rect 320744 564 320956 592
rect 319904 400 319956 406
rect 319904 342 319956 348
rect 320744 338 320772 564
rect 320928 480 320956 564
rect 321848 564 322152 592
rect 321560 536 321612 542
rect 321448 484 321560 490
rect 320732 332 320784 338
rect 320732 274 320784 280
rect 320640 128 320692 134
rect 320344 76 320640 82
rect 320344 70 320692 76
rect 320344 54 320680 70
rect 320886 -960 320998 480
rect 321448 478 321612 484
rect 321448 462 321600 478
rect 321848 270 321876 564
rect 322124 480 322152 564
rect 323136 564 323348 592
rect 321836 264 321888 270
rect 321836 206 321888 212
rect 322082 -960 322194 480
rect 322848 264 322900 270
rect 322644 212 322848 218
rect 322644 206 322900 212
rect 322644 190 322888 206
rect 323136 82 323164 564
rect 323320 480 323348 564
rect 324240 564 324452 592
rect 322860 66 323164 82
rect 322848 60 323164 66
rect 322900 54 323164 60
rect 322848 2 322900 8
rect 323278 -960 323390 480
rect 324240 474 324268 564
rect 324424 480 324452 564
rect 325608 546 325660 552
rect 324228 468 324280 474
rect 324228 410 324280 416
rect 323748 202 324084 218
rect 323748 196 324096 202
rect 323748 190 324044 196
rect 324044 138 324096 144
rect 324382 -960 324494 480
rect 324852 474 325188 490
rect 325620 480 325648 546
rect 326816 480 326844 614
rect 328000 604 328052 610
rect 328256 598 328500 614
rect 330392 604 330444 610
rect 328000 546 328052 552
rect 329024 564 329236 592
rect 328012 480 328040 546
rect 324852 468 325200 474
rect 324852 462 325148 468
rect 325148 410 325200 416
rect 325578 -960 325690 480
rect 326342 368 326398 377
rect 326048 326 326342 354
rect 326342 303 326398 312
rect 326774 -960 326886 480
rect 327448 400 327500 406
rect 327152 348 327448 354
rect 327152 342 327500 348
rect 327152 326 327488 342
rect 327970 -960 328082 480
rect 329024 134 329052 564
rect 329208 480 329236 564
rect 331660 598 331996 614
rect 332520 598 332732 626
rect 333960 598 334254 626
rect 330392 546 330444 552
rect 330404 480 330432 546
rect 329012 128 329064 134
rect 329012 70 329064 76
rect 329166 -960 329278 480
rect 329748 128 329800 134
rect 329452 76 329748 82
rect 329452 70 329800 76
rect 329452 54 329788 70
rect 330362 -960 330474 480
rect 331220 264 331272 270
rect 331558 218 331670 480
rect 331272 212 331670 218
rect 331220 206 331670 212
rect 331232 190 331670 206
rect 332520 202 332548 598
rect 332704 480 332732 598
rect 335064 598 335400 626
rect 336260 598 336596 626
rect 342168 672 342220 678
rect 337476 614 337528 620
rect 334254 575 334310 584
rect 335372 513 335400 598
rect 335358 504 335414 513
rect 330556 66 330892 82
rect 330556 60 330904 66
rect 330556 54 330852 60
rect 330852 2 330904 8
rect 331558 -960 331670 190
rect 332508 196 332560 202
rect 332508 138 332560 144
rect 332662 -960 332774 480
rect 333612 468 333664 474
rect 333612 410 333664 416
rect 333624 354 333652 410
rect 333858 354 333970 480
rect 332856 338 333192 354
rect 332856 332 333204 338
rect 332856 326 333152 332
rect 333624 326 333970 354
rect 333152 274 333204 280
rect 333858 -960 333970 326
rect 335054 354 335166 480
rect 335358 439 335414 448
rect 335266 368 335322 377
rect 335054 326 335266 354
rect 335054 -960 335166 326
rect 335266 303 335322 312
rect 336250 354 336362 480
rect 336464 400 336516 406
rect 336250 348 336464 354
rect 336568 377 336596 598
rect 337488 480 337516 614
rect 341964 610 342116 626
rect 348240 672 348292 678
rect 342168 614 342220 620
rect 343362 640 343418 649
rect 338672 604 338724 610
rect 338672 546 338724 552
rect 339868 604 339920 610
rect 339868 546 339920 552
rect 340972 604 341024 610
rect 341964 604 342128 610
rect 341964 598 342076 604
rect 340972 546 341024 552
rect 342076 546 342128 552
rect 338684 480 338712 546
rect 339880 480 339908 546
rect 340984 480 341012 546
rect 342180 480 342208 614
rect 344558 640 344614 649
rect 344172 610 344508 626
rect 344172 604 344520 610
rect 344172 598 344468 604
rect 343362 575 343418 584
rect 343180 536 343232 542
rect 343068 484 343180 490
rect 336250 342 336516 348
rect 336554 368 336610 377
rect 336250 326 336504 342
rect 336250 -960 336362 326
rect 336554 303 336610 312
rect 337200 264 337252 270
rect 337252 212 337364 218
rect 337200 206 337364 212
rect 337212 190 337364 206
rect 337446 -960 337558 480
rect 338316 202 338468 218
rect 338304 196 338468 202
rect 338356 190 338468 196
rect 338304 138 338356 144
rect 338642 -960 338754 480
rect 339512 66 339664 82
rect 339500 60 339664 66
rect 339552 54 339664 60
rect 339500 2 339552 8
rect 339838 -960 339950 480
rect 340616 338 340768 354
rect 340604 332 340768 338
rect 340656 326 340768 332
rect 340604 274 340656 280
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343068 478 343232 484
rect 343376 480 343404 575
rect 344558 575 344614 584
rect 345754 640 345810 649
rect 345754 575 345810 584
rect 345938 640 345994 649
rect 345938 575 345994 584
rect 346950 640 347006 649
rect 346950 575 347006 584
rect 347778 640 347834 649
rect 347778 575 347834 584
rect 347884 598 348096 626
rect 348240 614 348292 620
rect 349068 672 349120 678
rect 351644 672 351696 678
rect 350446 640 350502 649
rect 349120 620 349292 626
rect 349068 614 349292 620
rect 344468 546 344520 552
rect 344572 480 344600 575
rect 345768 480 345796 575
rect 343068 462 343220 478
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345572 264 345624 270
rect 345368 212 345572 218
rect 345368 206 345624 212
rect 345368 190 345612 206
rect 345726 -960 345838 480
rect 345952 202 345980 575
rect 346472 474 346808 490
rect 346964 480 346992 575
rect 346472 468 346820 474
rect 346472 462 346768 468
rect 346768 410 346820 416
rect 345940 196 345992 202
rect 345940 138 345992 144
rect 346922 -960 347034 480
rect 347792 338 347820 575
rect 347780 332 347832 338
rect 347780 274 347832 280
rect 347884 218 347912 598
rect 348068 480 348096 598
rect 347424 202 347576 218
rect 347412 196 347576 202
rect 347464 190 347576 196
rect 347700 190 347912 218
rect 347412 138 347464 144
rect 347700 134 347728 190
rect 347688 128 347740 134
rect 347688 70 347740 76
rect 348026 -960 348138 480
rect 348252 66 348280 614
rect 349080 598 349292 614
rect 349264 480 349292 598
rect 352472 672 352524 678
rect 351644 614 351696 620
rect 351826 640 351882 649
rect 350446 575 350502 584
rect 350460 480 350488 575
rect 351656 480 351684 614
rect 352176 620 352472 626
rect 361948 672 362000 678
rect 352176 614 352524 620
rect 352838 640 352894 649
rect 352176 598 352512 614
rect 351826 575 351882 584
rect 352838 575 352894 584
rect 354036 604 354088 610
rect 351840 542 351868 575
rect 351828 536 351880 542
rect 349068 400 349120 406
rect 348772 348 349068 354
rect 348772 342 349120 348
rect 348772 326 349108 342
rect 348240 60 348292 66
rect 348240 2 348292 8
rect 349222 -960 349334 480
rect 350172 128 350224 134
rect 349876 76 350172 82
rect 349876 70 350224 76
rect 349876 54 350212 70
rect 350418 -960 350530 480
rect 350980 338 351316 354
rect 350980 332 351328 338
rect 350980 326 351276 332
rect 351276 274 351328 280
rect 351614 -960 351726 480
rect 351828 478 351880 484
rect 352852 480 352880 575
rect 354036 546 354088 552
rect 354968 598 355272 626
rect 354048 480 354076 546
rect 354680 536 354732 542
rect 354384 484 354680 490
rect 352810 -960 352922 480
rect 353280 66 353616 82
rect 353280 60 353628 66
rect 353280 54 353576 60
rect 353576 2 353628 8
rect 354006 -960 354118 480
rect 354384 478 354732 484
rect 354384 462 354720 478
rect 354968 270 354996 598
rect 355244 480 355272 598
rect 356336 604 356388 610
rect 356336 546 356388 552
rect 357360 598 357572 626
rect 356348 480 356376 546
rect 354956 264 355008 270
rect 354956 206 355008 212
rect 355202 -960 355314 480
rect 355876 264 355928 270
rect 355580 212 355876 218
rect 355580 206 355928 212
rect 355580 190 355916 206
rect 356306 -960 356418 480
rect 356684 474 357020 490
rect 356684 468 357032 474
rect 356684 462 356980 468
rect 356980 410 357032 416
rect 357360 202 357388 598
rect 357544 480 357572 598
rect 358728 604 358780 610
rect 361192 598 361528 626
rect 369584 672 369636 678
rect 364430 640 364486 649
rect 361948 614 362000 620
rect 358728 546 358780 552
rect 359752 564 359964 592
rect 358740 480 358768 546
rect 359280 536 359332 542
rect 358984 484 359280 490
rect 357348 196 357400 202
rect 357348 138 357400 144
rect 357502 -960 357614 480
rect 357788 202 358124 218
rect 357788 196 358136 202
rect 357788 190 358084 196
rect 358084 138 358136 144
rect 358698 -960 358810 480
rect 358984 478 359332 484
rect 358984 462 359320 478
rect 359752 134 359780 564
rect 359936 480 359964 564
rect 359740 128 359792 134
rect 359740 70 359792 76
rect 359894 -960 360006 480
rect 360088 474 360424 490
rect 360088 468 360436 474
rect 360088 462 360384 468
rect 360384 410 360436 416
rect 361090 354 361202 480
rect 360856 338 361202 354
rect 360844 332 361202 338
rect 360896 326 361202 332
rect 360844 274 360896 280
rect 361090 -960 361202 326
rect 361500 202 361528 598
rect 361960 354 361988 614
rect 362388 598 362724 626
rect 363492 598 363828 626
rect 362696 542 362724 598
rect 362684 536 362736 542
rect 362286 354 362398 480
rect 362684 478 362736 484
rect 361960 326 362398 354
rect 361488 196 361540 202
rect 361488 138 361540 144
rect 362286 -960 362398 326
rect 363482 218 363594 480
rect 363800 338 363828 598
rect 364486 598 364596 626
rect 364800 604 364852 610
rect 364430 575 364486 584
rect 365792 598 366128 626
rect 364800 546 364852 552
rect 364586 354 364698 480
rect 364812 354 364840 546
rect 366100 513 366128 598
rect 367020 598 367324 626
rect 369196 610 369348 626
rect 369412 620 369584 626
rect 370412 672 370464 678
rect 369412 614 369636 620
rect 370300 620 370412 626
rect 370688 672 370740 678
rect 370300 614 370464 620
rect 370608 620 370688 626
rect 371608 672 371660 678
rect 370608 614 370740 620
rect 371496 620 371608 626
rect 375196 672 375248 678
rect 371496 614 371660 620
rect 366086 504 366142 513
rect 363788 332 363840 338
rect 363788 274 363840 280
rect 364586 326 364840 354
rect 363482 190 363736 218
rect 363482 -960 363594 190
rect 363708 66 363736 190
rect 363696 60 363748 66
rect 363696 2 363748 8
rect 364586 -960 364698 326
rect 365782 218 365894 480
rect 366744 474 366896 490
rect 367020 480 367048 598
rect 366086 439 366142 448
rect 366732 468 366896 474
rect 366784 462 366896 468
rect 366732 410 366784 416
rect 365996 264 366048 270
rect 365782 212 365996 218
rect 365782 206 366048 212
rect 365782 190 366036 206
rect 365782 -960 365894 190
rect 366978 -960 367090 480
rect 367296 406 367324 598
rect 368204 604 368256 610
rect 369196 604 369360 610
rect 369196 598 369308 604
rect 368204 546 368256 552
rect 369308 546 369360 552
rect 369412 598 369624 614
rect 370300 598 370452 614
rect 370608 598 370728 614
rect 371496 598 371648 614
rect 371712 598 372016 626
rect 368216 480 368244 546
rect 369412 480 369440 598
rect 370608 480 370636 598
rect 371712 480 371740 598
rect 367284 400 367336 406
rect 367284 342 367336 348
rect 367836 128 367888 134
rect 367888 76 368000 82
rect 367836 70 368000 76
rect 367848 54 368000 70
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 371988 202 372016 598
rect 372908 598 373120 626
rect 372908 480 372936 598
rect 373092 542 373120 598
rect 374104 598 374316 626
rect 374900 620 375196 626
rect 377404 672 377456 678
rect 374900 614 375248 620
rect 375286 640 375342 649
rect 374900 598 375236 614
rect 373080 536 373132 542
rect 372436 400 372488 406
rect 372488 348 372600 354
rect 372436 342 372600 348
rect 372448 326 372600 342
rect 371976 196 372028 202
rect 371976 138 372028 144
rect 372866 -960 372978 480
rect 373080 478 373132 484
rect 373704 474 373948 490
rect 374104 480 374132 598
rect 373704 468 373960 474
rect 373704 462 373908 468
rect 373908 410 373960 416
rect 374062 -960 374174 480
rect 374288 338 374316 598
rect 375286 575 375342 584
rect 376482 640 376538 649
rect 377108 620 377404 626
rect 382372 672 382424 678
rect 377108 614 377456 620
rect 377108 598 377444 614
rect 377508 598 377720 626
rect 376482 575 376538 584
rect 375300 480 375328 575
rect 376496 480 376524 575
rect 377404 536 377456 542
rect 377508 490 377536 598
rect 377456 484 377536 490
rect 374276 332 374328 338
rect 374276 274 374328 280
rect 375258 -960 375370 480
rect 376004 66 376340 82
rect 376004 60 376352 66
rect 376004 54 376300 60
rect 376300 2 376352 8
rect 376454 -960 376566 480
rect 377404 478 377536 484
rect 377692 480 377720 598
rect 378704 598 378916 626
rect 382372 614 382424 620
rect 385960 672 386012 678
rect 388812 672 388864 678
rect 385960 614 386012 620
rect 388516 620 388812 626
rect 396540 672 396592 678
rect 393778 640 393834 649
rect 388516 614 388864 620
rect 377416 462 377536 478
rect 377650 -960 377762 480
rect 378600 400 378652 406
rect 378304 348 378600 354
rect 378304 342 378652 348
rect 378304 326 378640 342
rect 378704 134 378732 598
rect 378888 480 378916 598
rect 379980 604 380032 610
rect 379980 546 380032 552
rect 381176 604 381228 610
rect 381176 546 381228 552
rect 379992 480 380020 546
rect 381188 480 381216 546
rect 382384 480 382412 614
rect 383304 564 383608 592
rect 378692 128 378744 134
rect 378692 70 378744 76
rect 378846 -960 378958 480
rect 379520 128 379572 134
rect 379408 76 379520 82
rect 379408 70 379572 76
rect 379408 54 379560 70
rect 379950 -960 380062 480
rect 380512 202 380848 218
rect 380512 196 380860 202
rect 380512 190 380808 196
rect 380808 138 380860 144
rect 381146 -960 381258 480
rect 382004 264 382056 270
rect 381708 212 382004 218
rect 381708 206 382056 212
rect 381708 190 382044 206
rect 382342 -960 382454 480
rect 383106 368 383162 377
rect 382812 326 383106 354
rect 383304 338 383332 564
rect 383580 480 383608 564
rect 384592 564 384804 592
rect 384210 504 384266 513
rect 383106 303 383162 312
rect 383292 332 383344 338
rect 383292 274 383344 280
rect 383538 -960 383650 480
rect 383916 462 384210 490
rect 384592 474 384620 564
rect 384776 480 384804 564
rect 385408 536 385460 542
rect 385112 484 385408 490
rect 384210 439 384266 448
rect 384580 468 384632 474
rect 384580 410 384632 416
rect 384734 -960 384846 480
rect 385112 478 385460 484
rect 385972 480 386000 614
rect 388260 604 388312 610
rect 386984 564 387196 592
rect 386984 490 387012 564
rect 385112 462 385448 478
rect 385774 232 385830 241
rect 385774 167 385776 176
rect 385828 167 385830 176
rect 385776 138 385828 144
rect 385930 -960 386042 480
rect 386800 462 387012 490
rect 387168 480 387196 564
rect 388516 598 388852 614
rect 389192 598 389496 626
rect 390724 610 391060 626
rect 390724 604 391072 610
rect 390724 598 391020 604
rect 388260 546 388312 552
rect 388272 480 388300 546
rect 386216 202 386552 218
rect 386216 196 386564 202
rect 386216 190 386512 196
rect 386512 138 386564 144
rect 386800 66 386828 462
rect 386970 368 387026 377
rect 386970 303 386972 312
rect 387024 303 387026 312
rect 386972 274 387024 280
rect 386788 60 386840 66
rect 386788 2 386840 8
rect 387126 -960 387238 480
rect 387320 66 387656 82
rect 387320 60 387668 66
rect 387320 54 387616 60
rect 387616 2 387668 8
rect 388230 -960 388342 480
rect 389192 406 389220 598
rect 389468 480 389496 598
rect 391920 598 392256 626
rect 393024 598 393360 626
rect 391020 546 391072 552
rect 389824 536 389876 542
rect 389822 504 389824 513
rect 392228 513 392256 598
rect 389876 504 389878 513
rect 389180 400 389232 406
rect 389180 342 389232 348
rect 389426 -960 389538 480
rect 392214 504 392270 513
rect 389822 439 389878 448
rect 389916 400 389968 406
rect 389620 348 389916 354
rect 389620 342 389968 348
rect 389620 326 389956 342
rect 390284 128 390336 134
rect 390622 82 390734 480
rect 391570 232 391626 241
rect 391818 218 391930 480
rect 392214 439 392270 448
rect 391626 190 391930 218
rect 391570 167 391626 176
rect 390336 76 390734 82
rect 390284 70 390734 76
rect 390296 54 390734 70
rect 390622 -960 390734 54
rect 391818 -960 391930 190
rect 393014 218 393126 480
rect 393332 474 393360 598
rect 393778 575 393834 584
rect 394252 598 394464 626
rect 395324 598 395660 626
rect 400036 672 400088 678
rect 396540 614 396592 620
rect 393320 468 393372 474
rect 393320 410 393372 416
rect 393792 406 393820 575
rect 394252 480 394280 598
rect 393780 400 393832 406
rect 393780 342 393832 348
rect 393228 264 393280 270
rect 393014 212 393228 218
rect 393014 206 393280 212
rect 393964 264 394016 270
rect 394016 212 394128 218
rect 393964 206 394128 212
rect 393014 190 393268 206
rect 393976 190 394128 206
rect 393014 -960 393126 190
rect 394210 -960 394322 480
rect 394436 338 394464 598
rect 394424 332 394476 338
rect 394424 274 394476 280
rect 395314 82 395426 480
rect 395632 474 395660 598
rect 396552 480 396580 614
rect 398728 610 398880 626
rect 399832 620 400036 626
rect 402520 672 402572 678
rect 399832 614 400088 620
rect 401322 640 401378 649
rect 397736 604 397788 610
rect 398728 604 398892 610
rect 398728 598 398840 604
rect 397736 546 397788 552
rect 399832 598 400076 614
rect 400220 604 400272 610
rect 398840 546 398892 552
rect 398944 564 399156 592
rect 397748 480 397776 546
rect 398944 480 398972 564
rect 395620 468 395672 474
rect 395620 410 395672 416
rect 395528 128 395580 134
rect 395314 76 395528 82
rect 395314 70 395580 76
rect 396264 128 396316 134
rect 396316 76 396428 82
rect 396264 70 396428 76
rect 395314 54 395568 70
rect 396276 54 396428 70
rect 395314 -960 395426 54
rect 396510 -960 396622 480
rect 397460 264 397512 270
rect 397512 212 397624 218
rect 397460 206 397624 212
rect 397472 190 397624 206
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 399128 66 399156 564
rect 400140 564 400220 592
rect 400140 480 400168 564
rect 400220 546 400272 552
rect 400312 604 400364 610
rect 403440 672 403492 678
rect 402520 614 402572 620
rect 403236 620 403440 626
rect 409236 672 409288 678
rect 403236 614 403492 620
rect 401322 575 401378 584
rect 400312 546 400364 552
rect 400324 513 400352 546
rect 400310 504 400366 513
rect 399116 60 399168 66
rect 399116 2 399168 8
rect 400098 -960 400210 480
rect 401336 480 401364 575
rect 402532 480 402560 614
rect 403236 598 403480 614
rect 403544 610 403664 626
rect 403532 604 403664 610
rect 403584 598 403664 604
rect 404432 610 404768 626
rect 405536 610 405688 626
rect 404432 604 404780 610
rect 404432 598 404728 604
rect 403532 546 403584 552
rect 403636 480 403664 598
rect 404728 546 404780 552
rect 404820 604 404872 610
rect 405536 604 405700 610
rect 405536 598 405648 604
rect 404820 546 404872 552
rect 405648 546 405700 552
rect 405752 598 406056 626
rect 404832 480 404860 546
rect 400310 439 400366 448
rect 401140 400 401192 406
rect 401028 348 401140 354
rect 401028 342 401192 348
rect 401028 326 401180 342
rect 401294 -960 401406 480
rect 402336 128 402388 134
rect 402132 76 402336 82
rect 402132 70 402388 76
rect 402132 54 402376 70
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405752 474 405780 598
rect 406028 480 406056 598
rect 408236 598 408448 626
rect 408940 620 409236 626
rect 410800 672 410852 678
rect 408940 614 409288 620
rect 408940 598 409276 614
rect 409432 598 409644 626
rect 416688 672 416740 678
rect 410800 614 410852 620
rect 407040 564 407252 592
rect 405740 468 405792 474
rect 405740 410 405792 416
rect 405986 -960 406098 480
rect 406640 338 406976 354
rect 406640 332 406988 338
rect 406640 326 406936 332
rect 406936 274 406988 280
rect 407040 66 407068 564
rect 407224 480 407252 564
rect 408236 542 408264 598
rect 408224 536 408276 542
rect 407028 60 407080 66
rect 407028 2 407080 8
rect 407182 -960 407294 480
rect 407836 474 408172 490
rect 408224 478 408276 484
rect 408420 480 408448 598
rect 407836 468 408184 474
rect 407836 462 408132 468
rect 408132 410 408184 416
rect 408378 -960 408490 480
rect 409432 202 409460 598
rect 409616 480 409644 598
rect 410340 536 410392 542
rect 410044 484 410340 490
rect 409420 196 409472 202
rect 409420 138 409472 144
rect 409574 -960 409686 480
rect 410044 478 410392 484
rect 410812 480 410840 614
rect 411732 598 411944 626
rect 412344 610 412680 626
rect 412344 604 412692 610
rect 412344 598 412640 604
rect 410044 462 410380 478
rect 410770 -960 410882 480
rect 411732 406 411760 598
rect 411916 480 411944 598
rect 412640 546 412692 552
rect 412928 598 413140 626
rect 413448 610 413784 626
rect 418344 672 418396 678
rect 416688 614 416740 620
rect 418048 620 418344 626
rect 421012 672 421064 678
rect 418048 614 418396 620
rect 413448 604 413796 610
rect 413448 598 413744 604
rect 411720 400 411772 406
rect 411720 342 411772 348
rect 411240 202 411576 218
rect 411240 196 411588 202
rect 411240 190 411536 196
rect 411536 138 411588 144
rect 411874 -960 411986 480
rect 412928 270 412956 598
rect 413112 480 413140 598
rect 413744 546 413796 552
rect 414296 604 414348 610
rect 414296 546 414348 552
rect 415492 604 415544 610
rect 415492 546 415544 552
rect 414308 480 414336 546
rect 415504 480 415532 546
rect 416700 480 416728 614
rect 417884 604 417936 610
rect 418048 598 418384 614
rect 418816 598 419028 626
rect 420256 598 420592 626
rect 421104 672 421156 678
rect 421012 614 421064 620
rect 421102 640 421104 649
rect 423496 672 423548 678
rect 421156 640 421158 649
rect 417884 546 417936 552
rect 417146 504 417202 513
rect 412916 264 412968 270
rect 412916 206 412968 212
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 414644 66 414980 82
rect 414644 60 414992 66
rect 414644 54 414940 60
rect 414940 2 414992 8
rect 415462 -960 415574 480
rect 415748 338 416084 354
rect 415748 332 416096 338
rect 415748 326 416044 332
rect 416044 274 416096 280
rect 416658 -960 416770 480
rect 416852 462 417146 490
rect 417896 480 417924 546
rect 417146 439 417202 448
rect 417854 -960 417966 480
rect 418816 270 418844 598
rect 419000 480 419028 598
rect 418804 264 418856 270
rect 418804 206 418856 212
rect 418958 -960 419070 480
rect 419908 468 419960 474
rect 419908 410 419960 416
rect 419920 354 419948 410
rect 420154 354 420266 480
rect 420564 474 420592 598
rect 420552 468 420604 474
rect 420552 410 420604 416
rect 419920 326 420266 354
rect 421024 354 421052 614
rect 421452 598 421788 626
rect 421102 575 421158 584
rect 421350 354 421462 480
rect 421024 326 421462 354
rect 419448 128 419500 134
rect 419152 76 419448 82
rect 419152 70 419500 76
rect 419152 54 419488 70
rect 420154 -960 420266 326
rect 421350 -960 421462 326
rect 421760 270 421788 598
rect 422404 598 422556 626
rect 425520 672 425572 678
rect 424966 640 425022 649
rect 423548 620 423660 626
rect 423496 614 423660 620
rect 423508 598 423660 614
rect 423772 604 423824 610
rect 421748 264 421800 270
rect 421748 206 421800 212
rect 422404 202 422432 598
rect 424966 575 425022 584
rect 425518 640 425520 649
rect 425612 672 425664 678
rect 425572 640 425574 649
rect 430856 672 430908 678
rect 426162 640 426218 649
rect 425664 620 425960 626
rect 425612 614 425960 620
rect 425624 598 425960 614
rect 425518 575 425574 584
rect 429658 640 429714 649
rect 428260 610 428412 626
rect 426162 575 426218 584
rect 427268 604 427320 610
rect 423772 546 423824 552
rect 422760 536 422812 542
rect 422546 354 422658 480
rect 422760 478 422812 484
rect 423784 480 423812 546
rect 424980 480 425008 575
rect 426176 480 426204 575
rect 428260 604 428424 610
rect 428260 598 428372 604
rect 427268 546 427320 552
rect 428372 546 428424 552
rect 428476 598 428688 626
rect 429364 610 429516 626
rect 429364 604 429528 610
rect 429364 598 429476 604
rect 427280 480 427308 546
rect 428476 480 428504 598
rect 422772 354 422800 478
rect 422546 326 422800 354
rect 422392 196 422444 202
rect 422392 138 422444 144
rect 422546 -960 422658 326
rect 423742 -960 423854 480
rect 424692 400 424744 406
rect 424744 348 424856 354
rect 424692 342 424856 348
rect 424704 326 424856 342
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427004 66 427156 82
rect 426992 60 427156 66
rect 427044 54 427156 60
rect 426992 2 427044 8
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 428660 338 428688 598
rect 431868 672 431920 678
rect 430856 614 430908 620
rect 431664 620 431868 626
rect 431664 614 431920 620
rect 432052 672 432104 678
rect 436468 672 436520 678
rect 432052 614 432104 620
rect 429658 575 429714 584
rect 429476 546 429528 552
rect 429672 480 429700 575
rect 428648 332 428700 338
rect 428648 274 428700 280
rect 429630 -960 429742 480
rect 430560 474 430712 490
rect 430868 480 430896 614
rect 431664 598 431908 614
rect 432064 480 432092 614
rect 433248 604 433300 610
rect 433248 546 433300 552
rect 434272 598 434484 626
rect 436172 620 436468 626
rect 436172 614 436520 620
rect 436744 672 436796 678
rect 437480 672 437532 678
rect 436744 614 436796 620
rect 437368 620 437480 626
rect 439872 672 439924 678
rect 437368 614 437532 620
rect 430560 468 430724 474
rect 430560 462 430672 468
rect 430672 410 430724 416
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 432768 474 433104 490
rect 433260 480 433288 546
rect 432768 468 433116 474
rect 432768 462 433064 468
rect 433064 410 433116 416
rect 433218 -960 433330 480
rect 434272 354 434300 598
rect 434456 480 434484 598
rect 434720 604 434772 610
rect 434720 546 434772 552
rect 435548 604 435600 610
rect 436172 598 436508 614
rect 435548 546 435600 552
rect 434088 326 434300 354
rect 434088 270 434116 326
rect 434076 264 434128 270
rect 434076 206 434128 212
rect 434260 128 434312 134
rect 433964 76 434260 82
rect 433964 70 434312 76
rect 433964 54 434300 70
rect 434414 -960 434526 480
rect 434732 202 434760 546
rect 435560 480 435588 546
rect 436756 480 436784 614
rect 437368 598 437520 614
rect 437768 598 437980 626
rect 439576 620 439872 626
rect 449992 672 450044 678
rect 445574 640 445630 649
rect 439576 614 439924 620
rect 435068 202 435404 218
rect 434720 196 434772 202
rect 435068 196 435416 202
rect 435068 190 435364 196
rect 434720 138 434772 144
rect 435364 138 435416 144
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437768 354 437796 598
rect 437952 480 437980 598
rect 439136 604 439188 610
rect 439576 598 439912 614
rect 440160 598 440372 626
rect 444176 610 444512 626
rect 439136 546 439188 552
rect 438768 536 438820 542
rect 438472 484 438768 490
rect 437584 338 437796 354
rect 437572 332 437796 338
rect 437624 326 437796 332
rect 437572 274 437624 280
rect 437910 -960 438022 480
rect 438472 478 438820 484
rect 439148 480 439176 546
rect 438472 462 438808 478
rect 439106 -960 439218 480
rect 440160 66 440188 598
rect 440344 480 440372 598
rect 441528 604 441580 610
rect 441528 546 441580 552
rect 442632 604 442684 610
rect 444176 604 444524 610
rect 444176 598 444472 604
rect 442632 546 442684 552
rect 443656 564 443868 592
rect 441540 480 441568 546
rect 442644 480 442672 546
rect 440148 60 440200 66
rect 440148 2 440200 8
rect 440302 -960 440414 480
rect 440772 66 441108 82
rect 440772 60 441120 66
rect 440772 54 441068 60
rect 441068 2 441120 8
rect 441498 -960 441610 480
rect 441876 338 442212 354
rect 441876 332 442224 338
rect 441876 326 442172 332
rect 442172 274 442224 280
rect 442602 -960 442714 480
rect 443656 406 443684 564
rect 443840 480 443868 564
rect 444472 546 444524 552
rect 445024 604 445076 610
rect 445280 598 445574 626
rect 449912 632 449992 660
rect 449912 626 449940 632
rect 446384 610 446720 626
rect 445574 575 445630 584
rect 446220 604 446272 610
rect 445024 546 445076 552
rect 446384 604 446732 610
rect 446384 598 446680 604
rect 446220 546 446272 552
rect 446680 546 446732 552
rect 447244 598 447456 626
rect 447580 610 447916 626
rect 447580 604 447928 610
rect 447580 598 447876 604
rect 445036 480 445064 546
rect 446232 480 446260 546
rect 447244 490 447272 598
rect 443644 400 443696 406
rect 443644 342 443696 348
rect 443276 264 443328 270
rect 442980 212 443276 218
rect 442980 206 443328 212
rect 442980 190 443316 206
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447152 462 447272 490
rect 447428 480 447456 598
rect 448684 598 449020 626
rect 447876 546 447928 552
rect 447152 134 447180 462
rect 447140 128 447192 134
rect 447140 70 447192 76
rect 447386 -960 447498 480
rect 448244 196 448296 202
rect 448244 138 448296 144
rect 448256 82 448284 138
rect 448582 82 448694 480
rect 448992 202 449020 598
rect 449636 598 449788 626
rect 449866 598 449940 626
rect 453580 672 453632 678
rect 449992 614 450044 620
rect 450984 598 451320 626
rect 452088 598 452424 626
rect 453284 620 453580 626
rect 453284 614 453632 620
rect 454224 672 454276 678
rect 454500 672 454552 678
rect 454276 620 454388 626
rect 454224 614 454388 620
rect 456892 672 456944 678
rect 454500 614 454552 620
rect 453284 598 453620 614
rect 454236 598 454388 614
rect 449636 406 449664 598
rect 449866 480 449894 598
rect 449624 400 449676 406
rect 449624 342 449676 348
rect 449778 326 449894 480
rect 450636 468 450688 474
rect 450636 410 450688 416
rect 450648 354 450676 410
rect 450882 354 450994 480
rect 450648 326 450994 354
rect 451292 338 451320 598
rect 452078 354 452190 480
rect 452396 406 452424 598
rect 454512 480 454540 614
rect 455708 598 455920 626
rect 460388 672 460440 678
rect 456892 614 456944 620
rect 459190 640 459246 649
rect 455708 480 455736 598
rect 455892 542 455920 598
rect 455880 536 455932 542
rect 452292 400 452344 406
rect 452078 348 452292 354
rect 452078 342 452344 348
rect 452384 400 452436 406
rect 452384 342 452436 348
rect 448980 196 449032 202
rect 448980 138 449032 144
rect 448256 54 448694 82
rect 448582 -960 448694 54
rect 449778 -960 449890 326
rect 450882 -960 450994 326
rect 451280 332 451332 338
rect 451280 274 451332 280
rect 452078 326 452332 342
rect 452078 -960 452190 326
rect 453274 82 453386 480
rect 453488 128 453540 134
rect 453274 76 453488 82
rect 453274 70 453540 76
rect 453274 54 453528 70
rect 453274 -960 453386 54
rect 454470 -960 454582 480
rect 455340 66 455492 82
rect 455328 60 455492 66
rect 455380 54 455492 60
rect 455328 2 455380 8
rect 455666 -960 455778 480
rect 455880 478 455932 484
rect 456904 480 456932 614
rect 458088 604 458140 610
rect 459190 575 459246 584
rect 459558 640 459614 649
rect 460388 614 460440 620
rect 460664 672 460716 678
rect 462136 672 462188 678
rect 461582 640 461638 649
rect 460664 614 460716 620
rect 459558 575 459614 584
rect 458088 546 458140 552
rect 458100 480 458128 546
rect 459008 536 459060 542
rect 458896 484 459008 490
rect 456524 128 456576 134
rect 456576 76 456688 82
rect 456524 70 456688 76
rect 456536 54 456688 70
rect 456862 -960 456974 480
rect 457904 400 457956 406
rect 457792 348 457904 354
rect 457792 342 457956 348
rect 457792 326 457944 342
rect 458058 -960 458170 480
rect 458896 478 459060 484
rect 459204 480 459232 575
rect 458896 462 459048 478
rect 459162 -960 459274 480
rect 459572 474 459600 575
rect 460092 474 460244 490
rect 460400 480 460428 614
rect 460676 513 460704 614
rect 461196 610 461532 626
rect 461196 604 461544 610
rect 461196 598 461492 604
rect 466368 672 466420 678
rect 463054 640 463110 649
rect 462188 620 462300 626
rect 462136 614 462300 620
rect 462148 598 462300 614
rect 462608 598 462820 626
rect 461582 575 461638 584
rect 461492 546 461544 552
rect 460662 504 460718 513
rect 459560 468 459612 474
rect 460092 468 460256 474
rect 460092 462 460204 468
rect 459560 410 459612 416
rect 460204 410 460256 416
rect 460358 -960 460470 480
rect 461596 480 461624 575
rect 460662 439 460718 448
rect 461554 -960 461666 480
rect 462608 218 462636 598
rect 462792 480 462820 598
rect 465170 640 465226 649
rect 463496 610 463648 626
rect 463496 604 463660 610
rect 463496 598 463608 604
rect 463054 575 463110 584
rect 462424 202 462636 218
rect 462412 196 462636 202
rect 462464 190 462636 196
rect 462412 138 462464 144
rect 462750 -960 462862 480
rect 463068 270 463096 575
rect 463608 546 463660 552
rect 463804 598 464016 626
rect 463804 513 463832 598
rect 463790 504 463846 513
rect 463988 480 464016 598
rect 465170 575 465226 584
rect 465354 640 465410 649
rect 465354 575 465410 584
rect 466182 640 466238 649
rect 466366 640 466368 649
rect 467196 672 467248 678
rect 466420 640 466422 649
rect 466238 598 466316 626
rect 466182 575 466238 584
rect 465184 480 465212 575
rect 463790 439 463846 448
rect 463056 264 463108 270
rect 463056 206 463108 212
rect 463946 -960 464058 480
rect 464896 264 464948 270
rect 464600 212 464896 218
rect 464600 206 464948 212
rect 464600 190 464936 206
rect 465142 -960 465254 480
rect 465368 338 465396 575
rect 466288 480 466316 598
rect 466900 620 467196 626
rect 468300 672 468352 678
rect 466900 614 467248 620
rect 467470 640 467526 649
rect 466900 598 467236 614
rect 466366 575 466422 584
rect 468004 620 468300 626
rect 468004 614 468352 620
rect 468668 672 468720 678
rect 477868 672 477920 678
rect 471058 640 471114 649
rect 468668 614 468720 620
rect 468004 598 468340 614
rect 467470 575 467526 584
rect 467484 480 467512 575
rect 467838 504 467894 513
rect 465356 332 465408 338
rect 465356 274 465408 280
rect 466000 128 466052 134
rect 465704 76 466000 82
rect 465704 70 466052 76
rect 465704 54 466040 70
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468680 480 468708 614
rect 469692 598 469904 626
rect 470304 610 470640 626
rect 470304 604 470652 610
rect 470304 598 470600 604
rect 467838 439 467894 448
rect 467852 202 467880 439
rect 467840 196 467892 202
rect 467840 138 467892 144
rect 468638 -960 468750 480
rect 469108 474 469260 490
rect 469108 468 469272 474
rect 469108 462 469220 468
rect 469220 410 469272 416
rect 469692 354 469720 598
rect 469876 480 469904 598
rect 475106 640 475162 649
rect 471408 610 471744 626
rect 471408 604 471756 610
rect 471408 598 471704 604
rect 471058 575 471114 584
rect 470600 546 470652 552
rect 471072 480 471100 575
rect 471704 546 471756 552
rect 472256 604 472308 610
rect 472256 546 472308 552
rect 473280 598 473492 626
rect 472268 480 472296 546
rect 469600 326 469720 354
rect 469600 66 469628 326
rect 469588 60 469640 66
rect 469588 2 469640 8
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473280 406 473308 598
rect 473464 480 473492 598
rect 474556 604 474608 610
rect 474812 598 475106 626
rect 482928 672 482980 678
rect 477868 614 477920 620
rect 475106 575 475162 584
rect 475752 604 475804 610
rect 474556 546 474608 552
rect 475752 546 475804 552
rect 476948 604 477000 610
rect 476948 546 477000 552
rect 474002 504 474058 513
rect 473268 400 473320 406
rect 472512 338 472848 354
rect 473268 342 473320 348
rect 472512 332 472860 338
rect 472512 326 472808 332
rect 472808 274 472860 280
rect 473422 -960 473534 480
rect 473708 462 474002 490
rect 474568 480 474596 546
rect 475764 480 475792 546
rect 476960 480 476988 546
rect 477408 536 477460 542
rect 477112 484 477408 490
rect 474002 439 474058 448
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 475916 66 476252 82
rect 475916 60 476264 66
rect 475916 54 476212 60
rect 476212 2 476264 8
rect 476918 -960 477030 480
rect 477112 478 477460 484
rect 477112 462 477448 478
rect 477880 218 477908 614
rect 478216 598 478552 626
rect 479320 598 479656 626
rect 480516 598 480852 626
rect 482816 620 482928 626
rect 482816 614 482980 620
rect 483020 672 483072 678
rect 483020 614 483072 620
rect 484032 672 484084 678
rect 486608 672 486660 678
rect 484032 614 484084 620
rect 478114 218 478226 480
rect 478524 270 478552 598
rect 477880 190 478226 218
rect 478512 264 478564 270
rect 478512 206 478564 212
rect 479310 218 479422 480
rect 479628 377 479656 598
rect 479614 368 479670 377
rect 479614 303 479670 312
rect 478114 -960 478226 190
rect 479310 202 479564 218
rect 479310 196 479576 202
rect 479310 190 479524 196
rect 479310 -960 479422 190
rect 479524 138 479576 144
rect 480506 82 480618 480
rect 480824 202 480852 598
rect 481732 604 481784 610
rect 482816 598 482968 614
rect 481732 546 481784 552
rect 481744 480 481772 546
rect 480812 196 480864 202
rect 480812 138 480864 144
rect 480720 128 480772 134
rect 480506 76 480720 82
rect 480506 70 480772 76
rect 481456 128 481508 134
rect 481508 76 481620 82
rect 481456 70 481620 76
rect 480506 54 480760 70
rect 481468 54 481620 70
rect 480506 -960 480618 54
rect 481702 -960 481814 480
rect 482806 354 482918 480
rect 483032 354 483060 614
rect 484044 480 484072 614
rect 485024 610 485176 626
rect 486220 610 486372 626
rect 486436 620 486608 626
rect 487436 672 487488 678
rect 486436 614 486660 620
rect 487324 620 487436 626
rect 487324 614 487488 620
rect 487620 672 487672 678
rect 487620 614 487672 620
rect 488264 672 488316 678
rect 492680 672 492732 678
rect 489918 640 489974 649
rect 488316 620 488428 626
rect 488264 614 488428 620
rect 485024 604 485188 610
rect 485024 598 485136 604
rect 485412 604 485464 610
rect 485136 546 485188 552
rect 485240 564 485412 592
rect 485240 480 485268 564
rect 486220 604 486384 610
rect 486220 598 486332 604
rect 485412 546 485464 552
rect 486332 546 486384 552
rect 486436 598 486648 614
rect 487324 598 487476 614
rect 486436 480 486464 598
rect 487632 480 487660 614
rect 488276 598 488428 614
rect 488644 598 488856 626
rect 488644 513 488672 598
rect 488630 504 488686 513
rect 482806 326 483060 354
rect 483768 338 483920 354
rect 483756 332 483920 338
rect 482806 -960 482918 326
rect 483808 326 483920 332
rect 483756 274 483808 280
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488828 480 488856 598
rect 492310 640 492366 649
rect 490728 610 490972 626
rect 490728 604 490984 610
rect 490728 598 490932 604
rect 489918 575 489974 584
rect 489276 536 489328 542
rect 489274 504 489276 513
rect 489328 504 489330 513
rect 488630 439 488686 448
rect 487804 400 487856 406
rect 487802 368 487804 377
rect 487856 368 487858 377
rect 487802 303 487858 312
rect 488786 -960 488898 480
rect 489932 480 489960 575
rect 490932 546 490984 552
rect 491116 604 491168 610
rect 492310 575 492366 584
rect 492678 640 492680 649
rect 496820 672 496872 678
rect 492732 640 492734 649
rect 495898 640 495954 649
rect 492678 575 492734 584
rect 493336 598 493548 626
rect 491116 546 491168 552
rect 491128 480 491156 546
rect 492324 480 492352 575
rect 492678 504 492734 513
rect 489274 439 489330 448
rect 489624 202 489776 218
rect 489624 196 489788 202
rect 489624 190 489736 196
rect 489736 138 489788 144
rect 489890 -960 490002 480
rect 490286 368 490342 377
rect 490286 303 490342 312
rect 490300 270 490328 303
rect 490288 264 490340 270
rect 490288 206 490340 212
rect 491086 -960 491198 480
rect 492128 264 492180 270
rect 491832 212 492128 218
rect 491832 206 492180 212
rect 491832 190 492168 206
rect 492282 -960 492394 480
rect 492600 462 492678 490
rect 492600 406 492628 462
rect 492678 439 492734 448
rect 492588 400 492640 406
rect 493336 377 493364 598
rect 493520 480 493548 598
rect 494532 598 494744 626
rect 494532 513 494560 598
rect 494518 504 494574 513
rect 492588 342 492640 348
rect 493322 368 493378 377
rect 493322 303 493378 312
rect 493028 66 493364 82
rect 493028 60 493376 66
rect 493028 54 493324 60
rect 493324 2 493376 8
rect 493478 -960 493590 480
rect 494716 480 494744 598
rect 495898 575 495954 584
rect 496818 640 496820 649
rect 498200 672 498252 678
rect 496872 640 496874 649
rect 496818 575 496874 584
rect 496924 598 497136 626
rect 498936 672 498988 678
rect 498200 614 498252 620
rect 498640 620 498936 626
rect 502340 672 502392 678
rect 500590 640 500646 649
rect 498640 614 498988 620
rect 495530 504 495586 513
rect 494518 439 494574 448
rect 494428 400 494480 406
rect 494132 348 494428 354
rect 494132 342 494480 348
rect 494132 326 494468 342
rect 494674 -960 494786 480
rect 495236 474 495388 490
rect 495236 468 495400 474
rect 495236 462 495348 468
rect 495912 480 495940 575
rect 496728 536 496780 542
rect 496432 484 496728 490
rect 495530 439 495586 448
rect 495348 410 495400 416
rect 495544 338 495572 439
rect 495532 332 495584 338
rect 495532 274 495584 280
rect 495870 -960 495982 480
rect 496432 478 496780 484
rect 496432 462 496768 478
rect 496924 354 496952 598
rect 497108 480 497136 598
rect 498212 480 498240 614
rect 498640 598 498976 614
rect 499224 598 499436 626
rect 499026 504 499082 513
rect 496832 326 496952 354
rect 496832 134 496860 326
rect 496820 128 496872 134
rect 496820 70 496872 76
rect 497066 -960 497178 480
rect 497536 338 497872 354
rect 497536 332 497884 338
rect 497536 326 497832 332
rect 497832 274 497884 280
rect 498170 -960 498282 480
rect 499224 490 499252 598
rect 499082 462 499252 490
rect 499408 480 499436 598
rect 502044 620 502340 626
rect 502044 614 502392 620
rect 502984 672 503036 678
rect 505744 672 505796 678
rect 502984 614 503036 620
rect 500590 575 500646 584
rect 501788 604 501840 610
rect 500604 480 500632 575
rect 502044 598 502380 614
rect 501788 546 501840 552
rect 501234 504 501290 513
rect 499026 439 499082 448
rect 499366 -960 499478 480
rect 500132 128 500184 134
rect 499836 76 500132 82
rect 499836 70 500184 76
rect 499836 54 500172 70
rect 500562 -960 500674 480
rect 500940 462 501234 490
rect 501800 480 501828 546
rect 502996 480 503024 614
rect 504008 598 504220 626
rect 505448 620 505744 626
rect 507860 672 507912 678
rect 507734 632 507860 660
rect 505448 614 505796 620
rect 505448 598 505784 614
rect 506216 598 506520 626
rect 507734 612 507762 632
rect 509884 672 509936 678
rect 509698 640 509754 649
rect 507860 614 507912 620
rect 508944 598 509280 626
rect 501234 439 501290 448
rect 501758 -960 501870 480
rect 502708 264 502760 270
rect 502706 232 502708 241
rect 502760 232 502762 241
rect 502706 167 502762 176
rect 502954 -960 503066 480
rect 504008 406 504036 598
rect 504192 480 504220 598
rect 503996 400 504048 406
rect 503996 342 504048 348
rect 503536 264 503588 270
rect 503240 212 503536 218
rect 503240 206 503588 212
rect 503240 190 503576 206
rect 504150 -960 504262 480
rect 504344 474 504680 490
rect 504344 468 504692 474
rect 504344 462 504640 468
rect 504640 410 504692 416
rect 505346 218 505458 480
rect 506216 474 506244 598
rect 506492 480 506520 598
rect 506938 504 506994 513
rect 506204 468 506256 474
rect 506204 410 506256 416
rect 505204 202 505458 218
rect 505192 196 505458 202
rect 505244 190 505458 196
rect 505192 138 505244 144
rect 505346 -960 505458 190
rect 506450 -960 506562 480
rect 506938 439 506940 448
rect 506992 439 506994 448
rect 506940 410 506992 416
rect 507306 232 507362 241
rect 506644 202 506980 218
rect 506644 196 506992 202
rect 506644 190 506940 196
rect 507646 218 507758 480
rect 507362 190 507758 218
rect 507306 167 507362 176
rect 506940 138 506992 144
rect 507646 -960 507758 190
rect 508842 82 508954 480
rect 509252 406 509280 598
rect 510034 660 510062 748
rect 563408 734 563744 762
rect 509936 632 510062 660
rect 510988 672 511040 678
rect 509884 614 509936 620
rect 512460 672 512512 678
rect 511040 620 511152 626
rect 510988 614 511152 620
rect 512460 614 512512 620
rect 514392 672 514444 678
rect 515956 672 516008 678
rect 514444 620 514556 626
rect 514392 614 514556 620
rect 516968 672 517020 678
rect 515956 614 516008 620
rect 516856 620 516968 626
rect 518256 672 518308 678
rect 516856 614 517020 620
rect 517960 620 518256 626
rect 509698 575 509754 584
rect 510252 604 510304 610
rect 509712 474 509740 575
rect 511000 598 511152 614
rect 510252 546 510304 552
rect 511276 564 511488 592
rect 509700 468 509752 474
rect 509700 410 509752 416
rect 509240 400 509292 406
rect 509240 342 509292 348
rect 508608 66 508954 82
rect 508596 60 508954 66
rect 508648 54 508954 60
rect 508596 2 508648 8
rect 508842 -960 508954 54
rect 510038 218 510150 480
rect 510264 218 510292 546
rect 511276 480 511304 564
rect 510038 190 510292 218
rect 510038 -960 510150 190
rect 511234 -960 511346 480
rect 511460 474 511488 564
rect 512472 480 512500 614
rect 513564 604 513616 610
rect 514404 598 514556 614
rect 513564 546 513616 552
rect 514772 564 514984 592
rect 511448 468 511500 474
rect 511448 410 511500 416
rect 512196 202 512348 218
rect 512184 196 512348 202
rect 512236 190 512348 196
rect 512184 138 512236 144
rect 512430 -960 512542 480
rect 513300 474 513452 490
rect 513576 480 513604 546
rect 514772 480 514800 564
rect 513288 468 513452 474
rect 513340 462 513452 468
rect 513288 410 513340 416
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 514956 474 514984 564
rect 515968 480 515996 614
rect 516856 598 517008 614
rect 517150 606 517206 615
rect 517960 614 518308 620
rect 518348 672 518400 678
rect 519452 672 519504 678
rect 518348 614 518400 620
rect 519156 620 519452 626
rect 519156 614 519504 620
rect 520740 672 520792 678
rect 521936 672 521988 678
rect 520740 614 520792 620
rect 521856 620 521936 626
rect 522856 672 522908 678
rect 521856 614 521988 620
rect 522560 620 522856 626
rect 522560 614 522908 620
rect 523500 672 523552 678
rect 530124 672 530176 678
rect 523552 620 523664 626
rect 523500 614 523664 620
rect 517960 598 518296 614
rect 517150 541 517206 550
rect 517164 480 517192 541
rect 518360 480 518388 614
rect 519156 598 519492 614
rect 519544 604 519596 610
rect 519544 546 519596 552
rect 519556 480 519584 546
rect 520752 480 520780 614
rect 521856 598 521976 614
rect 522560 598 522896 614
rect 523040 604 523092 610
rect 521856 480 521884 598
rect 523512 598 523664 614
rect 524768 610 525104 626
rect 524236 604 524288 610
rect 523040 546 523092 552
rect 524768 604 525116 610
rect 524768 598 525064 604
rect 524236 546 524288 552
rect 525064 546 525116 552
rect 525260 598 525472 626
rect 525964 610 526300 626
rect 525964 604 526312 610
rect 525964 598 526260 604
rect 523052 480 523080 546
rect 524248 480 524276 546
rect 514944 468 514996 474
rect 514944 410 514996 416
rect 515588 128 515640 134
rect 515640 76 515752 82
rect 515588 70 515752 76
rect 515600 54 515752 70
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520260 338 520412 354
rect 520260 332 520424 338
rect 520260 326 520372 332
rect 520372 274 520424 280
rect 520710 -960 520822 480
rect 521364 202 521608 218
rect 521364 196 521620 202
rect 521364 190 521568 196
rect 521568 138 521620 144
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525260 406 525288 598
rect 525444 480 525472 598
rect 526260 546 526312 552
rect 526456 598 526668 626
rect 526456 490 526484 598
rect 525248 400 525300 406
rect 525248 342 525300 348
rect 525402 -960 525514 480
rect 526272 462 526484 490
rect 526640 480 526668 598
rect 528848 598 529060 626
rect 531136 672 531188 678
rect 530124 614 530176 620
rect 531134 640 531136 649
rect 531320 672 531372 678
rect 531188 640 531190 649
rect 527560 564 527864 592
rect 526272 66 526300 462
rect 526260 60 526312 66
rect 526260 2 526312 8
rect 526598 -960 526710 480
rect 527560 474 527588 564
rect 527836 480 527864 564
rect 527548 468 527600 474
rect 527548 410 527600 416
rect 527180 400 527232 406
rect 527068 348 527180 354
rect 527068 342 527232 348
rect 527068 326 527220 342
rect 527794 -960 527906 480
rect 528848 270 528876 598
rect 529032 480 529060 598
rect 530136 480 530164 614
rect 531872 672 531924 678
rect 531320 614 531372 620
rect 531576 620 531872 626
rect 548340 672 548392 678
rect 533710 640 533766 649
rect 531576 614 531924 620
rect 531134 575 531190 584
rect 531332 480 531360 614
rect 531576 598 531912 614
rect 532344 598 532556 626
rect 528836 264 528888 270
rect 528836 206 528888 212
rect 528172 66 528508 82
rect 528172 60 528520 66
rect 528172 54 528468 60
rect 528468 2 528520 8
rect 528990 -960 529102 480
rect 529664 264 529716 270
rect 529368 212 529664 218
rect 529368 206 529716 212
rect 529368 190 529704 206
rect 530094 -960 530206 480
rect 530766 232 530822 241
rect 530472 190 530766 218
rect 530766 167 530822 176
rect 531290 -960 531402 480
rect 532344 134 532372 598
rect 532528 480 532556 598
rect 534170 640 534226 649
rect 533876 598 534170 626
rect 533710 575 533766 584
rect 548154 640 548210 649
rect 534980 598 535316 626
rect 536176 598 536512 626
rect 537280 598 537616 626
rect 538476 610 538812 626
rect 538476 604 538824 610
rect 538476 598 538772 604
rect 534170 575 534226 584
rect 533068 536 533120 542
rect 532772 484 533068 490
rect 532332 128 532384 134
rect 532332 70 532384 76
rect 532486 -960 532598 480
rect 532772 478 533120 484
rect 533724 480 533752 575
rect 532772 462 533108 478
rect 533682 -960 533794 480
rect 534540 128 534592 134
rect 534878 82 534990 480
rect 535288 105 535316 598
rect 535828 468 535880 474
rect 535828 410 535880 416
rect 535840 354 535868 410
rect 536074 354 536186 480
rect 536484 474 536512 598
rect 536472 468 536524 474
rect 536472 410 536524 416
rect 537178 354 537290 480
rect 537588 377 537616 598
rect 539580 598 539916 626
rect 542984 610 543136 626
rect 544088 610 544240 626
rect 545132 610 545284 626
rect 538772 546 538824 552
rect 539784 536 539836 542
rect 535840 326 536186 354
rect 536944 338 537290 354
rect 534592 76 534990 82
rect 534540 70 534990 76
rect 534552 54 534990 70
rect 534878 -960 534990 54
rect 535274 96 535330 105
rect 535274 31 535330 40
rect 536074 -960 536186 326
rect 536932 332 537290 338
rect 536984 326 537290 332
rect 536932 274 536984 280
rect 537178 -960 537290 326
rect 537574 368 537630 377
rect 537574 303 537630 312
rect 538374 218 538486 480
rect 538048 202 538486 218
rect 538036 196 538486 202
rect 538088 190 538486 196
rect 538036 138 538088 144
rect 538374 -960 538486 190
rect 539570 354 539682 480
rect 539784 478 539836 484
rect 539796 354 539824 478
rect 539570 326 539824 354
rect 539570 -960 539682 326
rect 539888 202 539916 598
rect 540796 604 540848 610
rect 540796 546 540848 552
rect 541992 604 542044 610
rect 542984 604 543148 610
rect 542984 598 543096 604
rect 541992 546 542044 552
rect 543372 604 543424 610
rect 543096 546 543148 552
rect 543200 564 543372 592
rect 540518 504 540574 513
rect 540574 462 540684 490
rect 540808 480 540836 546
rect 542004 480 542032 546
rect 543200 480 543228 564
rect 544088 604 544252 610
rect 544088 598 544200 604
rect 543372 546 543424 552
rect 544200 546 544252 552
rect 544384 604 544436 610
rect 544384 546 544436 552
rect 545120 604 545284 610
rect 545172 598 545284 604
rect 545488 604 545540 610
rect 545120 546 545172 552
rect 545488 546 545540 552
rect 546512 564 546724 592
rect 544396 480 544424 546
rect 545500 480 545528 546
rect 540518 439 540574 448
rect 539876 196 539928 202
rect 539876 138 539928 144
rect 540766 -960 540878 480
rect 541728 338 541880 354
rect 541716 332 541880 338
rect 541768 326 541880 332
rect 541716 274 541768 280
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546512 270 546540 564
rect 546696 480 546724 564
rect 547892 564 548104 592
rect 548338 640 548340 649
rect 548984 672 549036 678
rect 548392 640 548394 649
rect 548210 598 548288 626
rect 548154 575 548210 584
rect 547892 480 547920 564
rect 546500 264 546552 270
rect 546500 206 546552 212
rect 546388 66 546540 82
rect 546388 60 546552 66
rect 546388 54 546500 60
rect 546500 2 546552 8
rect 546654 -960 546766 480
rect 547696 400 547748 406
rect 547492 348 547696 354
rect 547492 342 547748 348
rect 547492 326 547736 342
rect 547850 -960 547962 480
rect 548076 241 548104 564
rect 548260 241 548288 598
rect 548688 620 548984 626
rect 551100 672 551152 678
rect 548688 614 549036 620
rect 549074 640 549130 649
rect 548688 598 549024 614
rect 548338 575 548394 584
rect 549074 575 549130 584
rect 549258 640 549314 649
rect 550896 620 551100 626
rect 552388 672 552440 678
rect 550896 614 551152 620
rect 552092 620 552388 626
rect 565636 672 565688 678
rect 552092 614 552440 620
rect 559746 640 559802 649
rect 550896 598 551140 614
rect 552092 598 552428 614
rect 549258 575 549314 584
rect 549088 480 549116 575
rect 549272 542 549300 575
rect 550284 564 550496 592
rect 549260 536 549312 542
rect 550088 536 550140 542
rect 548062 232 548118 241
rect 548062 167 548118 176
rect 548246 232 548302 241
rect 548246 167 548302 176
rect 549046 -960 549158 480
rect 549260 478 549312 484
rect 549792 484 550088 490
rect 549792 478 550140 484
rect 550284 480 550312 564
rect 549792 462 550128 478
rect 550242 -960 550354 480
rect 550468 134 550496 564
rect 551296 564 551508 592
rect 551296 241 551324 564
rect 551480 480 551508 564
rect 552492 564 552704 592
rect 551282 232 551338 241
rect 551282 167 551338 176
rect 550456 128 550508 134
rect 550456 70 550508 76
rect 551438 -960 551550 480
rect 552492 354 552520 564
rect 552676 480 552704 564
rect 553504 564 553808 592
rect 552400 326 552520 354
rect 552400 105 552428 326
rect 552386 96 552442 105
rect 552386 31 552442 40
rect 552634 -960 552746 480
rect 553504 474 553532 564
rect 553780 480 553808 564
rect 554792 564 555004 592
rect 554596 536 554648 542
rect 554300 484 554596 490
rect 553492 468 553544 474
rect 553492 410 553544 416
rect 553308 400 553360 406
rect 553196 348 553308 354
rect 553196 342 553360 348
rect 553196 326 553348 342
rect 553738 -960 553850 480
rect 554300 478 554648 484
rect 554300 462 554636 478
rect 554792 377 554820 564
rect 554976 480 555004 564
rect 555988 564 556200 592
rect 555792 536 555844 542
rect 555496 484 555792 490
rect 555988 490 556016 564
rect 554778 368 554834 377
rect 554778 303 554834 312
rect 554934 -960 555046 480
rect 555496 478 555844 484
rect 555496 462 555832 478
rect 555896 462 556016 490
rect 556172 480 556200 564
rect 557184 564 557396 592
rect 555896 338 555924 462
rect 555884 332 555936 338
rect 555884 274 555936 280
rect 556130 -960 556242 480
rect 556600 474 556936 490
rect 556600 468 556948 474
rect 556600 462 556896 468
rect 556896 410 556948 416
rect 557184 202 557212 564
rect 557368 480 557396 564
rect 558380 564 558592 592
rect 559746 575 559802 584
rect 560852 604 560904 610
rect 558380 513 558408 564
rect 558366 504 558422 513
rect 557172 196 557224 202
rect 557172 138 557224 144
rect 557326 -960 557438 480
rect 558564 480 558592 564
rect 559760 480 559788 575
rect 560852 546 560904 552
rect 562048 604 562100 610
rect 562048 546 562100 552
rect 563244 604 563296 610
rect 563244 546 563296 552
rect 564452 598 564664 626
rect 565636 614 565688 620
rect 560864 480 560892 546
rect 562060 480 562088 546
rect 563256 480 563284 546
rect 564452 480 564480 598
rect 558366 439 558422 448
rect 557704 338 558040 354
rect 557704 332 558052 338
rect 557704 326 558000 332
rect 558000 274 558052 280
rect 558522 -960 558634 480
rect 558900 338 559052 354
rect 558900 332 559064 338
rect 558900 326 559012 332
rect 559012 274 559064 280
rect 559718 -960 559830 480
rect 560004 202 560248 218
rect 560004 196 560260 202
rect 560004 190 560208 196
rect 560208 138 560260 144
rect 560822 -960 560934 480
rect 561108 66 561444 82
rect 561108 60 561456 66
rect 561108 54 561404 60
rect 561404 2 561456 8
rect 562018 -960 562130 480
rect 562600 264 562652 270
rect 562304 212 562600 218
rect 562304 206 562652 212
rect 562304 190 562640 206
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 564636 134 564664 598
rect 565648 480 565676 614
rect 566844 480 566872 818
rect 568028 808 568080 814
rect 568028 750 568080 756
rect 568040 480 568068 750
rect 569144 480 569172 886
rect 570328 740 570380 746
rect 570328 682 570380 688
rect 570340 480 570368 682
rect 571352 598 571564 626
rect 571352 490 571380 598
rect 564624 128 564676 134
rect 564624 70 564676 76
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571168 462 571380 490
rect 571536 480 571564 598
rect 572732 480 572760 2858
rect 576308 2848 576360 2854
rect 576308 2790 576360 2796
rect 573916 604 573968 610
rect 573916 546 573968 552
rect 575112 604 575164 610
rect 575112 546 575164 552
rect 573928 480 573956 546
rect 575124 480 575152 546
rect 576320 480 576348 2790
rect 577240 598 577452 626
rect 577240 490 577268 598
rect 571168 406 571196 462
rect 571156 400 571208 406
rect 571156 342 571208 348
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 576872 462 577268 490
rect 577424 480 577452 598
rect 578436 598 578648 626
rect 576872 354 576900 462
rect 576780 338 576900 354
rect 576768 332 576900 338
rect 576820 326 576900 332
rect 576768 274 576820 280
rect 577382 -960 577494 480
rect 578436 354 578464 598
rect 578620 480 578648 598
rect 580828 598 581040 626
rect 578344 326 578464 354
rect 578344 202 578372 326
rect 578332 196 578384 202
rect 578332 138 578384 144
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580828 218 580856 598
rect 581012 480 581040 598
rect 582024 598 582236 626
rect 580736 190 580856 218
rect 580736 66 580764 190
rect 580724 60 580776 66
rect 580724 2 580776 8
rect 580970 -960 581082 480
rect 582024 354 582052 598
rect 582208 480 582236 598
rect 583404 480 583432 2994
rect 581840 326 582052 354
rect 581840 270 581868 326
rect 581828 264 581880 270
rect 581828 206 581880 212
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 18 702072 74 702128
rect 662 700168 718 700224
rect 938 700576 994 700632
rect 1490 684256 1546 684312
rect 1582 632032 1638 632088
rect 938 606056 994 606112
rect 1766 698128 1822 698184
rect 1674 579944 1730 580000
rect 846 553832 902 553888
rect 2226 701392 2282 701448
rect 2042 701256 2098 701312
rect 1950 697856 2006 697912
rect 1858 527856 1914 527912
rect 1766 475632 1822 475688
rect 754 449520 810 449576
rect 1950 423544 2006 423600
rect 662 397432 718 397488
rect 570 254088 626 254144
rect 570 214920 626 214976
rect 570 188808 626 188864
rect 570 162832 626 162888
rect 202 111152 258 111208
rect 110 71848 166 71904
rect 18 19896 74 19952
rect 2134 699760 2190 699816
rect 4250 701800 4306 701856
rect 2502 697584 2558 697640
rect 2962 700440 3018 700496
rect 2686 697720 2742 697776
rect 3146 700304 3202 700360
rect 3054 658144 3110 658200
rect 2962 566888 3018 566944
rect 2778 514800 2834 514856
rect 3606 699896 3662 699952
rect 3422 699080 3478 699136
rect 3330 697992 3386 698048
rect 3238 671200 3294 671256
rect 3146 462576 3202 462632
rect 3330 501744 3386 501800
rect 3238 410488 3294 410544
rect 2686 371320 2742 371376
rect 2594 358400 2650 358456
rect 2502 345344 2558 345400
rect 2410 319232 2466 319288
rect 2318 267144 2374 267200
rect 3330 97552 3386 97608
rect 2226 58520 2282 58576
rect 3790 619112 3846 619168
rect 3698 201864 3754 201920
rect 3606 149776 3662 149832
rect 3514 136720 3570 136776
rect 4066 700032 4122 700088
rect 4434 701528 4490 701584
rect 21454 702480 21510 702536
rect 60646 701936 60702 701992
rect 46018 701664 46074 701720
rect 134430 701120 134486 701176
rect 286690 701120 286746 701176
rect 291474 701120 291530 701176
rect 6642 699352 6698 699408
rect 11610 699352 11666 699408
rect 16394 699352 16450 699408
rect 26146 699352 26202 699408
rect 31206 699352 31262 699408
rect 41050 699352 41106 699408
rect 379518 700576 379574 700632
rect 399022 700440 399078 700496
rect 428462 700304 428518 700360
rect 438628 700168 438684 700224
rect 433430 699488 433486 699544
rect 472714 700032 472770 700088
rect 526718 701800 526774 701856
rect 516966 699896 517022 699952
rect 531686 701528 531742 701584
rect 546498 701392 546554 701448
rect 556250 701256 556306 701312
rect 561126 702072 561182 702128
rect 565174 701936 565230 701992
rect 551282 699760 551338 699816
rect 408958 699352 409014 699408
rect 418710 699352 418766 699408
rect 444286 699352 444342 699408
rect 448150 699352 448206 699408
rect 453118 699352 453174 699408
rect 565082 698264 565138 698320
rect 4066 306176 4122 306232
rect 3974 293120 4030 293176
rect 3882 241032 3938 241088
rect 3790 84632 3846 84688
rect 3422 45464 3478 45520
rect 2134 32408 2190 32464
rect 571982 701664 572038 701720
rect 566646 698944 566702 699000
rect 565266 698672 565322 698728
rect 566462 698536 566518 698592
rect 569222 698400 569278 698456
rect 569406 698808 569462 698864
rect 576122 702480 576178 702536
rect 580170 697176 580226 697232
rect 580170 683848 580226 683904
rect 580170 670656 580226 670712
rect 578974 644000 579030 644056
rect 580170 630808 580226 630864
rect 580170 617480 580226 617536
rect 579802 577632 579858 577688
rect 580170 564340 580172 564360
rect 580172 564340 580224 564360
rect 580224 564340 580226 564360
rect 580170 564304 580226 564340
rect 580170 537784 580226 537840
rect 580170 511264 580226 511320
rect 579618 484608 579674 484664
rect 578882 431568 578938 431624
rect 579618 418240 579674 418296
rect 579802 404912 579858 404968
rect 579802 378392 579858 378448
rect 580170 351872 580226 351928
rect 580170 325216 580226 325272
rect 580170 312024 580226 312080
rect 580170 298696 580226 298752
rect 580170 272176 580226 272232
rect 579618 258848 579674 258904
rect 580170 245556 580172 245576
rect 580172 245556 580224 245576
rect 580224 245556 580226 245576
rect 580170 245520 580226 245556
rect 580170 232328 580226 232384
rect 580170 219000 580226 219056
rect 579894 205672 579950 205728
rect 579986 179152 580042 179208
rect 580170 165824 580226 165880
rect 580446 697992 580502 698048
rect 580814 590960 580870 591016
rect 580722 524456 580778 524512
rect 580630 471416 580686 471472
rect 580538 458088 580594 458144
rect 580446 365064 580502 365120
rect 580354 192480 580410 192536
rect 580262 152632 580318 152688
rect 580170 139340 580172 139360
rect 580172 139340 580224 139360
rect 580224 139340 580226 139360
rect 580170 139304 580226 139340
rect 580170 125976 580226 126032
rect 579802 112784 579858 112840
rect 580170 99456 580226 99512
rect 580170 86128 580226 86184
rect 580170 72936 580226 72992
rect 580170 59608 580226 59664
rect 580170 46280 580226 46336
rect 580170 33108 580226 33144
rect 580170 33088 580172 33108
rect 580172 33088 580224 33108
rect 580224 33088 580226 33108
rect 579986 19760 580042 19816
rect 580170 6568 580226 6624
rect 2042 6432 2098 6488
rect 4066 584 4122 640
rect 7838 584 7894 640
rect 9954 584 10010 640
rect 13266 584 13322 640
rect 18510 448 18566 504
rect 20626 584 20682 640
rect 23478 584 23534 640
rect 21270 448 21326 504
rect 26514 584 26570 640
rect 28722 620 28724 640
rect 28724 620 28776 640
rect 28776 620 28778 640
rect 28722 584 28778 620
rect 27894 448 27950 504
rect 30286 584 30342 640
rect 32402 584 32458 640
rect 33230 584 33286 640
rect 35990 584 36046 640
rect 38474 584 38530 640
rect 52550 584 52606 640
rect 56046 584 56102 640
rect 54206 448 54262 504
rect 57610 584 57666 640
rect 58438 584 58494 640
rect 57426 448 57482 504
rect 59818 584 59874 640
rect 58806 448 58862 504
rect 59450 448 59506 504
rect 62026 584 62082 640
rect 61106 448 61162 504
rect 63498 584 63554 640
rect 142066 584 142122 640
rect 143446 584 143502 640
rect 144734 584 144790 640
rect 145746 584 145802 640
rect 143722 448 143778 504
rect 147126 584 147182 640
rect 148966 584 149022 640
rect 147770 448 147826 504
rect 149334 448 149390 504
rect 150622 584 150678 640
rect 151818 584 151874 640
rect 150254 448 150310 504
rect 164790 584 164846 640
rect 167366 584 167422 640
rect 169482 584 169538 640
rect 168194 312 168250 368
rect 171966 584 172022 640
rect 172978 584 173034 640
rect 170954 312 171010 368
rect 171690 312 171746 368
rect 173898 448 173954 504
rect 175462 584 175518 640
rect 176382 584 176438 640
rect 173990 312 174046 368
rect 175186 312 175242 368
rect 176842 448 176898 504
rect 177486 448 177542 504
rect 179050 584 179106 640
rect 180246 584 180302 640
rect 177670 312 177726 368
rect 178682 312 178738 368
rect 182086 584 182142 640
rect 184938 584 184994 640
rect 191102 584 191158 640
rect 181258 312 181314 368
rect 186594 448 186650 504
rect 189906 448 189962 504
rect 194414 584 194470 640
rect 196714 584 196770 640
rect 195242 176 195298 232
rect 197726 312 197782 368
rect 200302 584 200358 640
rect 201498 584 201554 640
rect 203614 584 203670 640
rect 198922 176 198978 232
rect 198922 40 198978 96
rect 200026 312 200082 368
rect 201314 312 201370 368
rect 201866 448 201922 504
rect 201866 176 201922 232
rect 202418 176 202474 232
rect 202510 40 202566 96
rect 203706 448 203762 504
rect 204810 448 204866 504
rect 207386 584 207442 640
rect 208582 584 208638 640
rect 209318 584 209374 640
rect 204902 312 204958 368
rect 206006 176 206062 232
rect 206926 312 206982 368
rect 208214 448 208270 504
rect 210790 312 210846 368
rect 211986 448 212042 504
rect 213366 584 213422 640
rect 216126 448 216182 504
rect 222474 584 222530 640
rect 217230 312 217286 368
rect 220174 448 220230 504
rect 221738 312 221794 368
rect 223578 448 223634 504
rect 227534 584 227590 640
rect 228730 584 228786 640
rect 230938 584 230994 640
rect 235814 584 235870 640
rect 238850 584 238906 640
rect 244094 584 244150 640
rect 243358 448 243414 504
rect 249062 584 249118 640
rect 248970 448 249026 504
rect 249706 448 249762 504
rect 254674 584 254730 640
rect 255870 584 255926 640
rect 263138 584 263194 640
rect 264150 584 264206 640
rect 267278 584 267334 640
rect 273626 584 273682 640
rect 275834 584 275890 640
rect 275190 448 275246 504
rect 279238 312 279294 368
rect 283102 584 283158 640
rect 282182 448 282238 504
rect 285218 448 285274 504
rect 286598 584 286654 640
rect 287058 584 287114 640
rect 287794 584 287850 640
rect 291566 584 291622 640
rect 293682 584 293738 640
rect 293866 584 293922 640
rect 294878 584 294934 640
rect 292762 448 292818 504
rect 305826 584 305882 640
rect 307022 448 307078 504
rect 313830 584 313886 640
rect 315026 584 315082 640
rect 316590 584 316646 640
rect 317326 584 317382 640
rect 326342 312 326398 368
rect 334254 584 334310 640
rect 335358 448 335414 504
rect 335266 312 335322 368
rect 343362 584 343418 640
rect 336554 312 336610 368
rect 344558 584 344614 640
rect 345754 584 345810 640
rect 345938 584 345994 640
rect 346950 584 347006 640
rect 347778 584 347834 640
rect 350446 584 350502 640
rect 351826 584 351882 640
rect 352838 584 352894 640
rect 364430 584 364486 640
rect 366086 448 366142 504
rect 375286 584 375342 640
rect 376482 584 376538 640
rect 383106 312 383162 368
rect 384210 448 384266 504
rect 385774 196 385830 232
rect 385774 176 385776 196
rect 385776 176 385828 196
rect 385828 176 385830 196
rect 386970 332 387026 368
rect 386970 312 386972 332
rect 386972 312 387024 332
rect 387024 312 387026 332
rect 389822 484 389824 504
rect 389824 484 389876 504
rect 389876 484 389878 504
rect 389822 448 389878 484
rect 391570 176 391626 232
rect 392214 448 392270 504
rect 393778 584 393834 640
rect 401322 584 401378 640
rect 400310 448 400366 504
rect 421102 620 421104 640
rect 421104 620 421156 640
rect 421156 620 421158 640
rect 417146 448 417202 504
rect 421102 584 421158 620
rect 424966 584 425022 640
rect 425518 620 425520 640
rect 425520 620 425572 640
rect 425572 620 425574 640
rect 425518 584 425574 620
rect 426162 584 426218 640
rect 429658 584 429714 640
rect 445574 584 445630 640
rect 459190 584 459246 640
rect 459558 584 459614 640
rect 461582 584 461638 640
rect 460662 448 460718 504
rect 463054 584 463110 640
rect 463790 448 463846 504
rect 465170 584 465226 640
rect 465354 584 465410 640
rect 466182 584 466238 640
rect 466366 620 466368 640
rect 466368 620 466420 640
rect 466420 620 466422 640
rect 466366 584 466422 620
rect 467470 584 467526 640
rect 467838 448 467894 504
rect 471058 584 471114 640
rect 475106 584 475162 640
rect 474002 448 474058 504
rect 479614 312 479670 368
rect 488630 448 488686 504
rect 489918 584 489974 640
rect 489274 484 489276 504
rect 489276 484 489328 504
rect 489328 484 489330 504
rect 487802 348 487804 368
rect 487804 348 487856 368
rect 487856 348 487858 368
rect 487802 312 487858 348
rect 489274 448 489330 484
rect 492310 584 492366 640
rect 492678 620 492680 640
rect 492680 620 492732 640
rect 492732 620 492734 640
rect 492678 584 492734 620
rect 490286 312 490342 368
rect 492678 448 492734 504
rect 493322 312 493378 368
rect 494518 448 494574 504
rect 495898 584 495954 640
rect 496818 620 496820 640
rect 496820 620 496872 640
rect 496872 620 496874 640
rect 496818 584 496874 620
rect 495530 448 495586 504
rect 499026 448 499082 504
rect 500590 584 500646 640
rect 501234 448 501290 504
rect 502706 212 502708 232
rect 502708 212 502760 232
rect 502760 212 502762 232
rect 502706 176 502762 212
rect 506938 468 506994 504
rect 506938 448 506940 468
rect 506940 448 506992 468
rect 506992 448 506994 468
rect 507306 176 507362 232
rect 509698 584 509754 640
rect 517150 550 517206 606
rect 531134 620 531136 640
rect 531136 620 531188 640
rect 531188 620 531190 640
rect 531134 584 531190 620
rect 530766 176 530822 232
rect 533710 584 533766 640
rect 534170 584 534226 640
rect 535274 40 535330 96
rect 537574 312 537630 368
rect 540518 448 540574 504
rect 548154 584 548210 640
rect 548338 620 548340 640
rect 548340 620 548392 640
rect 548392 620 548394 640
rect 548338 584 548394 620
rect 549074 584 549130 640
rect 549258 584 549314 640
rect 548062 176 548118 232
rect 548246 176 548302 232
rect 551282 176 551338 232
rect 552386 40 552442 96
rect 554778 312 554834 368
rect 559746 584 559802 640
rect 558366 448 558422 504
<< metal3 >>
rect 21449 702538 21515 702541
rect 576117 702538 576183 702541
rect 21449 702536 576183 702538
rect 21449 702480 21454 702536
rect 21510 702480 576122 702536
rect 576178 702480 576183 702536
rect 21449 702478 576183 702480
rect 21449 702475 21515 702478
rect 576117 702475 576183 702478
rect 13 702130 79 702133
rect 561121 702130 561187 702133
rect 13 702128 561187 702130
rect 13 702072 18 702128
rect 74 702072 561126 702128
rect 561182 702072 561187 702128
rect 13 702070 561187 702072
rect 13 702067 79 702070
rect 561121 702067 561187 702070
rect 60641 701994 60707 701997
rect 565169 701994 565235 701997
rect 60641 701992 565235 701994
rect 60641 701936 60646 701992
rect 60702 701936 565174 701992
rect 565230 701936 565235 701992
rect 60641 701934 565235 701936
rect 60641 701931 60707 701934
rect 565169 701931 565235 701934
rect 4245 701858 4311 701861
rect 526713 701858 526779 701861
rect 4245 701856 526779 701858
rect 4245 701800 4250 701856
rect 4306 701800 526718 701856
rect 526774 701800 526779 701856
rect 4245 701798 526779 701800
rect 4245 701795 4311 701798
rect 526713 701795 526779 701798
rect 46013 701722 46079 701725
rect 571977 701722 572043 701725
rect 46013 701720 572043 701722
rect 46013 701664 46018 701720
rect 46074 701664 571982 701720
rect 572038 701664 572043 701720
rect 46013 701662 572043 701664
rect 46013 701659 46079 701662
rect 571977 701659 572043 701662
rect 4429 701586 4495 701589
rect 531681 701586 531747 701589
rect 4429 701584 531747 701586
rect 4429 701528 4434 701584
rect 4490 701528 531686 701584
rect 531742 701528 531747 701584
rect 4429 701526 531747 701528
rect 4429 701523 4495 701526
rect 531681 701523 531747 701526
rect 2221 701450 2287 701453
rect 546493 701450 546559 701453
rect 2221 701448 546559 701450
rect 2221 701392 2226 701448
rect 2282 701392 546498 701448
rect 546554 701392 546559 701448
rect 2221 701390 546559 701392
rect 2221 701387 2287 701390
rect 546493 701387 546559 701390
rect 2037 701314 2103 701317
rect 556245 701314 556311 701317
rect 2037 701312 556311 701314
rect 2037 701256 2042 701312
rect 2098 701256 556250 701312
rect 556306 701256 556311 701312
rect 2037 701254 556311 701256
rect 2037 701251 2103 701254
rect 556245 701251 556311 701254
rect 134425 701178 134491 701181
rect 164182 701178 164188 701180
rect 134425 701176 164188 701178
rect 134425 701120 134430 701176
rect 134486 701120 164188 701176
rect 134425 701118 164188 701120
rect 134425 701115 134491 701118
rect 164182 701116 164188 701118
rect 164252 701116 164258 701180
rect 286685 701178 286751 701181
rect 291469 701178 291535 701181
rect 286685 701176 291535 701178
rect 286685 701120 286690 701176
rect 286746 701120 291474 701176
rect 291530 701120 291535 701176
rect 286685 701118 291535 701120
rect 286685 701115 286751 701118
rect 291469 701115 291535 701118
rect 933 700634 999 700637
rect 379513 700634 379579 700637
rect 933 700632 379579 700634
rect 933 700576 938 700632
rect 994 700576 379518 700632
rect 379574 700576 379579 700632
rect 933 700574 379579 700576
rect 933 700571 999 700574
rect 379513 700571 379579 700574
rect 2957 700498 3023 700501
rect 399017 700498 399083 700501
rect 2957 700496 399083 700498
rect 2957 700440 2962 700496
rect 3018 700440 399022 700496
rect 399078 700440 399083 700496
rect 2957 700438 399083 700440
rect 2957 700435 3023 700438
rect 399017 700435 399083 700438
rect 3141 700362 3207 700365
rect 428457 700362 428523 700365
rect 3141 700360 428523 700362
rect 3141 700304 3146 700360
rect 3202 700304 428462 700360
rect 428518 700304 428523 700360
rect 3141 700302 428523 700304
rect 3141 700299 3207 700302
rect 428457 700299 428523 700302
rect 657 700226 723 700229
rect 438623 700226 438689 700229
rect 657 700224 438689 700226
rect 657 700168 662 700224
rect 718 700168 438628 700224
rect 438684 700168 438689 700224
rect 657 700166 438689 700168
rect 657 700163 723 700166
rect 438623 700163 438689 700166
rect 4061 700090 4127 700093
rect 472709 700090 472775 700093
rect 4061 700088 472775 700090
rect 4061 700032 4066 700088
rect 4122 700032 472714 700088
rect 472770 700032 472775 700088
rect 4061 700030 472775 700032
rect 4061 700027 4127 700030
rect 472709 700027 472775 700030
rect 3601 699954 3667 699957
rect 516961 699954 517027 699957
rect 3601 699952 517027 699954
rect 3601 699896 3606 699952
rect 3662 699896 516966 699952
rect 517022 699896 517027 699952
rect 3601 699894 517027 699896
rect 3601 699891 3667 699894
rect 516961 699891 517027 699894
rect 2129 699818 2195 699821
rect 551277 699818 551343 699821
rect 2129 699816 551343 699818
rect 2129 699760 2134 699816
rect 2190 699760 551282 699816
rect 551338 699760 551343 699816
rect 2129 699758 551343 699760
rect 2129 699755 2195 699758
rect 551277 699755 551343 699758
rect 433425 699548 433491 699549
rect 433374 699546 433380 699548
rect 433334 699486 433380 699546
rect 433444 699544 433491 699548
rect 433486 699488 433491 699544
rect 433374 699484 433380 699486
rect 433444 699484 433491 699488
rect 433425 699483 433491 699484
rect 6637 699410 6703 699413
rect 11462 699410 11468 699412
rect 6637 699408 11468 699410
rect 6637 699352 6642 699408
rect 6698 699352 11468 699408
rect 6637 699350 11468 699352
rect 6637 699347 6703 699350
rect 11462 699348 11468 699350
rect 11532 699348 11538 699412
rect 11605 699410 11671 699413
rect 13854 699410 13860 699412
rect 11605 699408 13860 699410
rect 11605 699352 11610 699408
rect 11666 699352 13860 699408
rect 11605 699350 13860 699352
rect 11605 699347 11671 699350
rect 13854 699348 13860 699350
rect 13924 699348 13930 699412
rect 16389 699410 16455 699413
rect 21398 699410 21404 699412
rect 16389 699408 21404 699410
rect 16389 699352 16394 699408
rect 16450 699352 21404 699408
rect 16389 699350 21404 699352
rect 16389 699347 16455 699350
rect 21398 699348 21404 699350
rect 21468 699348 21474 699412
rect 26141 699410 26207 699413
rect 30966 699410 30972 699412
rect 26141 699408 30972 699410
rect 26141 699352 26146 699408
rect 26202 699352 30972 699408
rect 26141 699350 30972 699352
rect 26141 699347 26207 699350
rect 30966 699348 30972 699350
rect 31036 699348 31042 699412
rect 31201 699410 31267 699413
rect 33358 699410 33364 699412
rect 31201 699408 33364 699410
rect 31201 699352 31206 699408
rect 31262 699352 33364 699408
rect 31201 699350 33364 699352
rect 31201 699347 31267 699350
rect 33358 699348 33364 699350
rect 33428 699348 33434 699412
rect 41045 699410 41111 699413
rect 408953 699412 409019 699413
rect 418705 699412 418771 699413
rect 43110 699410 43116 699412
rect 41045 699408 43116 699410
rect 41045 699352 41050 699408
rect 41106 699352 43116 699408
rect 41045 699350 43116 699352
rect 41045 699347 41111 699350
rect 43110 699348 43116 699350
rect 43180 699348 43186 699412
rect 408902 699410 408908 699412
rect 408862 699350 408908 699410
rect 408972 699408 409019 699412
rect 418654 699410 418660 699412
rect 409014 699352 409019 699408
rect 408902 699348 408908 699350
rect 408972 699348 409019 699352
rect 418614 699350 418660 699410
rect 418724 699408 418771 699412
rect 444281 699410 444347 699413
rect 448145 699412 448211 699413
rect 453113 699412 453179 699413
rect 448094 699410 448100 699412
rect 418766 699352 418771 699408
rect 418654 699348 418660 699350
rect 418724 699348 418771 699352
rect 408953 699347 409019 699348
rect 418705 699347 418771 699348
rect 431910 699408 444347 699410
rect 431910 699352 444286 699408
rect 444342 699352 444347 699408
rect 431910 699350 444347 699352
rect 448054 699350 448100 699410
rect 448164 699408 448211 699412
rect 453062 699410 453068 699412
rect 448206 699352 448211 699408
rect 164182 699212 164188 699276
rect 164252 699274 164258 699276
rect 409086 699274 409092 699276
rect 164252 699214 409092 699274
rect 164252 699212 164258 699214
rect 409086 699212 409092 699214
rect 409156 699212 409162 699276
rect 3417 699138 3483 699141
rect 431910 699138 431970 699350
rect 444281 699347 444347 699350
rect 448094 699348 448100 699350
rect 448164 699348 448211 699352
rect 453022 699350 453068 699410
rect 453132 699408 453179 699412
rect 453174 699352 453179 699408
rect 453062 699348 453068 699350
rect 453132 699348 453179 699352
rect 448145 699347 448211 699348
rect 453113 699347 453179 699348
rect 3417 699136 431970 699138
rect 3417 699080 3422 699136
rect 3478 699080 431970 699136
rect 3417 699078 431970 699080
rect 3417 699075 3483 699078
rect 43110 698940 43116 699004
rect 43180 699002 43186 699004
rect 566641 699002 566707 699005
rect 43180 699000 566707 699002
rect 43180 698944 566646 699000
rect 566702 698944 566707 699000
rect 43180 698942 566707 698944
rect 43180 698940 43186 698942
rect 566641 698939 566707 698942
rect 33358 698804 33364 698868
rect 33428 698866 33434 698868
rect 569401 698866 569467 698869
rect 33428 698864 569467 698866
rect 33428 698808 569406 698864
rect 569462 698808 569467 698864
rect 33428 698806 569467 698808
rect 33428 698804 33434 698806
rect 569401 698803 569467 698806
rect 30966 698668 30972 698732
rect 31036 698730 31042 698732
rect 565261 698730 565327 698733
rect 31036 698728 565327 698730
rect 31036 698672 565266 698728
rect 565322 698672 565327 698728
rect 31036 698670 565327 698672
rect 31036 698668 31042 698670
rect 565261 698667 565327 698670
rect 21398 698532 21404 698596
rect 21468 698594 21474 698596
rect 566457 698594 566523 698597
rect 21468 698592 566523 698594
rect 21468 698536 566462 698592
rect 566518 698536 566523 698592
rect 21468 698534 566523 698536
rect 21468 698532 21474 698534
rect 566457 698531 566523 698534
rect 13854 698396 13860 698460
rect 13924 698458 13930 698460
rect 569217 698458 569283 698461
rect 13924 698456 569283 698458
rect 13924 698400 569222 698456
rect 569278 698400 569283 698456
rect 13924 698398 569283 698400
rect 13924 698396 13930 698398
rect 569217 698395 569283 698398
rect 11462 698260 11468 698324
rect 11532 698322 11538 698324
rect 565077 698322 565143 698325
rect 11532 698320 565143 698322
rect 11532 698264 565082 698320
rect 565138 698264 565143 698320
rect 11532 698262 565143 698264
rect 11532 698260 11538 698262
rect 565077 698259 565143 698262
rect 1761 698186 1827 698189
rect 418654 698186 418660 698188
rect 1761 698184 418660 698186
rect 1761 698128 1766 698184
rect 1822 698128 418660 698184
rect 1761 698126 418660 698128
rect 1761 698123 1827 698126
rect 418654 698124 418660 698126
rect 418724 698124 418730 698188
rect 3325 698050 3391 698053
rect 408902 698050 408908 698052
rect 3325 698048 408908 698050
rect 3325 697992 3330 698048
rect 3386 697992 408908 698048
rect 3325 697990 408908 697992
rect 3325 697987 3391 697990
rect 408902 697988 408908 697990
rect 408972 697988 408978 698052
rect 409086 697988 409092 698052
rect 409156 698050 409162 698052
rect 580441 698050 580507 698053
rect 409156 698048 580507 698050
rect 409156 697992 580446 698048
rect 580502 697992 580507 698048
rect 409156 697990 580507 697992
rect 409156 697988 409162 697990
rect 580441 697987 580507 697990
rect 1945 697914 2011 697917
rect 433374 697914 433380 697916
rect 1945 697912 433380 697914
rect 1945 697856 1950 697912
rect 2006 697856 433380 697912
rect 1945 697854 433380 697856
rect 1945 697851 2011 697854
rect 433374 697852 433380 697854
rect 433444 697852 433450 697916
rect 2681 697778 2747 697781
rect 448094 697778 448100 697780
rect 2681 697776 448100 697778
rect 2681 697720 2686 697776
rect 2742 697720 448100 697776
rect 2681 697718 448100 697720
rect 2681 697715 2747 697718
rect 448094 697716 448100 697718
rect 448164 697716 448170 697780
rect 2497 697642 2563 697645
rect 453062 697642 453068 697644
rect 2497 697640 453068 697642
rect 2497 697584 2502 697640
rect 2558 697584 453068 697640
rect 2497 697582 453068 697584
rect 2497 697579 2563 697582
rect 453062 697580 453068 697582
rect 453132 697580 453138 697644
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 1485 684314 1551 684317
rect -960 684312 1551 684314
rect -960 684256 1490 684312
rect 1546 684256 1551 684312
rect -960 684254 1551 684256
rect -960 684164 480 684254
rect 1485 684251 1551 684254
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3233 671258 3299 671261
rect -960 671256 3299 671258
rect -960 671200 3238 671256
rect 3294 671200 3299 671256
rect -960 671198 3299 671200
rect -960 671108 480 671198
rect 3233 671195 3299 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3049 658202 3115 658205
rect -960 658200 3115 658202
rect -960 658144 3054 658200
rect 3110 658144 3115 658200
rect -960 658142 3115 658144
rect -960 658052 480 658142
rect 3049 658139 3115 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 578969 644058 579035 644061
rect 583520 644058 584960 644148
rect 578969 644056 584960 644058
rect 578969 644000 578974 644056
rect 579030 644000 584960 644056
rect 578969 643998 584960 644000
rect 578969 643995 579035 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 1577 632090 1643 632093
rect -960 632088 1643 632090
rect -960 632032 1582 632088
rect 1638 632032 1643 632088
rect -960 632030 1643 632032
rect -960 631940 480 632030
rect 1577 632027 1643 632030
rect 580165 630866 580231 630869
rect 583520 630866 584960 630956
rect 580165 630864 584960 630866
rect 580165 630808 580170 630864
rect 580226 630808 584960 630864
rect 580165 630806 584960 630808
rect 580165 630803 580231 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3785 619170 3851 619173
rect -960 619168 3851 619170
rect -960 619112 3790 619168
rect 3846 619112 3851 619168
rect -960 619110 3851 619112
rect -960 619020 480 619110
rect 3785 619107 3851 619110
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 933 606114 999 606117
rect -960 606112 999 606114
rect -960 606056 938 606112
rect 994 606056 999 606112
rect -960 606054 999 606056
rect -960 605964 480 606054
rect 933 606051 999 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 580809 591018 580875 591021
rect 583520 591018 584960 591108
rect 580809 591016 584960 591018
rect 580809 590960 580814 591016
rect 580870 590960 584960 591016
rect 580809 590958 584960 590960
rect 580809 590955 580875 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 1669 580002 1735 580005
rect -960 580000 1735 580002
rect -960 579944 1674 580000
rect 1730 579944 1735 580000
rect -960 579942 1735 579944
rect -960 579852 480 579942
rect 1669 579939 1735 579942
rect 579797 577690 579863 577693
rect 583520 577690 584960 577780
rect 579797 577688 584960 577690
rect 579797 577632 579802 577688
rect 579858 577632 584960 577688
rect 579797 577630 584960 577632
rect 579797 577627 579863 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 2957 566946 3023 566949
rect -960 566944 3023 566946
rect -960 566888 2962 566944
rect 3018 566888 3023 566944
rect -960 566886 3023 566888
rect -960 566796 480 566886
rect 2957 566883 3023 566886
rect 580165 564362 580231 564365
rect 583520 564362 584960 564452
rect 580165 564360 584960 564362
rect 580165 564304 580170 564360
rect 580226 564304 584960 564360
rect 580165 564302 584960 564304
rect 580165 564299 580231 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 841 553890 907 553893
rect -960 553888 907 553890
rect -960 553832 846 553888
rect 902 553832 907 553888
rect -960 553830 907 553832
rect -960 553740 480 553830
rect 841 553827 907 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 580165 537842 580231 537845
rect 583520 537842 584960 537932
rect 580165 537840 584960 537842
rect 580165 537784 580170 537840
rect 580226 537784 584960 537840
rect 580165 537782 584960 537784
rect 580165 537779 580231 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 1853 527914 1919 527917
rect -960 527912 1919 527914
rect -960 527856 1858 527912
rect 1914 527856 1919 527912
rect -960 527854 1919 527856
rect -960 527764 480 527854
rect 1853 527851 1919 527854
rect 580717 524514 580783 524517
rect 583520 524514 584960 524604
rect 580717 524512 584960 524514
rect 580717 524456 580722 524512
rect 580778 524456 584960 524512
rect 580717 524454 584960 524456
rect 580717 524451 580783 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 2773 514858 2839 514861
rect -960 514856 2839 514858
rect -960 514800 2778 514856
rect 2834 514800 2839 514856
rect -960 514798 2839 514800
rect -960 514708 480 514798
rect 2773 514795 2839 514798
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 3325 501802 3391 501805
rect -960 501800 3391 501802
rect -960 501744 3330 501800
rect 3386 501744 3391 501800
rect -960 501742 3391 501744
rect -960 501652 480 501742
rect 3325 501739 3391 501742
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 579613 484666 579679 484669
rect 583520 484666 584960 484756
rect 579613 484664 584960 484666
rect 579613 484608 579618 484664
rect 579674 484608 584960 484664
rect 579613 484606 584960 484608
rect 579613 484603 579679 484606
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect 1761 475690 1827 475693
rect -960 475688 1827 475690
rect -960 475632 1766 475688
rect 1822 475632 1827 475688
rect -960 475630 1827 475632
rect -960 475540 480 475630
rect 1761 475627 1827 475630
rect 580625 471474 580691 471477
rect 583520 471474 584960 471564
rect 580625 471472 584960 471474
rect 580625 471416 580630 471472
rect 580686 471416 584960 471472
rect 580625 471414 584960 471416
rect 580625 471411 580691 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 3141 462634 3207 462637
rect -960 462632 3207 462634
rect -960 462576 3146 462632
rect 3202 462576 3207 462632
rect -960 462574 3207 462576
rect -960 462484 480 462574
rect 3141 462571 3207 462574
rect 580533 458146 580599 458149
rect 583520 458146 584960 458236
rect 580533 458144 584960 458146
rect 580533 458088 580538 458144
rect 580594 458088 584960 458144
rect 580533 458086 584960 458088
rect 580533 458083 580599 458086
rect 583520 457996 584960 458086
rect -960 449578 480 449668
rect 749 449578 815 449581
rect -960 449576 815 449578
rect -960 449520 754 449576
rect 810 449520 815 449576
rect -960 449518 815 449520
rect -960 449428 480 449518
rect 749 449515 815 449518
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 578877 431626 578943 431629
rect 583520 431626 584960 431716
rect 578877 431624 584960 431626
rect 578877 431568 578882 431624
rect 578938 431568 584960 431624
rect 578877 431566 584960 431568
rect 578877 431563 578943 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 1945 423602 2011 423605
rect -960 423600 2011 423602
rect -960 423544 1950 423600
rect 2006 423544 2011 423600
rect -960 423542 2011 423544
rect -960 423452 480 423542
rect 1945 423539 2011 423542
rect 579613 418298 579679 418301
rect 583520 418298 584960 418388
rect 579613 418296 584960 418298
rect 579613 418240 579618 418296
rect 579674 418240 584960 418296
rect 579613 418238 584960 418240
rect 579613 418235 579679 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 3233 410546 3299 410549
rect -960 410544 3299 410546
rect -960 410488 3238 410544
rect 3294 410488 3299 410544
rect -960 410486 3299 410488
rect -960 410396 480 410486
rect 3233 410483 3299 410486
rect 579797 404970 579863 404973
rect 583520 404970 584960 405060
rect 579797 404968 584960 404970
rect 579797 404912 579802 404968
rect 579858 404912 584960 404968
rect 579797 404910 584960 404912
rect 579797 404907 579863 404910
rect 583520 404820 584960 404910
rect -960 397490 480 397580
rect 657 397490 723 397493
rect -960 397488 723 397490
rect -960 397432 662 397488
rect 718 397432 723 397488
rect -960 397430 723 397432
rect -960 397340 480 397430
rect 657 397427 723 397430
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 579797 378450 579863 378453
rect 583520 378450 584960 378540
rect 579797 378448 584960 378450
rect 579797 378392 579802 378448
rect 579858 378392 584960 378448
rect 579797 378390 584960 378392
rect 579797 378387 579863 378390
rect 583520 378300 584960 378390
rect -960 371378 480 371468
rect 2681 371378 2747 371381
rect -960 371376 2747 371378
rect -960 371320 2686 371376
rect 2742 371320 2747 371376
rect -960 371318 2747 371320
rect -960 371228 480 371318
rect 2681 371315 2747 371318
rect 580441 365122 580507 365125
rect 583520 365122 584960 365212
rect 580441 365120 584960 365122
rect 580441 365064 580446 365120
rect 580502 365064 584960 365120
rect 580441 365062 584960 365064
rect 580441 365059 580507 365062
rect 583520 364972 584960 365062
rect -960 358458 480 358548
rect 2589 358458 2655 358461
rect -960 358456 2655 358458
rect -960 358400 2594 358456
rect 2650 358400 2655 358456
rect -960 358398 2655 358400
rect -960 358308 480 358398
rect 2589 358395 2655 358398
rect 580165 351930 580231 351933
rect 583520 351930 584960 352020
rect 580165 351928 584960 351930
rect 580165 351872 580170 351928
rect 580226 351872 584960 351928
rect 580165 351870 584960 351872
rect 580165 351867 580231 351870
rect 583520 351780 584960 351870
rect -960 345402 480 345492
rect 2497 345402 2563 345405
rect -960 345400 2563 345402
rect -960 345344 2502 345400
rect 2558 345344 2563 345400
rect -960 345342 2563 345344
rect -960 345252 480 345342
rect 2497 345339 2563 345342
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 580165 325274 580231 325277
rect 583520 325274 584960 325364
rect 580165 325272 584960 325274
rect 580165 325216 580170 325272
rect 580226 325216 584960 325272
rect 580165 325214 584960 325216
rect 580165 325211 580231 325214
rect 583520 325124 584960 325214
rect -960 319290 480 319380
rect 2405 319290 2471 319293
rect -960 319288 2471 319290
rect -960 319232 2410 319288
rect 2466 319232 2471 319288
rect -960 319230 2471 319232
rect -960 319140 480 319230
rect 2405 319227 2471 319230
rect 580165 312082 580231 312085
rect 583520 312082 584960 312172
rect 580165 312080 584960 312082
rect 580165 312024 580170 312080
rect 580226 312024 584960 312080
rect 580165 312022 584960 312024
rect 580165 312019 580231 312022
rect 583520 311932 584960 312022
rect -960 306234 480 306324
rect 4061 306234 4127 306237
rect -960 306232 4127 306234
rect -960 306176 4066 306232
rect 4122 306176 4127 306232
rect -960 306174 4127 306176
rect -960 306084 480 306174
rect 4061 306171 4127 306174
rect 580165 298754 580231 298757
rect 583520 298754 584960 298844
rect 580165 298752 584960 298754
rect 580165 298696 580170 298752
rect 580226 298696 584960 298752
rect 580165 298694 584960 298696
rect 580165 298691 580231 298694
rect 583520 298604 584960 298694
rect -960 293178 480 293268
rect 3969 293178 4035 293181
rect -960 293176 4035 293178
rect -960 293120 3974 293176
rect 4030 293120 4035 293176
rect -960 293118 4035 293120
rect -960 293028 480 293118
rect 3969 293115 4035 293118
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 580165 272234 580231 272237
rect 583520 272234 584960 272324
rect 580165 272232 584960 272234
rect 580165 272176 580170 272232
rect 580226 272176 584960 272232
rect 580165 272174 584960 272176
rect 580165 272171 580231 272174
rect 583520 272084 584960 272174
rect -960 267202 480 267292
rect 2313 267202 2379 267205
rect -960 267200 2379 267202
rect -960 267144 2318 267200
rect 2374 267144 2379 267200
rect -960 267142 2379 267144
rect -960 267052 480 267142
rect 2313 267139 2379 267142
rect 579613 258906 579679 258909
rect 583520 258906 584960 258996
rect 579613 258904 584960 258906
rect 579613 258848 579618 258904
rect 579674 258848 584960 258904
rect 579613 258846 584960 258848
rect 579613 258843 579679 258846
rect 583520 258756 584960 258846
rect -960 254146 480 254236
rect 565 254146 631 254149
rect -960 254144 631 254146
rect -960 254088 570 254144
rect 626 254088 631 254144
rect -960 254086 631 254088
rect -960 253996 480 254086
rect 565 254083 631 254086
rect 580165 245578 580231 245581
rect 583520 245578 584960 245668
rect 580165 245576 584960 245578
rect 580165 245520 580170 245576
rect 580226 245520 584960 245576
rect 580165 245518 584960 245520
rect 580165 245515 580231 245518
rect 583520 245428 584960 245518
rect -960 241090 480 241180
rect 3877 241090 3943 241093
rect -960 241088 3943 241090
rect -960 241032 3882 241088
rect 3938 241032 3943 241088
rect -960 241030 3943 241032
rect -960 240940 480 241030
rect 3877 241027 3943 241030
rect 580165 232386 580231 232389
rect 583520 232386 584960 232476
rect 580165 232384 584960 232386
rect 580165 232328 580170 232384
rect 580226 232328 584960 232384
rect 580165 232326 584960 232328
rect 580165 232323 580231 232326
rect 583520 232236 584960 232326
rect -960 227884 480 228124
rect 580165 219058 580231 219061
rect 583520 219058 584960 219148
rect 580165 219056 584960 219058
rect 580165 219000 580170 219056
rect 580226 219000 584960 219056
rect 580165 218998 584960 219000
rect 580165 218995 580231 218998
rect 583520 218908 584960 218998
rect -960 214978 480 215068
rect 565 214978 631 214981
rect -960 214976 631 214978
rect -960 214920 570 214976
rect 626 214920 631 214976
rect -960 214918 631 214920
rect -960 214828 480 214918
rect 565 214915 631 214918
rect 579889 205730 579955 205733
rect 583520 205730 584960 205820
rect 579889 205728 584960 205730
rect 579889 205672 579894 205728
rect 579950 205672 584960 205728
rect 579889 205670 584960 205672
rect 579889 205667 579955 205670
rect 583520 205580 584960 205670
rect -960 201922 480 202012
rect 3693 201922 3759 201925
rect -960 201920 3759 201922
rect -960 201864 3698 201920
rect 3754 201864 3759 201920
rect -960 201862 3759 201864
rect -960 201772 480 201862
rect 3693 201859 3759 201862
rect 580349 192538 580415 192541
rect 583520 192538 584960 192628
rect 580349 192536 584960 192538
rect 580349 192480 580354 192536
rect 580410 192480 584960 192536
rect 580349 192478 584960 192480
rect 580349 192475 580415 192478
rect 583520 192388 584960 192478
rect -960 188866 480 188956
rect 565 188866 631 188869
rect -960 188864 631 188866
rect -960 188808 570 188864
rect 626 188808 631 188864
rect -960 188806 631 188808
rect -960 188716 480 188806
rect 565 188803 631 188806
rect 579981 179210 580047 179213
rect 583520 179210 584960 179300
rect 579981 179208 584960 179210
rect 579981 179152 579986 179208
rect 580042 179152 584960 179208
rect 579981 179150 584960 179152
rect 579981 179147 580047 179150
rect 583520 179060 584960 179150
rect -960 175796 480 176036
rect 580165 165882 580231 165885
rect 583520 165882 584960 165972
rect 580165 165880 584960 165882
rect 580165 165824 580170 165880
rect 580226 165824 584960 165880
rect 580165 165822 584960 165824
rect 580165 165819 580231 165822
rect 583520 165732 584960 165822
rect -960 162890 480 162980
rect 565 162890 631 162893
rect -960 162888 631 162890
rect -960 162832 570 162888
rect 626 162832 631 162888
rect -960 162830 631 162832
rect -960 162740 480 162830
rect 565 162827 631 162830
rect 580257 152690 580323 152693
rect 583520 152690 584960 152780
rect 580257 152688 584960 152690
rect 580257 152632 580262 152688
rect 580318 152632 584960 152688
rect 580257 152630 584960 152632
rect 580257 152627 580323 152630
rect 583520 152540 584960 152630
rect -960 149834 480 149924
rect 3601 149834 3667 149837
rect -960 149832 3667 149834
rect -960 149776 3606 149832
rect 3662 149776 3667 149832
rect -960 149774 3667 149776
rect -960 149684 480 149774
rect 3601 149771 3667 149774
rect 580165 139362 580231 139365
rect 583520 139362 584960 139452
rect 580165 139360 584960 139362
rect 580165 139304 580170 139360
rect 580226 139304 584960 139360
rect 580165 139302 584960 139304
rect 580165 139299 580231 139302
rect 583520 139212 584960 139302
rect -960 136778 480 136868
rect 3509 136778 3575 136781
rect -960 136776 3575 136778
rect -960 136720 3514 136776
rect 3570 136720 3575 136776
rect -960 136718 3575 136720
rect -960 136628 480 136718
rect 3509 136715 3575 136718
rect 580165 126034 580231 126037
rect 583520 126034 584960 126124
rect 580165 126032 584960 126034
rect 580165 125976 580170 126032
rect 580226 125976 584960 126032
rect 580165 125974 584960 125976
rect 580165 125971 580231 125974
rect 583520 125884 584960 125974
rect -960 123572 480 123812
rect 579797 112842 579863 112845
rect 583520 112842 584960 112932
rect 579797 112840 584960 112842
rect 579797 112784 579802 112840
rect 579858 112784 584960 112840
rect 579797 112782 584960 112784
rect 579797 112779 579863 112782
rect 583520 112692 584960 112782
rect 197 111210 263 111213
rect 197 111208 306 111210
rect 197 111152 202 111208
rect 258 111152 306 111208
rect 197 111147 306 111152
rect 246 110802 306 111147
rect 246 110756 674 110802
rect -960 110742 674 110756
rect -960 110666 480 110742
rect 614 110666 674 110742
rect -960 110606 674 110666
rect -960 110516 480 110606
rect 580165 99514 580231 99517
rect 583520 99514 584960 99604
rect 580165 99512 584960 99514
rect 580165 99456 580170 99512
rect 580226 99456 584960 99512
rect 580165 99454 584960 99456
rect 580165 99451 580231 99454
rect 583520 99364 584960 99454
rect -960 97610 480 97700
rect 3325 97610 3391 97613
rect -960 97608 3391 97610
rect -960 97552 3330 97608
rect 3386 97552 3391 97608
rect -960 97550 3391 97552
rect -960 97460 480 97550
rect 3325 97547 3391 97550
rect 580165 86186 580231 86189
rect 583520 86186 584960 86276
rect 580165 86184 584960 86186
rect 580165 86128 580170 86184
rect 580226 86128 584960 86184
rect 580165 86126 584960 86128
rect 580165 86123 580231 86126
rect 583520 86036 584960 86126
rect -960 84690 480 84780
rect 3785 84690 3851 84693
rect -960 84688 3851 84690
rect -960 84632 3790 84688
rect 3846 84632 3851 84688
rect -960 84630 3851 84632
rect -960 84540 480 84630
rect 3785 84627 3851 84630
rect 580165 72994 580231 72997
rect 583520 72994 584960 73084
rect 580165 72992 584960 72994
rect 580165 72936 580170 72992
rect 580226 72936 584960 72992
rect 580165 72934 584960 72936
rect 580165 72931 580231 72934
rect 583520 72844 584960 72934
rect 105 71906 171 71909
rect 62 71904 171 71906
rect 62 71848 110 71904
rect 166 71848 171 71904
rect 62 71843 171 71848
rect 62 71770 122 71843
rect 62 71724 674 71770
rect -960 71710 674 71724
rect -960 71634 480 71710
rect 614 71634 674 71710
rect -960 71574 674 71634
rect -960 71484 480 71574
rect 580165 59666 580231 59669
rect 583520 59666 584960 59756
rect 580165 59664 584960 59666
rect 580165 59608 580170 59664
rect 580226 59608 584960 59664
rect 580165 59606 584960 59608
rect 580165 59603 580231 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 2221 58578 2287 58581
rect -960 58576 2287 58578
rect -960 58520 2226 58576
rect 2282 58520 2287 58576
rect -960 58518 2287 58520
rect -960 58428 480 58518
rect 2221 58515 2287 58518
rect 580165 46338 580231 46341
rect 583520 46338 584960 46428
rect 580165 46336 584960 46338
rect 580165 46280 580170 46336
rect 580226 46280 584960 46336
rect 580165 46278 584960 46280
rect 580165 46275 580231 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3417 45522 3483 45525
rect -960 45520 3483 45522
rect -960 45464 3422 45520
rect 3478 45464 3483 45520
rect -960 45462 3483 45464
rect -960 45372 480 45462
rect 3417 45459 3483 45462
rect 580165 33146 580231 33149
rect 583520 33146 584960 33236
rect 580165 33144 584960 33146
rect 580165 33088 580170 33144
rect 580226 33088 584960 33144
rect 580165 33086 584960 33088
rect 580165 33083 580231 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 2129 32466 2195 32469
rect -960 32464 2195 32466
rect -960 32408 2134 32464
rect 2190 32408 2195 32464
rect -960 32406 2195 32408
rect -960 32316 480 32406
rect 2129 32403 2195 32406
rect 13 19954 79 19957
rect 13 19952 122 19954
rect 13 19896 18 19952
rect 74 19896 122 19952
rect 13 19891 122 19896
rect 62 19546 122 19891
rect 579981 19818 580047 19821
rect 583520 19818 584960 19908
rect 579981 19816 584960 19818
rect 579981 19760 579986 19816
rect 580042 19760 584960 19816
rect 579981 19758 584960 19760
rect 579981 19755 580047 19758
rect 583520 19668 584960 19758
rect 62 19500 674 19546
rect -960 19486 674 19500
rect -960 19410 480 19486
rect 614 19410 674 19486
rect -960 19350 674 19410
rect -960 19260 480 19350
rect 580165 6626 580231 6629
rect 583520 6626 584960 6716
rect 580165 6624 584960 6626
rect -960 6490 480 6580
rect 580165 6568 580170 6624
rect 580226 6568 584960 6624
rect 580165 6566 584960 6568
rect 580165 6563 580231 6566
rect 2037 6490 2103 6493
rect -960 6488 2103 6490
rect -960 6432 2042 6488
rect 2098 6432 2103 6488
rect 583520 6476 584960 6566
rect -960 6430 2103 6432
rect -960 6340 480 6430
rect 2037 6427 2103 6430
rect 550590 718 553410 778
rect 4061 642 4127 645
rect 7833 642 7899 645
rect 4061 640 7899 642
rect 4061 584 4066 640
rect 4122 584 7838 640
rect 7894 584 7899 640
rect 4061 582 7899 584
rect 4061 579 4127 582
rect 7833 579 7899 582
rect 9949 642 10015 645
rect 13261 642 13327 645
rect 9949 640 13327 642
rect 9949 584 9954 640
rect 10010 584 13266 640
rect 13322 584 13327 640
rect 9949 582 13327 584
rect 9949 579 10015 582
rect 13261 579 13327 582
rect 20621 642 20687 645
rect 23473 642 23539 645
rect 20621 640 23539 642
rect 20621 584 20626 640
rect 20682 584 23478 640
rect 23534 584 23539 640
rect 20621 582 23539 584
rect 20621 579 20687 582
rect 23473 579 23539 582
rect 26509 642 26575 645
rect 28717 642 28783 645
rect 30281 642 30347 645
rect 26509 640 28783 642
rect 26509 584 26514 640
rect 26570 584 28722 640
rect 28778 584 28783 640
rect 26509 582 28783 584
rect 26509 579 26575 582
rect 28717 579 28783 582
rect 29134 640 30347 642
rect 29134 584 30286 640
rect 30342 584 30347 640
rect 29134 582 30347 584
rect 18505 506 18571 509
rect 21265 506 21331 509
rect 18505 504 21331 506
rect 18505 448 18510 504
rect 18566 448 21270 504
rect 21326 448 21331 504
rect 18505 446 21331 448
rect 18505 443 18571 446
rect 21265 443 21331 446
rect 27889 506 27955 509
rect 29134 506 29194 582
rect 30281 579 30347 582
rect 32397 642 32463 645
rect 33225 642 33291 645
rect 32397 640 33291 642
rect 32397 584 32402 640
rect 32458 584 33230 640
rect 33286 584 33291 640
rect 32397 582 33291 584
rect 32397 579 32463 582
rect 33225 579 33291 582
rect 35985 642 36051 645
rect 38469 642 38535 645
rect 35985 640 38535 642
rect 35985 584 35990 640
rect 36046 584 38474 640
rect 38530 584 38535 640
rect 35985 582 38535 584
rect 35985 579 36051 582
rect 38469 579 38535 582
rect 52545 642 52611 645
rect 56041 642 56107 645
rect 57605 642 57671 645
rect 52545 640 53850 642
rect 52545 584 52550 640
rect 52606 584 53850 640
rect 52545 582 53850 584
rect 52545 579 52611 582
rect 27889 504 29194 506
rect 27889 448 27894 504
rect 27950 448 29194 504
rect 27889 446 29194 448
rect 53790 506 53850 582
rect 56041 640 57671 642
rect 56041 584 56046 640
rect 56102 584 57610 640
rect 57666 584 57671 640
rect 56041 582 57671 584
rect 56041 579 56107 582
rect 57605 579 57671 582
rect 58433 642 58499 645
rect 59813 642 59879 645
rect 58433 640 59879 642
rect 58433 584 58438 640
rect 58494 584 59818 640
rect 59874 584 59879 640
rect 58433 582 59879 584
rect 58433 579 58499 582
rect 59813 579 59879 582
rect 62021 642 62087 645
rect 63493 642 63559 645
rect 62021 640 63559 642
rect 62021 584 62026 640
rect 62082 584 63498 640
rect 63554 584 63559 640
rect 62021 582 63559 584
rect 62021 579 62087 582
rect 63493 579 63559 582
rect 142061 642 142127 645
rect 143441 642 143507 645
rect 144729 642 144795 645
rect 142061 640 142170 642
rect 142061 584 142066 640
rect 142122 584 142170 640
rect 142061 579 142170 584
rect 143441 640 144795 642
rect 143441 584 143446 640
rect 143502 584 144734 640
rect 144790 584 144795 640
rect 143441 582 144795 584
rect 143441 579 143507 582
rect 144729 579 144795 582
rect 145741 642 145807 645
rect 147121 642 147187 645
rect 145741 640 147187 642
rect 145741 584 145746 640
rect 145802 584 147126 640
rect 147182 584 147187 640
rect 145741 582 147187 584
rect 145741 579 145807 582
rect 147121 579 147187 582
rect 148961 642 149027 645
rect 150617 642 150683 645
rect 151813 642 151879 645
rect 148961 640 150683 642
rect 148961 584 148966 640
rect 149022 584 150622 640
rect 150678 584 150683 640
rect 148961 582 150683 584
rect 148961 579 149027 582
rect 150617 579 150683 582
rect 151678 640 151879 642
rect 151678 584 151818 640
rect 151874 584 151879 640
rect 151678 582 151879 584
rect 54201 506 54267 509
rect 53790 504 54267 506
rect 53790 448 54206 504
rect 54262 448 54267 504
rect 53790 446 54267 448
rect 27889 443 27955 446
rect 54201 443 54267 446
rect 57421 506 57487 509
rect 58801 506 58867 509
rect 57421 504 58867 506
rect 57421 448 57426 504
rect 57482 448 58806 504
rect 58862 448 58867 504
rect 57421 446 58867 448
rect 57421 443 57487 446
rect 58801 443 58867 446
rect 59445 506 59511 509
rect 61101 506 61167 509
rect 59445 504 61167 506
rect 59445 448 59450 504
rect 59506 448 61106 504
rect 61162 448 61167 504
rect 59445 446 61167 448
rect 142110 506 142170 579
rect 143717 506 143783 509
rect 142110 504 143783 506
rect 142110 448 143722 504
rect 143778 448 143783 504
rect 142110 446 143783 448
rect 59445 443 59511 446
rect 61101 443 61167 446
rect 143717 443 143783 446
rect 147765 506 147831 509
rect 149329 506 149395 509
rect 147765 504 149395 506
rect 147765 448 147770 504
rect 147826 448 149334 504
rect 149390 448 149395 504
rect 147765 446 149395 448
rect 147765 443 147831 446
rect 149329 443 149395 446
rect 150249 506 150315 509
rect 151678 506 151738 582
rect 151813 579 151879 582
rect 164785 642 164851 645
rect 167361 642 167427 645
rect 164785 640 167427 642
rect 164785 584 164790 640
rect 164846 584 167366 640
rect 167422 584 167427 640
rect 164785 582 167427 584
rect 164785 579 164851 582
rect 167361 579 167427 582
rect 169477 642 169543 645
rect 171961 642 172027 645
rect 169477 640 172027 642
rect 169477 584 169482 640
rect 169538 584 171966 640
rect 172022 584 172027 640
rect 169477 582 172027 584
rect 169477 579 169543 582
rect 171961 579 172027 582
rect 172973 642 173039 645
rect 175457 642 175523 645
rect 172973 640 175523 642
rect 172973 584 172978 640
rect 173034 584 175462 640
rect 175518 584 175523 640
rect 172973 582 175523 584
rect 172973 579 173039 582
rect 175457 579 175523 582
rect 176377 642 176443 645
rect 179045 642 179111 645
rect 180241 642 180307 645
rect 176377 640 179111 642
rect 176377 584 176382 640
rect 176438 584 179050 640
rect 179106 584 179111 640
rect 176377 582 179111 584
rect 176377 579 176443 582
rect 179045 579 179111 582
rect 179370 640 180307 642
rect 179370 584 180246 640
rect 180302 584 180307 640
rect 179370 582 180307 584
rect 150249 504 151738 506
rect 150249 448 150254 504
rect 150310 448 151738 504
rect 150249 446 151738 448
rect 173893 506 173959 509
rect 176837 506 176903 509
rect 173893 504 176903 506
rect 173893 448 173898 504
rect 173954 448 176842 504
rect 176898 448 176903 504
rect 173893 446 176903 448
rect 150249 443 150315 446
rect 173893 443 173959 446
rect 176837 443 176903 446
rect 177481 506 177547 509
rect 179370 506 179430 582
rect 180241 579 180307 582
rect 182081 642 182147 645
rect 184933 642 184999 645
rect 182081 640 184999 642
rect 182081 584 182086 640
rect 182142 584 184938 640
rect 184994 584 184999 640
rect 182081 582 184999 584
rect 182081 579 182147 582
rect 184933 579 184999 582
rect 191097 642 191163 645
rect 194409 642 194475 645
rect 191097 640 194475 642
rect 191097 584 191102 640
rect 191158 584 194414 640
rect 194470 584 194475 640
rect 191097 582 194475 584
rect 191097 579 191163 582
rect 194409 579 194475 582
rect 196709 642 196775 645
rect 200297 642 200363 645
rect 201493 642 201559 645
rect 196709 640 200363 642
rect 196709 584 196714 640
rect 196770 584 200302 640
rect 200358 584 200363 640
rect 196709 582 200363 584
rect 196709 579 196775 582
rect 200297 579 200363 582
rect 201358 640 201559 642
rect 201358 584 201498 640
rect 201554 584 201559 640
rect 201358 582 201559 584
rect 177481 504 179430 506
rect 177481 448 177486 504
rect 177542 448 179430 504
rect 177481 446 179430 448
rect 186589 506 186655 509
rect 189901 506 189967 509
rect 201358 506 201418 582
rect 201493 579 201559 582
rect 203609 642 203675 645
rect 207381 642 207447 645
rect 208577 642 208643 645
rect 203609 640 207447 642
rect 203609 584 203614 640
rect 203670 584 207386 640
rect 207442 584 207447 640
rect 203609 582 207447 584
rect 203609 579 203675 582
rect 207381 579 207447 582
rect 207982 640 208643 642
rect 207982 584 208582 640
rect 208638 584 208643 640
rect 207982 582 208643 584
rect 186589 504 189967 506
rect 186589 448 186594 504
rect 186650 448 189906 504
rect 189962 448 189967 504
rect 186589 446 189967 448
rect 177481 443 177547 446
rect 186589 443 186655 446
rect 189901 443 189967 446
rect 198782 446 201418 506
rect 201861 506 201927 509
rect 203701 506 203767 509
rect 201861 504 203767 506
rect 201861 448 201866 504
rect 201922 448 203706 504
rect 203762 448 203767 504
rect 201861 446 203767 448
rect 168189 370 168255 373
rect 170949 370 171015 373
rect 168189 368 171015 370
rect 168189 312 168194 368
rect 168250 312 170954 368
rect 171010 312 171015 368
rect 168189 310 171015 312
rect 168189 307 168255 310
rect 170949 307 171015 310
rect 171685 370 171751 373
rect 173985 370 174051 373
rect 171685 368 174051 370
rect 171685 312 171690 368
rect 171746 312 173990 368
rect 174046 312 174051 368
rect 171685 310 174051 312
rect 171685 307 171751 310
rect 173985 307 174051 310
rect 175181 370 175247 373
rect 177665 370 177731 373
rect 175181 368 177731 370
rect 175181 312 175186 368
rect 175242 312 177670 368
rect 177726 312 177731 368
rect 175181 310 177731 312
rect 175181 307 175247 310
rect 177665 307 177731 310
rect 178677 370 178743 373
rect 181253 370 181319 373
rect 178677 368 181319 370
rect 178677 312 178682 368
rect 178738 312 181258 368
rect 181314 312 181319 368
rect 178677 310 181319 312
rect 178677 307 178743 310
rect 181253 307 181319 310
rect 197721 370 197787 373
rect 198782 370 198842 446
rect 201861 443 201927 446
rect 203701 443 203767 446
rect 204805 506 204871 509
rect 207982 506 208042 582
rect 208577 579 208643 582
rect 209313 642 209379 645
rect 213361 642 213427 645
rect 209313 640 213427 642
rect 209313 584 209318 640
rect 209374 584 213366 640
rect 213422 584 213427 640
rect 209313 582 213427 584
rect 209313 579 209379 582
rect 213361 579 213427 582
rect 222469 642 222535 645
rect 227529 642 227595 645
rect 228725 642 228791 645
rect 222469 640 227595 642
rect 222469 584 222474 640
rect 222530 584 227534 640
rect 227590 584 227595 640
rect 222469 582 227595 584
rect 222469 579 222535 582
rect 227529 579 227595 582
rect 227670 640 228791 642
rect 227670 584 228730 640
rect 228786 584 228791 640
rect 227670 582 228791 584
rect 204805 504 208042 506
rect 204805 448 204810 504
rect 204866 448 208042 504
rect 204805 446 208042 448
rect 208209 506 208275 509
rect 211981 506 212047 509
rect 208209 504 212047 506
rect 208209 448 208214 504
rect 208270 448 211986 504
rect 212042 448 212047 504
rect 208209 446 212047 448
rect 204805 443 204871 446
rect 208209 443 208275 446
rect 211981 443 212047 446
rect 216121 506 216187 509
rect 220169 506 220235 509
rect 216121 504 220235 506
rect 216121 448 216126 504
rect 216182 448 220174 504
rect 220230 448 220235 504
rect 216121 446 220235 448
rect 216121 443 216187 446
rect 220169 443 220235 446
rect 223573 506 223639 509
rect 227670 506 227730 582
rect 228725 579 228791 582
rect 230933 642 230999 645
rect 235809 642 235875 645
rect 230933 640 235875 642
rect 230933 584 230938 640
rect 230994 584 235814 640
rect 235870 584 235875 640
rect 230933 582 235875 584
rect 230933 579 230999 582
rect 235809 579 235875 582
rect 238845 642 238911 645
rect 244089 642 244155 645
rect 238845 640 244155 642
rect 238845 584 238850 640
rect 238906 584 244094 640
rect 244150 584 244155 640
rect 238845 582 244155 584
rect 238845 579 238911 582
rect 244089 579 244155 582
rect 249057 642 249123 645
rect 254669 642 254735 645
rect 255865 642 255931 645
rect 249057 640 254735 642
rect 249057 584 249062 640
rect 249118 584 254674 640
rect 254730 584 254735 640
rect 249057 582 254735 584
rect 249057 579 249123 582
rect 254669 579 254735 582
rect 255822 640 255931 642
rect 255822 584 255870 640
rect 255926 584 255931 640
rect 255822 579 255931 584
rect 263133 642 263199 645
rect 264145 642 264211 645
rect 263133 640 264211 642
rect 263133 584 263138 640
rect 263194 584 264150 640
rect 264206 584 264211 640
rect 263133 582 264211 584
rect 263133 579 263199 582
rect 264145 579 264211 582
rect 267273 642 267339 645
rect 273621 642 273687 645
rect 267273 640 273687 642
rect 267273 584 267278 640
rect 267334 584 273626 640
rect 273682 584 273687 640
rect 267273 582 273687 584
rect 267273 579 267339 582
rect 273621 579 273687 582
rect 275829 642 275895 645
rect 283097 642 283163 645
rect 286593 642 286659 645
rect 275829 640 283163 642
rect 275829 584 275834 640
rect 275890 584 283102 640
rect 283158 584 283163 640
rect 275829 582 283163 584
rect 275829 579 275895 582
rect 283097 579 283163 582
rect 283238 640 286659 642
rect 283238 584 286598 640
rect 286654 584 286659 640
rect 283238 582 286659 584
rect 223573 504 227730 506
rect 223573 448 223578 504
rect 223634 448 227730 504
rect 223573 446 227730 448
rect 243353 506 243419 509
rect 248965 506 249031 509
rect 243353 504 249031 506
rect 243353 448 243358 504
rect 243414 448 248970 504
rect 249026 448 249031 504
rect 243353 446 249031 448
rect 223573 443 223639 446
rect 243353 443 243419 446
rect 248965 443 249031 446
rect 249701 506 249767 509
rect 255822 506 255882 579
rect 249701 504 255882 506
rect 249701 448 249706 504
rect 249762 448 255882 504
rect 249701 446 255882 448
rect 275185 506 275251 509
rect 282177 506 282243 509
rect 275185 504 282243 506
rect 275185 448 275190 504
rect 275246 448 282182 504
rect 282238 448 282243 504
rect 275185 446 282243 448
rect 249701 443 249767 446
rect 275185 443 275251 446
rect 282177 443 282243 446
rect 197721 368 198842 370
rect 197721 312 197726 368
rect 197782 312 198842 368
rect 197721 310 198842 312
rect 200021 370 200087 373
rect 201309 370 201375 373
rect 204897 370 204963 373
rect 200021 368 200130 370
rect 200021 312 200026 368
rect 200082 312 200130 368
rect 197721 307 197787 310
rect 200021 307 200130 312
rect 201309 368 204963 370
rect 201309 312 201314 368
rect 201370 312 204902 368
rect 204958 312 204963 368
rect 201309 310 204963 312
rect 201309 307 201375 310
rect 204897 307 204963 310
rect 206921 370 206987 373
rect 210785 370 210851 373
rect 206921 368 210851 370
rect 206921 312 206926 368
rect 206982 312 210790 368
rect 210846 312 210851 368
rect 206921 310 210851 312
rect 206921 307 206987 310
rect 210785 307 210851 310
rect 217225 370 217291 373
rect 221733 370 221799 373
rect 217225 368 221799 370
rect 217225 312 217230 368
rect 217286 312 221738 368
rect 221794 312 221799 368
rect 217225 310 221799 312
rect 217225 307 217291 310
rect 221733 307 221799 310
rect 279233 370 279299 373
rect 283238 370 283298 582
rect 286593 579 286659 582
rect 287053 642 287119 645
rect 287789 642 287855 645
rect 287053 640 287855 642
rect 287053 584 287058 640
rect 287114 584 287794 640
rect 287850 584 287855 640
rect 287053 582 287855 584
rect 287053 579 287119 582
rect 287789 579 287855 582
rect 291561 642 291627 645
rect 293677 642 293743 645
rect 291561 640 293743 642
rect 291561 584 291566 640
rect 291622 584 293682 640
rect 293738 584 293743 640
rect 291561 582 293743 584
rect 291561 579 291627 582
rect 293677 579 293743 582
rect 293861 642 293927 645
rect 294873 642 294939 645
rect 293861 640 294939 642
rect 293861 584 293866 640
rect 293922 584 294878 640
rect 294934 584 294939 640
rect 293861 582 294939 584
rect 293861 579 293927 582
rect 294873 579 294939 582
rect 305821 642 305887 645
rect 313825 642 313891 645
rect 305821 640 313891 642
rect 305821 584 305826 640
rect 305882 584 313830 640
rect 313886 584 313891 640
rect 305821 582 313891 584
rect 305821 579 305887 582
rect 313825 579 313891 582
rect 315021 640 315087 645
rect 315021 584 315026 640
rect 315082 584 315087 640
rect 315021 579 315087 584
rect 316585 642 316651 645
rect 317321 642 317387 645
rect 316585 640 317387 642
rect 316585 584 316590 640
rect 316646 584 317326 640
rect 317382 584 317387 640
rect 316585 582 317387 584
rect 316585 579 316651 582
rect 317321 579 317387 582
rect 334249 642 334315 645
rect 343357 642 343423 645
rect 344553 642 344619 645
rect 345749 642 345815 645
rect 334249 640 343423 642
rect 334249 584 334254 640
rect 334310 584 343362 640
rect 343418 584 343423 640
rect 334249 582 343423 584
rect 334249 579 334315 582
rect 343357 579 343423 582
rect 343590 640 344619 642
rect 343590 584 344558 640
rect 344614 584 344619 640
rect 343590 582 344619 584
rect 285213 506 285279 509
rect 292757 506 292823 509
rect 285213 504 292823 506
rect 285213 448 285218 504
rect 285274 448 292762 504
rect 292818 448 292823 504
rect 285213 446 292823 448
rect 285213 443 285279 446
rect 292757 443 292823 446
rect 307017 506 307083 509
rect 315024 506 315084 579
rect 307017 504 315084 506
rect 307017 448 307022 504
rect 307078 448 315084 504
rect 307017 446 315084 448
rect 335353 506 335419 509
rect 343590 506 343650 582
rect 344553 579 344619 582
rect 344970 640 345815 642
rect 344970 584 345754 640
rect 345810 584 345815 640
rect 344970 582 345815 584
rect 335353 504 343650 506
rect 335353 448 335358 504
rect 335414 448 343650 504
rect 335353 446 343650 448
rect 307017 443 307083 446
rect 335353 443 335419 446
rect 279233 368 283298 370
rect 279233 312 279238 368
rect 279294 312 283298 368
rect 279233 310 283298 312
rect 326337 370 326403 373
rect 335261 370 335327 373
rect 326337 368 335327 370
rect 326337 312 326342 368
rect 326398 312 335266 368
rect 335322 312 335327 368
rect 326337 310 335327 312
rect 279233 307 279299 310
rect 326337 307 326403 310
rect 335261 307 335327 310
rect 336549 370 336615 373
rect 344970 370 345030 582
rect 345749 579 345815 582
rect 345933 642 345999 645
rect 346945 642 347011 645
rect 345933 640 347011 642
rect 345933 584 345938 640
rect 345994 584 346950 640
rect 347006 584 347011 640
rect 345933 582 347011 584
rect 345933 579 345999 582
rect 346945 579 347011 582
rect 347773 642 347839 645
rect 350441 642 350507 645
rect 347773 640 350507 642
rect 347773 584 347778 640
rect 347834 584 350446 640
rect 350502 584 350507 640
rect 347773 582 350507 584
rect 347773 579 347839 582
rect 350441 579 350507 582
rect 351821 642 351887 645
rect 352833 642 352899 645
rect 351821 640 352899 642
rect 351821 584 351826 640
rect 351882 584 352838 640
rect 352894 584 352899 640
rect 351821 582 352899 584
rect 351821 579 351887 582
rect 352833 579 352899 582
rect 364425 642 364491 645
rect 375281 642 375347 645
rect 376477 642 376543 645
rect 364425 640 375347 642
rect 364425 584 364430 640
rect 364486 584 375286 640
rect 375342 584 375347 640
rect 364425 582 375347 584
rect 364425 579 364491 582
rect 375281 579 375347 582
rect 375422 640 376543 642
rect 375422 584 376482 640
rect 376538 584 376543 640
rect 375422 582 376543 584
rect 366081 506 366147 509
rect 375422 506 375482 582
rect 376477 579 376543 582
rect 393773 642 393839 645
rect 401317 642 401383 645
rect 393773 640 401383 642
rect 393773 584 393778 640
rect 393834 584 401322 640
rect 401378 584 401383 640
rect 393773 582 401383 584
rect 393773 579 393839 582
rect 401317 579 401383 582
rect 421097 642 421163 645
rect 424961 642 425027 645
rect 421097 640 425027 642
rect 421097 584 421102 640
rect 421158 584 424966 640
rect 425022 584 425027 640
rect 421097 582 425027 584
rect 421097 579 421163 582
rect 424961 579 425027 582
rect 425513 642 425579 645
rect 426157 642 426223 645
rect 429653 642 429719 645
rect 425513 640 426223 642
rect 425513 584 425518 640
rect 425574 584 426162 640
rect 426218 584 426223 640
rect 425513 582 426223 584
rect 425513 579 425579 582
rect 426157 579 426223 582
rect 426390 640 429719 642
rect 426390 584 429658 640
rect 429714 584 429719 640
rect 426390 582 429719 584
rect 366081 504 375482 506
rect 366081 448 366086 504
rect 366142 448 375482 504
rect 366081 446 375482 448
rect 384205 506 384271 509
rect 389817 506 389883 509
rect 384205 504 389883 506
rect 384205 448 384210 504
rect 384266 448 389822 504
rect 389878 448 389883 504
rect 384205 446 389883 448
rect 366081 443 366147 446
rect 384205 443 384271 446
rect 389817 443 389883 446
rect 392209 506 392275 509
rect 400305 506 400371 509
rect 392209 504 400371 506
rect 392209 448 392214 504
rect 392270 448 400310 504
rect 400366 448 400371 504
rect 392209 446 400371 448
rect 392209 443 392275 446
rect 400305 443 400371 446
rect 417141 506 417207 509
rect 426390 506 426450 582
rect 429653 579 429719 582
rect 445569 642 445635 645
rect 459185 642 459251 645
rect 445569 640 459251 642
rect 445569 584 445574 640
rect 445630 584 459190 640
rect 459246 584 459251 640
rect 445569 582 459251 584
rect 445569 579 445635 582
rect 459185 579 459251 582
rect 459553 642 459619 645
rect 461577 642 461643 645
rect 459553 640 461643 642
rect 459553 584 459558 640
rect 459614 584 461582 640
rect 461638 584 461643 640
rect 459553 582 461643 584
rect 459553 579 459619 582
rect 461577 579 461643 582
rect 463049 642 463115 645
rect 465165 642 465231 645
rect 463049 640 465231 642
rect 463049 584 463054 640
rect 463110 584 465170 640
rect 465226 584 465231 640
rect 463049 582 465231 584
rect 463049 579 463115 582
rect 465165 579 465231 582
rect 465349 642 465415 645
rect 466177 642 466243 645
rect 465349 640 466243 642
rect 465349 584 465354 640
rect 465410 584 466182 640
rect 466238 584 466243 640
rect 465349 582 466243 584
rect 465349 579 465415 582
rect 466177 579 466243 582
rect 466361 642 466427 645
rect 467465 642 467531 645
rect 471053 642 471119 645
rect 466361 640 467531 642
rect 466361 584 466366 640
rect 466422 584 467470 640
rect 467526 584 467531 640
rect 466361 582 467531 584
rect 466361 579 466427 582
rect 467465 579 467531 582
rect 469170 640 471119 642
rect 469170 584 471058 640
rect 471114 584 471119 640
rect 469170 582 471119 584
rect 417141 504 426450 506
rect 417141 448 417146 504
rect 417202 448 426450 504
rect 417141 446 426450 448
rect 460657 506 460723 509
rect 463785 506 463851 509
rect 460657 504 463851 506
rect 460657 448 460662 504
rect 460718 448 463790 504
rect 463846 448 463851 504
rect 460657 446 463851 448
rect 417141 443 417207 446
rect 460657 443 460723 446
rect 463785 443 463851 446
rect 467833 506 467899 509
rect 469170 506 469230 582
rect 471053 579 471119 582
rect 475101 642 475167 645
rect 489913 642 489979 645
rect 492305 642 492371 645
rect 475101 640 489979 642
rect 475101 584 475106 640
rect 475162 584 489918 640
rect 489974 584 489979 640
rect 475101 582 489979 584
rect 475101 579 475167 582
rect 489913 579 489979 582
rect 492262 640 492371 642
rect 492262 584 492310 640
rect 492366 584 492371 640
rect 492262 579 492371 584
rect 492673 642 492739 645
rect 495893 642 495959 645
rect 492673 640 495959 642
rect 492673 584 492678 640
rect 492734 584 495898 640
rect 495954 584 495959 640
rect 492673 582 495959 584
rect 492673 579 492739 582
rect 495893 579 495959 582
rect 496813 642 496879 645
rect 500585 642 500651 645
rect 496813 640 500651 642
rect 496813 584 496818 640
rect 496874 584 500590 640
rect 500646 584 500651 640
rect 496813 582 500651 584
rect 496813 579 496879 582
rect 500585 579 500651 582
rect 509693 642 509759 645
rect 531129 642 531195 645
rect 533705 642 533771 645
rect 509693 640 517162 642
rect 509693 584 509698 640
rect 509754 611 517162 640
rect 531129 640 533771 642
rect 509754 606 517211 611
rect 509754 584 517150 606
rect 509693 582 517150 584
rect 509693 579 509759 582
rect 467833 504 469230 506
rect 467833 448 467838 504
rect 467894 448 469230 504
rect 467833 446 469230 448
rect 473997 506 474063 509
rect 488625 506 488691 509
rect 473997 504 488691 506
rect 473997 448 474002 504
rect 474058 448 488630 504
rect 488686 448 488691 504
rect 473997 446 488691 448
rect 467833 443 467899 446
rect 473997 443 474063 446
rect 488625 443 488691 446
rect 489269 506 489335 509
rect 492262 506 492322 579
rect 517102 550 517150 582
rect 517206 550 517211 606
rect 531129 584 531134 640
rect 531190 584 533710 640
rect 533766 584 533771 640
rect 531129 582 533771 584
rect 531129 579 531195 582
rect 533705 579 533771 582
rect 534165 642 534231 645
rect 548149 642 548215 645
rect 534165 640 548215 642
rect 534165 584 534170 640
rect 534226 584 548154 640
rect 548210 584 548215 640
rect 534165 582 548215 584
rect 534165 579 534231 582
rect 548149 579 548215 582
rect 548333 642 548399 645
rect 549069 642 549135 645
rect 548333 640 549135 642
rect 548333 584 548338 640
rect 548394 584 549074 640
rect 549130 584 549135 640
rect 548333 582 549135 584
rect 548333 579 548399 582
rect 549069 579 549135 582
rect 549253 642 549319 645
rect 550590 642 550650 718
rect 549253 640 550650 642
rect 549253 584 549258 640
rect 549314 584 550650 640
rect 549253 582 550650 584
rect 553350 642 553410 718
rect 559741 642 559807 645
rect 553350 640 559807 642
rect 553350 584 559746 640
rect 559802 584 559807 640
rect 553350 582 559807 584
rect 549253 579 549319 582
rect 559741 579 559807 582
rect 517102 548 517211 550
rect 517145 545 517211 548
rect 489269 504 492322 506
rect 489269 448 489274 504
rect 489330 448 492322 504
rect 489269 446 492322 448
rect 492673 506 492739 509
rect 494513 506 494579 509
rect 492673 504 494579 506
rect 492673 448 492678 504
rect 492734 448 494518 504
rect 494574 448 494579 504
rect 492673 446 494579 448
rect 489269 443 489335 446
rect 492673 443 492739 446
rect 494513 443 494579 446
rect 495525 506 495591 509
rect 499021 506 499087 509
rect 495525 504 499087 506
rect 495525 448 495530 504
rect 495586 448 499026 504
rect 499082 448 499087 504
rect 495525 446 499087 448
rect 495525 443 495591 446
rect 499021 443 499087 446
rect 501229 506 501295 509
rect 506933 506 506999 509
rect 501229 504 506999 506
rect 501229 448 501234 504
rect 501290 448 506938 504
rect 506994 448 506999 504
rect 501229 446 506999 448
rect 501229 443 501295 446
rect 506933 443 506999 446
rect 540513 506 540579 509
rect 558361 506 558427 509
rect 540513 504 558427 506
rect 540513 448 540518 504
rect 540574 448 558366 504
rect 558422 448 558427 504
rect 540513 446 558427 448
rect 540513 443 540579 446
rect 558361 443 558427 446
rect 336549 368 345030 370
rect 336549 312 336554 368
rect 336610 312 345030 368
rect 336549 310 345030 312
rect 383101 370 383167 373
rect 386965 370 387031 373
rect 383101 368 387031 370
rect 383101 312 383106 368
rect 383162 312 386970 368
rect 387026 312 387031 368
rect 383101 310 387031 312
rect 336549 307 336615 310
rect 383101 307 383167 310
rect 386965 307 387031 310
rect 479609 370 479675 373
rect 487797 370 487863 373
rect 479609 368 487863 370
rect 479609 312 479614 368
rect 479670 312 487802 368
rect 487858 312 487863 368
rect 479609 310 487863 312
rect 479609 307 479675 310
rect 487797 307 487863 310
rect 490281 370 490347 373
rect 493317 370 493383 373
rect 490281 368 493383 370
rect 490281 312 490286 368
rect 490342 312 493322 368
rect 493378 312 493383 368
rect 490281 310 493383 312
rect 490281 307 490347 310
rect 493317 307 493383 310
rect 537569 370 537635 373
rect 554773 370 554839 373
rect 537569 368 554839 370
rect 537569 312 537574 368
rect 537630 312 554778 368
rect 554834 312 554839 368
rect 537569 310 554839 312
rect 537569 307 537635 310
rect 554773 307 554839 310
rect 195237 234 195303 237
rect 198917 234 198983 237
rect 195237 232 198983 234
rect 195237 176 195242 232
rect 195298 176 198922 232
rect 198978 176 198983 232
rect 195237 174 198983 176
rect 200070 234 200130 307
rect 201861 234 201927 237
rect 200070 232 201927 234
rect 200070 176 201866 232
rect 201922 176 201927 232
rect 200070 174 201927 176
rect 195237 171 195303 174
rect 198917 171 198983 174
rect 201861 171 201927 174
rect 202413 234 202479 237
rect 206001 234 206067 237
rect 202413 232 206067 234
rect 202413 176 202418 232
rect 202474 176 206006 232
rect 206062 176 206067 232
rect 202413 174 206067 176
rect 202413 171 202479 174
rect 206001 171 206067 174
rect 385769 234 385835 237
rect 391565 234 391631 237
rect 385769 232 391631 234
rect 385769 176 385774 232
rect 385830 176 391570 232
rect 391626 176 391631 232
rect 385769 174 391631 176
rect 385769 171 385835 174
rect 391565 171 391631 174
rect 502701 234 502767 237
rect 507301 234 507367 237
rect 502701 232 507367 234
rect 502701 176 502706 232
rect 502762 176 507306 232
rect 507362 176 507367 232
rect 502701 174 507367 176
rect 502701 171 502767 174
rect 507301 171 507367 174
rect 530761 234 530827 237
rect 548057 234 548123 237
rect 530761 232 548123 234
rect 530761 176 530766 232
rect 530822 176 548062 232
rect 548118 176 548123 232
rect 530761 174 548123 176
rect 530761 171 530827 174
rect 548057 171 548123 174
rect 548241 234 548307 237
rect 551277 234 551343 237
rect 548241 232 551343 234
rect 548241 176 548246 232
rect 548302 176 551282 232
rect 551338 176 551343 232
rect 548241 174 551343 176
rect 548241 171 548307 174
rect 551277 171 551343 174
rect 198917 98 198983 101
rect 202505 98 202571 101
rect 198917 96 202571 98
rect 198917 40 198922 96
rect 198978 40 202510 96
rect 202566 40 202571 96
rect 198917 38 202571 40
rect 198917 35 198983 38
rect 202505 35 202571 38
rect 535269 98 535335 101
rect 552381 98 552447 101
rect 535269 96 552447 98
rect 535269 40 535274 96
rect 535330 40 552386 96
rect 552442 40 552447 96
rect 535269 38 552447 40
rect 535269 35 535335 38
rect 552381 35 552447 38
<< via3 >>
rect 164188 701116 164252 701180
rect 433380 699544 433444 699548
rect 433380 699488 433430 699544
rect 433430 699488 433444 699544
rect 433380 699484 433444 699488
rect 11468 699348 11532 699412
rect 13860 699348 13924 699412
rect 21404 699348 21468 699412
rect 30972 699348 31036 699412
rect 33364 699348 33428 699412
rect 43116 699348 43180 699412
rect 408908 699408 408972 699412
rect 408908 699352 408958 699408
rect 408958 699352 408972 699408
rect 408908 699348 408972 699352
rect 418660 699408 418724 699412
rect 418660 699352 418710 699408
rect 418710 699352 418724 699408
rect 418660 699348 418724 699352
rect 448100 699408 448164 699412
rect 448100 699352 448150 699408
rect 448150 699352 448164 699408
rect 164188 699212 164252 699276
rect 409092 699212 409156 699276
rect 448100 699348 448164 699352
rect 453068 699408 453132 699412
rect 453068 699352 453118 699408
rect 453118 699352 453132 699408
rect 453068 699348 453132 699352
rect 43116 698940 43180 699004
rect 33364 698804 33428 698868
rect 30972 698668 31036 698732
rect 21404 698532 21468 698596
rect 13860 698396 13924 698460
rect 11468 698260 11532 698324
rect 418660 698124 418724 698188
rect 408908 697988 408972 698052
rect 409092 697988 409156 698052
rect 433380 697852 433444 697916
rect 448100 697716 448164 697780
rect 453068 697580 453132 697644
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 680614 -8106 711002
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 -8106 680614
rect -8726 680294 -8106 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 -8106 680294
rect -8726 644614 -8106 680058
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 -8106 644614
rect -8726 644294 -8106 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 -8106 644294
rect -8726 608614 -8106 644058
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 -8106 608614
rect -8726 608294 -8106 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 -8106 608294
rect -8726 572614 -8106 608058
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 -8106 572614
rect -8726 572294 -8106 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 -8106 572294
rect -8726 536614 -8106 572058
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 -8106 536614
rect -8726 536294 -8106 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 -8106 536294
rect -8726 500614 -8106 536058
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 -8106 500614
rect -8726 500294 -8106 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 -8106 500294
rect -8726 464614 -8106 500058
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 -8106 464614
rect -8726 464294 -8106 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 -8106 464294
rect -8726 428614 -8106 464058
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 -8106 428614
rect -8726 428294 -8106 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 -8106 428294
rect -8726 392614 -8106 428058
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 -8106 392614
rect -8726 392294 -8106 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 -8106 392294
rect -8726 356614 -8106 392058
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 -8106 356614
rect -8726 356294 -8106 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 -8106 356294
rect -8726 320614 -8106 356058
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 -8106 320614
rect -8726 320294 -8106 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 -8106 320294
rect -8726 284614 -8106 320058
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 -8106 284614
rect -8726 284294 -8106 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 -8106 284294
rect -8726 248614 -8106 284058
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 -8106 248614
rect -8726 248294 -8106 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 -8106 248294
rect -8726 212614 -8106 248058
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 -8106 212614
rect -8726 212294 -8106 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 -8106 212294
rect -8726 176614 -8106 212058
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 -8106 176614
rect -8726 176294 -8106 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 -8106 176294
rect -8726 140614 -8106 176058
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 -8106 140614
rect -8726 140294 -8106 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 -8106 140294
rect -8726 104614 -8106 140058
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 -8106 104614
rect -8726 104294 -8106 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 -8106 104294
rect -8726 68614 -8106 104058
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 -8106 68614
rect -8726 68294 -8106 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 -8106 68294
rect -8726 32614 -8106 68058
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 -8106 32614
rect -8726 32294 -8106 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 -8106 32294
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 13574 710598
rect 12954 710278 13574 710362
rect 12954 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 13574 710278
rect -7766 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 -7146 698614
rect -7766 698294 -7146 698378
rect -7766 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 -7146 698294
rect -7766 662614 -7146 698058
rect -7766 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 -7146 662614
rect -7766 662294 -7146 662378
rect -7766 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 -7146 662294
rect -7766 626614 -7146 662058
rect -7766 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 -7146 626614
rect -7766 626294 -7146 626378
rect -7766 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 -7146 626294
rect -7766 590614 -7146 626058
rect -7766 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 -7146 590614
rect -7766 590294 -7146 590378
rect -7766 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 -7146 590294
rect -7766 554614 -7146 590058
rect -7766 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 -7146 554614
rect -7766 554294 -7146 554378
rect -7766 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 -7146 554294
rect -7766 518614 -7146 554058
rect -7766 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 -7146 518614
rect -7766 518294 -7146 518378
rect -7766 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 -7146 518294
rect -7766 482614 -7146 518058
rect -7766 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 -7146 482614
rect -7766 482294 -7146 482378
rect -7766 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 -7146 482294
rect -7766 446614 -7146 482058
rect -7766 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 -7146 446614
rect -7766 446294 -7146 446378
rect -7766 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 -7146 446294
rect -7766 410614 -7146 446058
rect -7766 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 -7146 410614
rect -7766 410294 -7146 410378
rect -7766 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 -7146 410294
rect -7766 374614 -7146 410058
rect -7766 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 -7146 374614
rect -7766 374294 -7146 374378
rect -7766 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 -7146 374294
rect -7766 338614 -7146 374058
rect -7766 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 -7146 338614
rect -7766 338294 -7146 338378
rect -7766 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 -7146 338294
rect -7766 302614 -7146 338058
rect -7766 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 -7146 302614
rect -7766 302294 -7146 302378
rect -7766 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 -7146 302294
rect -7766 266614 -7146 302058
rect -7766 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 -7146 266614
rect -7766 266294 -7146 266378
rect -7766 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 -7146 266294
rect -7766 230614 -7146 266058
rect -7766 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 -7146 230614
rect -7766 230294 -7146 230378
rect -7766 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 -7146 230294
rect -7766 194614 -7146 230058
rect -7766 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 -7146 194614
rect -7766 194294 -7146 194378
rect -7766 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 -7146 194294
rect -7766 158614 -7146 194058
rect -7766 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 -7146 158614
rect -7766 158294 -7146 158378
rect -7766 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 -7146 158294
rect -7766 122614 -7146 158058
rect -7766 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 -7146 122614
rect -7766 122294 -7146 122378
rect -7766 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 -7146 122294
rect -7766 86614 -7146 122058
rect -7766 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 -7146 86614
rect -7766 86294 -7146 86378
rect -7766 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 -7146 86294
rect -7766 50614 -7146 86058
rect -7766 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 -7146 50614
rect -7766 50294 -7146 50378
rect -7766 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 -7146 50294
rect -7766 14614 -7146 50058
rect -7766 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 -7146 14614
rect -7766 14294 -7146 14378
rect -7766 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 -7146 14294
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 676894 -6186 709082
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 -6186 676894
rect -6806 676574 -6186 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 -6186 676574
rect -6806 640894 -6186 676338
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 -6186 640894
rect -6806 640574 -6186 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 -6186 640574
rect -6806 604894 -6186 640338
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 -6186 604894
rect -6806 604574 -6186 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 -6186 604574
rect -6806 568894 -6186 604338
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 -6186 568894
rect -6806 568574 -6186 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 -6186 568574
rect -6806 532894 -6186 568338
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 -6186 532894
rect -6806 532574 -6186 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 -6186 532574
rect -6806 496894 -6186 532338
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 -6186 496894
rect -6806 496574 -6186 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 -6186 496574
rect -6806 460894 -6186 496338
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 -6186 460894
rect -6806 460574 -6186 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 -6186 460574
rect -6806 424894 -6186 460338
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 -6186 424894
rect -6806 424574 -6186 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 -6186 424574
rect -6806 388894 -6186 424338
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 -6186 388894
rect -6806 388574 -6186 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 -6186 388574
rect -6806 352894 -6186 388338
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 -6186 352894
rect -6806 352574 -6186 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 -6186 352574
rect -6806 316894 -6186 352338
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 -6186 316894
rect -6806 316574 -6186 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 -6186 316574
rect -6806 280894 -6186 316338
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 -6186 280894
rect -6806 280574 -6186 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 -6186 280574
rect -6806 244894 -6186 280338
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 -6186 244894
rect -6806 244574 -6186 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 -6186 244574
rect -6806 208894 -6186 244338
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 -6186 208894
rect -6806 208574 -6186 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 -6186 208574
rect -6806 172894 -6186 208338
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 -6186 172894
rect -6806 172574 -6186 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 -6186 172574
rect -6806 136894 -6186 172338
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 -6186 136894
rect -6806 136574 -6186 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 -6186 136574
rect -6806 100894 -6186 136338
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 -6186 100894
rect -6806 100574 -6186 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 -6186 100574
rect -6806 64894 -6186 100338
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 -6186 64894
rect -6806 64574 -6186 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 -6186 64574
rect -6806 28894 -6186 64338
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 -6186 28894
rect -6806 28574 -6186 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 -6186 28574
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 9854 708678
rect 9234 708358 9854 708442
rect 9234 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 9854 708358
rect -5846 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 -5226 694894
rect -5846 694574 -5226 694658
rect -5846 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 -5226 694574
rect -5846 658894 -5226 694338
rect -5846 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 -5226 658894
rect -5846 658574 -5226 658658
rect -5846 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 -5226 658574
rect -5846 622894 -5226 658338
rect -5846 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 -5226 622894
rect -5846 622574 -5226 622658
rect -5846 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 -5226 622574
rect -5846 586894 -5226 622338
rect -5846 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 -5226 586894
rect -5846 586574 -5226 586658
rect -5846 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 -5226 586574
rect -5846 550894 -5226 586338
rect -5846 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 -5226 550894
rect -5846 550574 -5226 550658
rect -5846 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 -5226 550574
rect -5846 514894 -5226 550338
rect -5846 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 -5226 514894
rect -5846 514574 -5226 514658
rect -5846 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 -5226 514574
rect -5846 478894 -5226 514338
rect -5846 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 -5226 478894
rect -5846 478574 -5226 478658
rect -5846 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 -5226 478574
rect -5846 442894 -5226 478338
rect -5846 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 -5226 442894
rect -5846 442574 -5226 442658
rect -5846 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 -5226 442574
rect -5846 406894 -5226 442338
rect -5846 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 -5226 406894
rect -5846 406574 -5226 406658
rect -5846 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 -5226 406574
rect -5846 370894 -5226 406338
rect -5846 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 -5226 370894
rect -5846 370574 -5226 370658
rect -5846 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 -5226 370574
rect -5846 334894 -5226 370338
rect -5846 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 -5226 334894
rect -5846 334574 -5226 334658
rect -5846 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 -5226 334574
rect -5846 298894 -5226 334338
rect -5846 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 -5226 298894
rect -5846 298574 -5226 298658
rect -5846 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 -5226 298574
rect -5846 262894 -5226 298338
rect -5846 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 -5226 262894
rect -5846 262574 -5226 262658
rect -5846 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 -5226 262574
rect -5846 226894 -5226 262338
rect -5846 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 -5226 226894
rect -5846 226574 -5226 226658
rect -5846 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 -5226 226574
rect -5846 190894 -5226 226338
rect -5846 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 -5226 190894
rect -5846 190574 -5226 190658
rect -5846 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 -5226 190574
rect -5846 154894 -5226 190338
rect -5846 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 -5226 154894
rect -5846 154574 -5226 154658
rect -5846 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 -5226 154574
rect -5846 118894 -5226 154338
rect -5846 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 -5226 118894
rect -5846 118574 -5226 118658
rect -5846 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 -5226 118574
rect -5846 82894 -5226 118338
rect -5846 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 -5226 82894
rect -5846 82574 -5226 82658
rect -5846 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 -5226 82574
rect -5846 46894 -5226 82338
rect -5846 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 -5226 46894
rect -5846 46574 -5226 46658
rect -5846 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 -5226 46574
rect -5846 10894 -5226 46338
rect -5846 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 -5226 10894
rect -5846 10574 -5226 10658
rect -5846 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 -5226 10574
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 673174 -4266 707162
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 -4266 673174
rect -4886 672854 -4266 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 -4266 672854
rect -4886 637174 -4266 672618
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 -4266 637174
rect -4886 636854 -4266 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 -4266 636854
rect -4886 601174 -4266 636618
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 -4266 601174
rect -4886 600854 -4266 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 -4266 600854
rect -4886 565174 -4266 600618
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 -4266 565174
rect -4886 564854 -4266 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 -4266 564854
rect -4886 529174 -4266 564618
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 -4266 529174
rect -4886 528854 -4266 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 -4266 528854
rect -4886 493174 -4266 528618
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 -4266 493174
rect -4886 492854 -4266 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 -4266 492854
rect -4886 457174 -4266 492618
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 -4266 457174
rect -4886 456854 -4266 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 -4266 456854
rect -4886 421174 -4266 456618
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 -4266 421174
rect -4886 420854 -4266 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 -4266 420854
rect -4886 385174 -4266 420618
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 -4266 385174
rect -4886 384854 -4266 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 -4266 384854
rect -4886 349174 -4266 384618
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 -4266 349174
rect -4886 348854 -4266 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 -4266 348854
rect -4886 313174 -4266 348618
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 -4266 313174
rect -4886 312854 -4266 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 -4266 312854
rect -4886 277174 -4266 312618
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 -4266 277174
rect -4886 276854 -4266 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 -4266 276854
rect -4886 241174 -4266 276618
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 -4266 241174
rect -4886 240854 -4266 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 -4266 240854
rect -4886 205174 -4266 240618
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 -4266 205174
rect -4886 204854 -4266 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 -4266 204854
rect -4886 169174 -4266 204618
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 -4266 169174
rect -4886 168854 -4266 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 -4266 168854
rect -4886 133174 -4266 168618
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 -4266 133174
rect -4886 132854 -4266 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 -4266 132854
rect -4886 97174 -4266 132618
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 -4266 97174
rect -4886 96854 -4266 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 -4266 96854
rect -4886 61174 -4266 96618
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 -4266 61174
rect -4886 60854 -4266 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 -4266 60854
rect -4886 25174 -4266 60618
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 -4266 25174
rect -4886 24854 -4266 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 -4266 24854
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 6134 706758
rect 5514 706438 6134 706522
rect 5514 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 6134 706438
rect -3926 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 -3306 691174
rect -3926 690854 -3306 690938
rect -3926 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 -3306 690854
rect -3926 655174 -3306 690618
rect -3926 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 -3306 655174
rect -3926 654854 -3306 654938
rect -3926 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 -3306 654854
rect -3926 619174 -3306 654618
rect -3926 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 -3306 619174
rect -3926 618854 -3306 618938
rect -3926 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 -3306 618854
rect -3926 583174 -3306 618618
rect -3926 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 -3306 583174
rect -3926 582854 -3306 582938
rect -3926 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 -3306 582854
rect -3926 547174 -3306 582618
rect -3926 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 -3306 547174
rect -3926 546854 -3306 546938
rect -3926 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 -3306 546854
rect -3926 511174 -3306 546618
rect -3926 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 -3306 511174
rect -3926 510854 -3306 510938
rect -3926 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 -3306 510854
rect -3926 475174 -3306 510618
rect -3926 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 -3306 475174
rect -3926 474854 -3306 474938
rect -3926 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 -3306 474854
rect -3926 439174 -3306 474618
rect -3926 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 -3306 439174
rect -3926 438854 -3306 438938
rect -3926 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 -3306 438854
rect -3926 403174 -3306 438618
rect -3926 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 -3306 403174
rect -3926 402854 -3306 402938
rect -3926 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 -3306 402854
rect -3926 367174 -3306 402618
rect -3926 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 -3306 367174
rect -3926 366854 -3306 366938
rect -3926 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 -3306 366854
rect -3926 331174 -3306 366618
rect -3926 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 -3306 331174
rect -3926 330854 -3306 330938
rect -3926 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 -3306 330854
rect -3926 295174 -3306 330618
rect -3926 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 -3306 295174
rect -3926 294854 -3306 294938
rect -3926 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 -3306 294854
rect -3926 259174 -3306 294618
rect -3926 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 -3306 259174
rect -3926 258854 -3306 258938
rect -3926 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 -3306 258854
rect -3926 223174 -3306 258618
rect -3926 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 -3306 223174
rect -3926 222854 -3306 222938
rect -3926 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 -3306 222854
rect -3926 187174 -3306 222618
rect -3926 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 -3306 187174
rect -3926 186854 -3306 186938
rect -3926 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 -3306 186854
rect -3926 151174 -3306 186618
rect -3926 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 -3306 151174
rect -3926 150854 -3306 150938
rect -3926 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 -3306 150854
rect -3926 115174 -3306 150618
rect -3926 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 -3306 115174
rect -3926 114854 -3306 114938
rect -3926 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 -3306 114854
rect -3926 79174 -3306 114618
rect -3926 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 -3306 79174
rect -3926 78854 -3306 78938
rect -3926 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 -3306 78854
rect -3926 43174 -3306 78618
rect -3926 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 -3306 43174
rect -3926 42854 -3306 42938
rect -3926 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 -3306 42854
rect -3926 7174 -3306 42618
rect -3926 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 -3306 7174
rect -3926 6854 -3306 6938
rect -3926 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 -3306 6854
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 702000 2414 704282
rect 5514 702000 6134 706202
rect 9234 702000 9854 708122
rect 12954 702000 13574 710042
rect 30954 711558 31574 711590
rect 30954 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 31574 711558
rect 30954 711238 31574 711322
rect 30954 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 31574 711238
rect 27234 709638 27854 709670
rect 27234 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 27854 709638
rect 27234 709318 27854 709402
rect 27234 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 27854 709318
rect 23514 707718 24134 707750
rect 23514 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 24134 707718
rect 23514 707398 24134 707482
rect 23514 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 24134 707398
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 19794 702000 20414 705242
rect 23514 702000 24134 707162
rect 27234 702000 27854 709082
rect 30954 702000 31574 711002
rect 48954 710598 49574 711590
rect 48954 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 49574 710598
rect 48954 710278 49574 710362
rect 48954 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 49574 710278
rect 45234 708678 45854 709670
rect 45234 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 45854 708678
rect 45234 708358 45854 708442
rect 45234 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 45854 708358
rect 41514 706758 42134 707750
rect 41514 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 42134 706758
rect 41514 706438 42134 706522
rect 41514 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 42134 706438
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 702000 38414 704282
rect 41514 702000 42134 706202
rect 45234 702000 45854 708122
rect 48954 702000 49574 710042
rect 66954 711558 67574 711590
rect 66954 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 67574 711558
rect 66954 711238 67574 711322
rect 66954 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 67574 711238
rect 63234 709638 63854 709670
rect 63234 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 63854 709638
rect 63234 709318 63854 709402
rect 63234 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 63854 709318
rect 59514 707718 60134 707750
rect 59514 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 60134 707718
rect 59514 707398 60134 707482
rect 59514 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 60134 707398
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 702000 56414 705242
rect 59514 702000 60134 707162
rect 63234 702000 63854 709082
rect 66954 702000 67574 711002
rect 84954 710598 85574 711590
rect 84954 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 85574 710598
rect 84954 710278 85574 710362
rect 84954 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 85574 710278
rect 81234 708678 81854 709670
rect 81234 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 81854 708678
rect 81234 708358 81854 708442
rect 81234 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 81854 708358
rect 77514 706758 78134 707750
rect 77514 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 78134 706758
rect 77514 706438 78134 706522
rect 77514 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 78134 706438
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 702000 74414 704282
rect 77514 702000 78134 706202
rect 81234 702000 81854 708122
rect 84954 702000 85574 710042
rect 102954 711558 103574 711590
rect 102954 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 103574 711558
rect 102954 711238 103574 711322
rect 102954 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 103574 711238
rect 99234 709638 99854 709670
rect 99234 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 99854 709638
rect 99234 709318 99854 709402
rect 99234 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 99854 709318
rect 95514 707718 96134 707750
rect 95514 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 96134 707718
rect 95514 707398 96134 707482
rect 95514 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 96134 707398
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 702000 92414 705242
rect 95514 702000 96134 707162
rect 99234 702000 99854 709082
rect 102954 702000 103574 711002
rect 120954 710598 121574 711590
rect 120954 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 121574 710598
rect 120954 710278 121574 710362
rect 120954 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 121574 710278
rect 117234 708678 117854 709670
rect 117234 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 117854 708678
rect 117234 708358 117854 708442
rect 117234 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 117854 708358
rect 113514 706758 114134 707750
rect 113514 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 114134 706758
rect 113514 706438 114134 706522
rect 113514 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 114134 706438
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 702000 110414 704282
rect 113514 702000 114134 706202
rect 117234 702000 117854 708122
rect 120954 702000 121574 710042
rect 138954 711558 139574 711590
rect 138954 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 139574 711558
rect 138954 711238 139574 711322
rect 138954 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 139574 711238
rect 135234 709638 135854 709670
rect 135234 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 135854 709638
rect 135234 709318 135854 709402
rect 135234 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 135854 709318
rect 131514 707718 132134 707750
rect 131514 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 132134 707718
rect 131514 707398 132134 707482
rect 131514 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 132134 707398
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 127794 702000 128414 705242
rect 131514 702000 132134 707162
rect 135234 702000 135854 709082
rect 138954 702000 139574 711002
rect 156954 710598 157574 711590
rect 156954 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 157574 710598
rect 156954 710278 157574 710362
rect 156954 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 157574 710278
rect 153234 708678 153854 709670
rect 153234 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 153854 708678
rect 153234 708358 153854 708442
rect 153234 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 153854 708358
rect 149514 706758 150134 707750
rect 149514 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 150134 706758
rect 149514 706438 150134 706522
rect 149514 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 150134 706438
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 702000 146414 704282
rect 149514 702000 150134 706202
rect 153234 702000 153854 708122
rect 156954 702000 157574 710042
rect 174954 711558 175574 711590
rect 174954 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 175574 711558
rect 174954 711238 175574 711322
rect 174954 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 175574 711238
rect 171234 709638 171854 709670
rect 171234 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 171854 709638
rect 171234 709318 171854 709402
rect 171234 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 171854 709318
rect 167514 707718 168134 707750
rect 167514 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 168134 707718
rect 167514 707398 168134 707482
rect 167514 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 168134 707398
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 702000 164414 705242
rect 167514 702000 168134 707162
rect 171234 702000 171854 709082
rect 174954 702000 175574 711002
rect 192954 710598 193574 711590
rect 192954 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 193574 710598
rect 192954 710278 193574 710362
rect 192954 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 193574 710278
rect 189234 708678 189854 709670
rect 189234 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 189854 708678
rect 189234 708358 189854 708442
rect 189234 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 189854 708358
rect 185514 706758 186134 707750
rect 185514 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 186134 706758
rect 185514 706438 186134 706522
rect 185514 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 186134 706438
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 702000 182414 704282
rect 185514 702000 186134 706202
rect 189234 702000 189854 708122
rect 192954 702000 193574 710042
rect 210954 711558 211574 711590
rect 210954 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 211574 711558
rect 210954 711238 211574 711322
rect 210954 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 211574 711238
rect 207234 709638 207854 709670
rect 207234 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 207854 709638
rect 207234 709318 207854 709402
rect 207234 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 207854 709318
rect 203514 707718 204134 707750
rect 203514 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 204134 707718
rect 203514 707398 204134 707482
rect 203514 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 204134 707398
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 702000 200414 705242
rect 203514 702000 204134 707162
rect 207234 702000 207854 709082
rect 210954 702000 211574 711002
rect 228954 710598 229574 711590
rect 228954 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 229574 710598
rect 228954 710278 229574 710362
rect 228954 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 229574 710278
rect 225234 708678 225854 709670
rect 225234 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 225854 708678
rect 225234 708358 225854 708442
rect 225234 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 225854 708358
rect 221514 706758 222134 707750
rect 221514 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 222134 706758
rect 221514 706438 222134 706522
rect 221514 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 222134 706438
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 702000 218414 704282
rect 221514 702000 222134 706202
rect 225234 702000 225854 708122
rect 228954 702000 229574 710042
rect 246954 711558 247574 711590
rect 246954 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 247574 711558
rect 246954 711238 247574 711322
rect 246954 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 247574 711238
rect 243234 709638 243854 709670
rect 243234 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 243854 709638
rect 243234 709318 243854 709402
rect 243234 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 243854 709318
rect 239514 707718 240134 707750
rect 239514 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 240134 707718
rect 239514 707398 240134 707482
rect 239514 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 240134 707398
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 235794 702000 236414 705242
rect 239514 702000 240134 707162
rect 243234 702000 243854 709082
rect 246954 702000 247574 711002
rect 264954 710598 265574 711590
rect 264954 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 265574 710598
rect 264954 710278 265574 710362
rect 264954 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 265574 710278
rect 261234 708678 261854 709670
rect 261234 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 261854 708678
rect 261234 708358 261854 708442
rect 261234 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 261854 708358
rect 257514 706758 258134 707750
rect 257514 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 258134 706758
rect 257514 706438 258134 706522
rect 257514 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 258134 706438
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 702000 254414 704282
rect 257514 702000 258134 706202
rect 261234 702000 261854 708122
rect 264954 702000 265574 710042
rect 282954 711558 283574 711590
rect 282954 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 283574 711558
rect 282954 711238 283574 711322
rect 282954 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 283574 711238
rect 279234 709638 279854 709670
rect 279234 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 279854 709638
rect 279234 709318 279854 709402
rect 279234 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 279854 709318
rect 275514 707718 276134 707750
rect 275514 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 276134 707718
rect 275514 707398 276134 707482
rect 275514 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 276134 707398
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 271794 702000 272414 705242
rect 275514 702000 276134 707162
rect 279234 702000 279854 709082
rect 282954 702000 283574 711002
rect 300954 710598 301574 711590
rect 300954 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 301574 710598
rect 300954 710278 301574 710362
rect 300954 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 301574 710278
rect 297234 708678 297854 709670
rect 297234 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 297854 708678
rect 297234 708358 297854 708442
rect 297234 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 297854 708358
rect 293514 706758 294134 707750
rect 293514 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 294134 706758
rect 293514 706438 294134 706522
rect 293514 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 294134 706438
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 702000 290414 704282
rect 293514 702000 294134 706202
rect 297234 702000 297854 708122
rect 300954 702000 301574 710042
rect 318954 711558 319574 711590
rect 318954 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 319574 711558
rect 318954 711238 319574 711322
rect 318954 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 319574 711238
rect 315234 709638 315854 709670
rect 315234 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 315854 709638
rect 315234 709318 315854 709402
rect 315234 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 315854 709318
rect 311514 707718 312134 707750
rect 311514 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 312134 707718
rect 311514 707398 312134 707482
rect 311514 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 312134 707398
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 702000 308414 705242
rect 311514 702000 312134 707162
rect 315234 702000 315854 709082
rect 318954 702000 319574 711002
rect 336954 710598 337574 711590
rect 336954 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 337574 710598
rect 336954 710278 337574 710362
rect 336954 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 337574 710278
rect 333234 708678 333854 709670
rect 333234 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 333854 708678
rect 333234 708358 333854 708442
rect 333234 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 333854 708358
rect 329514 706758 330134 707750
rect 329514 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 330134 706758
rect 329514 706438 330134 706522
rect 329514 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 330134 706438
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 702000 326414 704282
rect 329514 702000 330134 706202
rect 333234 702000 333854 708122
rect 336954 702000 337574 710042
rect 354954 711558 355574 711590
rect 354954 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 355574 711558
rect 354954 711238 355574 711322
rect 354954 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 355574 711238
rect 351234 709638 351854 709670
rect 351234 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 351854 709638
rect 351234 709318 351854 709402
rect 351234 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 351854 709318
rect 347514 707718 348134 707750
rect 347514 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 348134 707718
rect 347514 707398 348134 707482
rect 347514 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 348134 707398
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 343794 702000 344414 705242
rect 347514 702000 348134 707162
rect 351234 702000 351854 709082
rect 354954 702000 355574 711002
rect 372954 710598 373574 711590
rect 372954 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 373574 710598
rect 372954 710278 373574 710362
rect 372954 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 373574 710278
rect 369234 708678 369854 709670
rect 369234 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 369854 708678
rect 369234 708358 369854 708442
rect 369234 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 369854 708358
rect 365514 706758 366134 707750
rect 365514 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 366134 706758
rect 365514 706438 366134 706522
rect 365514 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 366134 706438
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 702000 362414 704282
rect 365514 702000 366134 706202
rect 369234 702000 369854 708122
rect 372954 702000 373574 710042
rect 390954 711558 391574 711590
rect 390954 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 391574 711558
rect 390954 711238 391574 711322
rect 390954 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 391574 711238
rect 387234 709638 387854 709670
rect 387234 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 387854 709638
rect 387234 709318 387854 709402
rect 387234 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 387854 709318
rect 383514 707718 384134 707750
rect 383514 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 384134 707718
rect 383514 707398 384134 707482
rect 383514 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 384134 707398
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 379794 702000 380414 705242
rect 383514 702000 384134 707162
rect 387234 702000 387854 709082
rect 390954 702000 391574 711002
rect 408954 710598 409574 711590
rect 408954 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 409574 710598
rect 408954 710278 409574 710362
rect 408954 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 409574 710278
rect 405234 708678 405854 709670
rect 405234 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 405854 708678
rect 405234 708358 405854 708442
rect 405234 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 405854 708358
rect 401514 706758 402134 707750
rect 401514 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 402134 706758
rect 401514 706438 402134 706522
rect 401514 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 402134 706438
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 702000 398414 704282
rect 401514 702000 402134 706202
rect 405234 702000 405854 708122
rect 408954 702000 409574 710042
rect 426954 711558 427574 711590
rect 426954 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 427574 711558
rect 426954 711238 427574 711322
rect 426954 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 427574 711238
rect 423234 709638 423854 709670
rect 423234 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 423854 709638
rect 423234 709318 423854 709402
rect 423234 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 423854 709318
rect 419514 707718 420134 707750
rect 419514 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 420134 707718
rect 419514 707398 420134 707482
rect 419514 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 420134 707398
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 415794 702000 416414 705242
rect 419514 702000 420134 707162
rect 423234 702000 423854 709082
rect 426954 702000 427574 711002
rect 444954 710598 445574 711590
rect 444954 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 445574 710598
rect 444954 710278 445574 710362
rect 444954 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 445574 710278
rect 441234 708678 441854 709670
rect 441234 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 441854 708678
rect 441234 708358 441854 708442
rect 441234 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 441854 708358
rect 437514 706758 438134 707750
rect 437514 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 438134 706758
rect 437514 706438 438134 706522
rect 437514 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 438134 706438
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 702000 434414 704282
rect 437514 702000 438134 706202
rect 441234 702000 441854 708122
rect 444954 702000 445574 710042
rect 462954 711558 463574 711590
rect 462954 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 463574 711558
rect 462954 711238 463574 711322
rect 462954 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 463574 711238
rect 459234 709638 459854 709670
rect 459234 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 459854 709638
rect 459234 709318 459854 709402
rect 459234 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 459854 709318
rect 455514 707718 456134 707750
rect 455514 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 456134 707718
rect 455514 707398 456134 707482
rect 455514 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 456134 707398
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 702000 452414 705242
rect 455514 702000 456134 707162
rect 459234 702000 459854 709082
rect 462954 702000 463574 711002
rect 480954 710598 481574 711590
rect 480954 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 481574 710598
rect 480954 710278 481574 710362
rect 480954 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 481574 710278
rect 477234 708678 477854 709670
rect 477234 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 477854 708678
rect 477234 708358 477854 708442
rect 477234 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 477854 708358
rect 473514 706758 474134 707750
rect 473514 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 474134 706758
rect 473514 706438 474134 706522
rect 473514 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 474134 706438
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 702000 470414 704282
rect 473514 702000 474134 706202
rect 477234 702000 477854 708122
rect 480954 702000 481574 710042
rect 498954 711558 499574 711590
rect 498954 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 499574 711558
rect 498954 711238 499574 711322
rect 498954 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 499574 711238
rect 495234 709638 495854 709670
rect 495234 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 495854 709638
rect 495234 709318 495854 709402
rect 495234 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 495854 709318
rect 491514 707718 492134 707750
rect 491514 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 492134 707718
rect 491514 707398 492134 707482
rect 491514 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 492134 707398
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 487794 702000 488414 705242
rect 491514 702000 492134 707162
rect 495234 702000 495854 709082
rect 498954 702000 499574 711002
rect 516954 710598 517574 711590
rect 516954 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 517574 710598
rect 516954 710278 517574 710362
rect 516954 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 517574 710278
rect 513234 708678 513854 709670
rect 513234 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 513854 708678
rect 513234 708358 513854 708442
rect 513234 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 513854 708358
rect 509514 706758 510134 707750
rect 509514 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 510134 706758
rect 509514 706438 510134 706522
rect 509514 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 510134 706438
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 702000 506414 704282
rect 509514 702000 510134 706202
rect 513234 702000 513854 708122
rect 516954 702000 517574 710042
rect 534954 711558 535574 711590
rect 534954 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 535574 711558
rect 534954 711238 535574 711322
rect 534954 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 535574 711238
rect 531234 709638 531854 709670
rect 531234 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 531854 709638
rect 531234 709318 531854 709402
rect 531234 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 531854 709318
rect 527514 707718 528134 707750
rect 527514 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 528134 707718
rect 527514 707398 528134 707482
rect 527514 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 528134 707398
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 702000 524414 705242
rect 527514 702000 528134 707162
rect 531234 702000 531854 709082
rect 534954 702000 535574 711002
rect 552954 710598 553574 711590
rect 552954 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 553574 710598
rect 552954 710278 553574 710362
rect 552954 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 553574 710278
rect 549234 708678 549854 709670
rect 549234 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 549854 708678
rect 549234 708358 549854 708442
rect 549234 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 549854 708358
rect 545514 706758 546134 707750
rect 545514 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 546134 706758
rect 545514 706438 546134 706522
rect 545514 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 546134 706438
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 702000 542414 704282
rect 545514 702000 546134 706202
rect 549234 702000 549854 708122
rect 552954 702000 553574 710042
rect 570954 711558 571574 711590
rect 570954 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 571574 711558
rect 570954 711238 571574 711322
rect 570954 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 571574 711238
rect 567234 709638 567854 709670
rect 567234 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 567854 709638
rect 567234 709318 567854 709402
rect 567234 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 567854 709318
rect 563514 707718 564134 707750
rect 563514 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 564134 707718
rect 563514 707398 564134 707482
rect 563514 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 564134 707398
rect 559794 705798 560414 705830
rect 559794 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 560414 705798
rect 559794 705478 560414 705562
rect 559794 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 560414 705478
rect 559794 702000 560414 705242
rect 563514 702000 564134 707162
rect 164187 701180 164253 701181
rect 164187 701116 164188 701180
rect 164252 701116 164253 701180
rect 164187 701115 164253 701116
rect 11467 699412 11533 699413
rect 11467 699348 11468 699412
rect 11532 699348 11533 699412
rect 11467 699347 11533 699348
rect 13859 699412 13925 699413
rect 13859 699348 13860 699412
rect 13924 699348 13925 699412
rect 13859 699347 13925 699348
rect 21403 699412 21469 699413
rect 21403 699348 21404 699412
rect 21468 699348 21469 699412
rect 21403 699347 21469 699348
rect 30971 699412 31037 699413
rect 30971 699348 30972 699412
rect 31036 699348 31037 699412
rect 30971 699347 31037 699348
rect 33363 699412 33429 699413
rect 33363 699348 33364 699412
rect 33428 699348 33429 699412
rect 33363 699347 33429 699348
rect 43115 699412 43181 699413
rect 43115 699348 43116 699412
rect 43180 699348 43181 699412
rect 43115 699347 43181 699348
rect 11470 698325 11530 699347
rect 13862 698461 13922 699347
rect 21406 698597 21466 699347
rect 30974 698733 31034 699347
rect 33366 698869 33426 699347
rect 43118 699005 43178 699347
rect 164190 699277 164250 701115
rect 433379 699548 433445 699549
rect 433379 699484 433380 699548
rect 433444 699484 433445 699548
rect 433379 699483 433445 699484
rect 408907 699412 408973 699413
rect 408907 699348 408908 699412
rect 408972 699348 408973 699412
rect 408907 699347 408973 699348
rect 418659 699412 418725 699413
rect 418659 699348 418660 699412
rect 418724 699348 418725 699412
rect 418659 699347 418725 699348
rect 164187 699276 164253 699277
rect 164187 699212 164188 699276
rect 164252 699212 164253 699276
rect 164187 699211 164253 699212
rect 43115 699004 43181 699005
rect 43115 698940 43116 699004
rect 43180 698940 43181 699004
rect 43115 698939 43181 698940
rect 33363 698868 33429 698869
rect 33363 698804 33364 698868
rect 33428 698804 33429 698868
rect 33363 698803 33429 698804
rect 30971 698732 31037 698733
rect 30971 698668 30972 698732
rect 31036 698668 31037 698732
rect 30971 698667 31037 698668
rect 21403 698596 21469 698597
rect 21403 698532 21404 698596
rect 21468 698532 21469 698596
rect 21403 698531 21469 698532
rect 13859 698460 13925 698461
rect 13859 698396 13860 698460
rect 13924 698396 13925 698460
rect 13859 698395 13925 698396
rect 11467 698324 11533 698325
rect 11467 698260 11468 698324
rect 11532 698260 11533 698324
rect 11467 698259 11533 698260
rect 408910 698053 408970 699347
rect 409091 699276 409157 699277
rect 409091 699212 409092 699276
rect 409156 699212 409157 699276
rect 409091 699211 409157 699212
rect 409094 698053 409154 699211
rect 418662 698189 418722 699347
rect 418659 698188 418725 698189
rect 418659 698124 418660 698188
rect 418724 698124 418725 698188
rect 418659 698123 418725 698124
rect 408907 698052 408973 698053
rect 408907 697988 408908 698052
rect 408972 697988 408973 698052
rect 408907 697987 408973 697988
rect 409091 698052 409157 698053
rect 409091 697988 409092 698052
rect 409156 697988 409157 698052
rect 409091 697987 409157 697988
rect 433382 697917 433442 699483
rect 448099 699412 448165 699413
rect 448099 699348 448100 699412
rect 448164 699348 448165 699412
rect 448099 699347 448165 699348
rect 453067 699412 453133 699413
rect 453067 699348 453068 699412
rect 453132 699348 453133 699412
rect 453067 699347 453133 699348
rect 433379 697916 433445 697917
rect 433379 697852 433380 697916
rect 433444 697852 433445 697916
rect 433379 697851 433445 697852
rect 448102 697781 448162 699347
rect 448099 697780 448165 697781
rect 448099 697716 448100 697780
rect 448164 697716 448165 697780
rect 448099 697715 448165 697716
rect 453070 697645 453130 699347
rect 453067 697644 453133 697645
rect 453067 697580 453068 697644
rect 453132 697580 453133 697644
rect 453067 697579 453133 697580
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect 8208 687454 8528 687486
rect 8208 687218 8250 687454
rect 8486 687218 8528 687454
rect 8208 687134 8528 687218
rect 8208 686898 8250 687134
rect 8486 686898 8528 687134
rect 8208 686866 8528 686898
rect 38928 687454 39248 687486
rect 38928 687218 38970 687454
rect 39206 687218 39248 687454
rect 38928 687134 39248 687218
rect 38928 686898 38970 687134
rect 39206 686898 39248 687134
rect 38928 686866 39248 686898
rect 69648 687454 69968 687486
rect 69648 687218 69690 687454
rect 69926 687218 69968 687454
rect 69648 687134 69968 687218
rect 69648 686898 69690 687134
rect 69926 686898 69968 687134
rect 69648 686866 69968 686898
rect 100368 687454 100688 687486
rect 100368 687218 100410 687454
rect 100646 687218 100688 687454
rect 100368 687134 100688 687218
rect 100368 686898 100410 687134
rect 100646 686898 100688 687134
rect 100368 686866 100688 686898
rect 131088 687454 131408 687486
rect 131088 687218 131130 687454
rect 131366 687218 131408 687454
rect 131088 687134 131408 687218
rect 131088 686898 131130 687134
rect 131366 686898 131408 687134
rect 131088 686866 131408 686898
rect 161808 687454 162128 687486
rect 161808 687218 161850 687454
rect 162086 687218 162128 687454
rect 161808 687134 162128 687218
rect 161808 686898 161850 687134
rect 162086 686898 162128 687134
rect 161808 686866 162128 686898
rect 192528 687454 192848 687486
rect 192528 687218 192570 687454
rect 192806 687218 192848 687454
rect 192528 687134 192848 687218
rect 192528 686898 192570 687134
rect 192806 686898 192848 687134
rect 192528 686866 192848 686898
rect 223248 687454 223568 687486
rect 223248 687218 223290 687454
rect 223526 687218 223568 687454
rect 223248 687134 223568 687218
rect 223248 686898 223290 687134
rect 223526 686898 223568 687134
rect 223248 686866 223568 686898
rect 253968 687454 254288 687486
rect 253968 687218 254010 687454
rect 254246 687218 254288 687454
rect 253968 687134 254288 687218
rect 253968 686898 254010 687134
rect 254246 686898 254288 687134
rect 253968 686866 254288 686898
rect 284688 687454 285008 687486
rect 284688 687218 284730 687454
rect 284966 687218 285008 687454
rect 284688 687134 285008 687218
rect 284688 686898 284730 687134
rect 284966 686898 285008 687134
rect 284688 686866 285008 686898
rect 315408 687454 315728 687486
rect 315408 687218 315450 687454
rect 315686 687218 315728 687454
rect 315408 687134 315728 687218
rect 315408 686898 315450 687134
rect 315686 686898 315728 687134
rect 315408 686866 315728 686898
rect 346128 687454 346448 687486
rect 346128 687218 346170 687454
rect 346406 687218 346448 687454
rect 346128 687134 346448 687218
rect 346128 686898 346170 687134
rect 346406 686898 346448 687134
rect 346128 686866 346448 686898
rect 376848 687454 377168 687486
rect 376848 687218 376890 687454
rect 377126 687218 377168 687454
rect 376848 687134 377168 687218
rect 376848 686898 376890 687134
rect 377126 686898 377168 687134
rect 376848 686866 377168 686898
rect 407568 687454 407888 687486
rect 407568 687218 407610 687454
rect 407846 687218 407888 687454
rect 407568 687134 407888 687218
rect 407568 686898 407610 687134
rect 407846 686898 407888 687134
rect 407568 686866 407888 686898
rect 438288 687454 438608 687486
rect 438288 687218 438330 687454
rect 438566 687218 438608 687454
rect 438288 687134 438608 687218
rect 438288 686898 438330 687134
rect 438566 686898 438608 687134
rect 438288 686866 438608 686898
rect 469008 687454 469328 687486
rect 469008 687218 469050 687454
rect 469286 687218 469328 687454
rect 469008 687134 469328 687218
rect 469008 686898 469050 687134
rect 469286 686898 469328 687134
rect 469008 686866 469328 686898
rect 499728 687454 500048 687486
rect 499728 687218 499770 687454
rect 500006 687218 500048 687454
rect 499728 687134 500048 687218
rect 499728 686898 499770 687134
rect 500006 686898 500048 687134
rect 499728 686866 500048 686898
rect 530448 687454 530768 687486
rect 530448 687218 530490 687454
rect 530726 687218 530768 687454
rect 530448 687134 530768 687218
rect 530448 686898 530490 687134
rect 530726 686898 530768 687134
rect 530448 686866 530768 686898
rect 561168 687454 561488 687486
rect 561168 687218 561210 687454
rect 561446 687218 561488 687454
rect 561168 687134 561488 687218
rect 561168 686898 561210 687134
rect 561446 686898 561488 687134
rect 561168 686866 561488 686898
rect 567234 676894 567854 709082
rect 567234 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 567854 676894
rect 567234 676574 567854 676658
rect 567234 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 567854 676574
rect 23568 669454 23888 669486
rect 23568 669218 23610 669454
rect 23846 669218 23888 669454
rect 23568 669134 23888 669218
rect 23568 668898 23610 669134
rect 23846 668898 23888 669134
rect 23568 668866 23888 668898
rect 54288 669454 54608 669486
rect 54288 669218 54330 669454
rect 54566 669218 54608 669454
rect 54288 669134 54608 669218
rect 54288 668898 54330 669134
rect 54566 668898 54608 669134
rect 54288 668866 54608 668898
rect 85008 669454 85328 669486
rect 85008 669218 85050 669454
rect 85286 669218 85328 669454
rect 85008 669134 85328 669218
rect 85008 668898 85050 669134
rect 85286 668898 85328 669134
rect 85008 668866 85328 668898
rect 115728 669454 116048 669486
rect 115728 669218 115770 669454
rect 116006 669218 116048 669454
rect 115728 669134 116048 669218
rect 115728 668898 115770 669134
rect 116006 668898 116048 669134
rect 115728 668866 116048 668898
rect 146448 669454 146768 669486
rect 146448 669218 146490 669454
rect 146726 669218 146768 669454
rect 146448 669134 146768 669218
rect 146448 668898 146490 669134
rect 146726 668898 146768 669134
rect 146448 668866 146768 668898
rect 177168 669454 177488 669486
rect 177168 669218 177210 669454
rect 177446 669218 177488 669454
rect 177168 669134 177488 669218
rect 177168 668898 177210 669134
rect 177446 668898 177488 669134
rect 177168 668866 177488 668898
rect 207888 669454 208208 669486
rect 207888 669218 207930 669454
rect 208166 669218 208208 669454
rect 207888 669134 208208 669218
rect 207888 668898 207930 669134
rect 208166 668898 208208 669134
rect 207888 668866 208208 668898
rect 238608 669454 238928 669486
rect 238608 669218 238650 669454
rect 238886 669218 238928 669454
rect 238608 669134 238928 669218
rect 238608 668898 238650 669134
rect 238886 668898 238928 669134
rect 238608 668866 238928 668898
rect 269328 669454 269648 669486
rect 269328 669218 269370 669454
rect 269606 669218 269648 669454
rect 269328 669134 269648 669218
rect 269328 668898 269370 669134
rect 269606 668898 269648 669134
rect 269328 668866 269648 668898
rect 300048 669454 300368 669486
rect 300048 669218 300090 669454
rect 300326 669218 300368 669454
rect 300048 669134 300368 669218
rect 300048 668898 300090 669134
rect 300326 668898 300368 669134
rect 300048 668866 300368 668898
rect 330768 669454 331088 669486
rect 330768 669218 330810 669454
rect 331046 669218 331088 669454
rect 330768 669134 331088 669218
rect 330768 668898 330810 669134
rect 331046 668898 331088 669134
rect 330768 668866 331088 668898
rect 361488 669454 361808 669486
rect 361488 669218 361530 669454
rect 361766 669218 361808 669454
rect 361488 669134 361808 669218
rect 361488 668898 361530 669134
rect 361766 668898 361808 669134
rect 361488 668866 361808 668898
rect 392208 669454 392528 669486
rect 392208 669218 392250 669454
rect 392486 669218 392528 669454
rect 392208 669134 392528 669218
rect 392208 668898 392250 669134
rect 392486 668898 392528 669134
rect 392208 668866 392528 668898
rect 422928 669454 423248 669486
rect 422928 669218 422970 669454
rect 423206 669218 423248 669454
rect 422928 669134 423248 669218
rect 422928 668898 422970 669134
rect 423206 668898 423248 669134
rect 422928 668866 423248 668898
rect 453648 669454 453968 669486
rect 453648 669218 453690 669454
rect 453926 669218 453968 669454
rect 453648 669134 453968 669218
rect 453648 668898 453690 669134
rect 453926 668898 453968 669134
rect 453648 668866 453968 668898
rect 484368 669454 484688 669486
rect 484368 669218 484410 669454
rect 484646 669218 484688 669454
rect 484368 669134 484688 669218
rect 484368 668898 484410 669134
rect 484646 668898 484688 669134
rect 484368 668866 484688 668898
rect 515088 669454 515408 669486
rect 515088 669218 515130 669454
rect 515366 669218 515408 669454
rect 515088 669134 515408 669218
rect 515088 668898 515130 669134
rect 515366 668898 515408 669134
rect 515088 668866 515408 668898
rect 545808 669454 546128 669486
rect 545808 669218 545850 669454
rect 546086 669218 546128 669454
rect 545808 669134 546128 669218
rect 545808 668898 545850 669134
rect 546086 668898 546128 669134
rect 545808 668866 546128 668898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect 8208 651454 8528 651486
rect 8208 651218 8250 651454
rect 8486 651218 8528 651454
rect 8208 651134 8528 651218
rect 8208 650898 8250 651134
rect 8486 650898 8528 651134
rect 8208 650866 8528 650898
rect 38928 651454 39248 651486
rect 38928 651218 38970 651454
rect 39206 651218 39248 651454
rect 38928 651134 39248 651218
rect 38928 650898 38970 651134
rect 39206 650898 39248 651134
rect 38928 650866 39248 650898
rect 69648 651454 69968 651486
rect 69648 651218 69690 651454
rect 69926 651218 69968 651454
rect 69648 651134 69968 651218
rect 69648 650898 69690 651134
rect 69926 650898 69968 651134
rect 69648 650866 69968 650898
rect 100368 651454 100688 651486
rect 100368 651218 100410 651454
rect 100646 651218 100688 651454
rect 100368 651134 100688 651218
rect 100368 650898 100410 651134
rect 100646 650898 100688 651134
rect 100368 650866 100688 650898
rect 131088 651454 131408 651486
rect 131088 651218 131130 651454
rect 131366 651218 131408 651454
rect 131088 651134 131408 651218
rect 131088 650898 131130 651134
rect 131366 650898 131408 651134
rect 131088 650866 131408 650898
rect 161808 651454 162128 651486
rect 161808 651218 161850 651454
rect 162086 651218 162128 651454
rect 161808 651134 162128 651218
rect 161808 650898 161850 651134
rect 162086 650898 162128 651134
rect 161808 650866 162128 650898
rect 192528 651454 192848 651486
rect 192528 651218 192570 651454
rect 192806 651218 192848 651454
rect 192528 651134 192848 651218
rect 192528 650898 192570 651134
rect 192806 650898 192848 651134
rect 192528 650866 192848 650898
rect 223248 651454 223568 651486
rect 223248 651218 223290 651454
rect 223526 651218 223568 651454
rect 223248 651134 223568 651218
rect 223248 650898 223290 651134
rect 223526 650898 223568 651134
rect 223248 650866 223568 650898
rect 253968 651454 254288 651486
rect 253968 651218 254010 651454
rect 254246 651218 254288 651454
rect 253968 651134 254288 651218
rect 253968 650898 254010 651134
rect 254246 650898 254288 651134
rect 253968 650866 254288 650898
rect 284688 651454 285008 651486
rect 284688 651218 284730 651454
rect 284966 651218 285008 651454
rect 284688 651134 285008 651218
rect 284688 650898 284730 651134
rect 284966 650898 285008 651134
rect 284688 650866 285008 650898
rect 315408 651454 315728 651486
rect 315408 651218 315450 651454
rect 315686 651218 315728 651454
rect 315408 651134 315728 651218
rect 315408 650898 315450 651134
rect 315686 650898 315728 651134
rect 315408 650866 315728 650898
rect 346128 651454 346448 651486
rect 346128 651218 346170 651454
rect 346406 651218 346448 651454
rect 346128 651134 346448 651218
rect 346128 650898 346170 651134
rect 346406 650898 346448 651134
rect 346128 650866 346448 650898
rect 376848 651454 377168 651486
rect 376848 651218 376890 651454
rect 377126 651218 377168 651454
rect 376848 651134 377168 651218
rect 376848 650898 376890 651134
rect 377126 650898 377168 651134
rect 376848 650866 377168 650898
rect 407568 651454 407888 651486
rect 407568 651218 407610 651454
rect 407846 651218 407888 651454
rect 407568 651134 407888 651218
rect 407568 650898 407610 651134
rect 407846 650898 407888 651134
rect 407568 650866 407888 650898
rect 438288 651454 438608 651486
rect 438288 651218 438330 651454
rect 438566 651218 438608 651454
rect 438288 651134 438608 651218
rect 438288 650898 438330 651134
rect 438566 650898 438608 651134
rect 438288 650866 438608 650898
rect 469008 651454 469328 651486
rect 469008 651218 469050 651454
rect 469286 651218 469328 651454
rect 469008 651134 469328 651218
rect 469008 650898 469050 651134
rect 469286 650898 469328 651134
rect 469008 650866 469328 650898
rect 499728 651454 500048 651486
rect 499728 651218 499770 651454
rect 500006 651218 500048 651454
rect 499728 651134 500048 651218
rect 499728 650898 499770 651134
rect 500006 650898 500048 651134
rect 499728 650866 500048 650898
rect 530448 651454 530768 651486
rect 530448 651218 530490 651454
rect 530726 651218 530768 651454
rect 530448 651134 530768 651218
rect 530448 650898 530490 651134
rect 530726 650898 530768 651134
rect 530448 650866 530768 650898
rect 561168 651454 561488 651486
rect 561168 651218 561210 651454
rect 561446 651218 561488 651454
rect 561168 651134 561488 651218
rect 561168 650898 561210 651134
rect 561446 650898 561488 651134
rect 561168 650866 561488 650898
rect 567234 640894 567854 676338
rect 567234 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 567854 640894
rect 567234 640574 567854 640658
rect 567234 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 567854 640574
rect 23568 633454 23888 633486
rect 23568 633218 23610 633454
rect 23846 633218 23888 633454
rect 23568 633134 23888 633218
rect 23568 632898 23610 633134
rect 23846 632898 23888 633134
rect 23568 632866 23888 632898
rect 54288 633454 54608 633486
rect 54288 633218 54330 633454
rect 54566 633218 54608 633454
rect 54288 633134 54608 633218
rect 54288 632898 54330 633134
rect 54566 632898 54608 633134
rect 54288 632866 54608 632898
rect 85008 633454 85328 633486
rect 85008 633218 85050 633454
rect 85286 633218 85328 633454
rect 85008 633134 85328 633218
rect 85008 632898 85050 633134
rect 85286 632898 85328 633134
rect 85008 632866 85328 632898
rect 115728 633454 116048 633486
rect 115728 633218 115770 633454
rect 116006 633218 116048 633454
rect 115728 633134 116048 633218
rect 115728 632898 115770 633134
rect 116006 632898 116048 633134
rect 115728 632866 116048 632898
rect 146448 633454 146768 633486
rect 146448 633218 146490 633454
rect 146726 633218 146768 633454
rect 146448 633134 146768 633218
rect 146448 632898 146490 633134
rect 146726 632898 146768 633134
rect 146448 632866 146768 632898
rect 177168 633454 177488 633486
rect 177168 633218 177210 633454
rect 177446 633218 177488 633454
rect 177168 633134 177488 633218
rect 177168 632898 177210 633134
rect 177446 632898 177488 633134
rect 177168 632866 177488 632898
rect 207888 633454 208208 633486
rect 207888 633218 207930 633454
rect 208166 633218 208208 633454
rect 207888 633134 208208 633218
rect 207888 632898 207930 633134
rect 208166 632898 208208 633134
rect 207888 632866 208208 632898
rect 238608 633454 238928 633486
rect 238608 633218 238650 633454
rect 238886 633218 238928 633454
rect 238608 633134 238928 633218
rect 238608 632898 238650 633134
rect 238886 632898 238928 633134
rect 238608 632866 238928 632898
rect 269328 633454 269648 633486
rect 269328 633218 269370 633454
rect 269606 633218 269648 633454
rect 269328 633134 269648 633218
rect 269328 632898 269370 633134
rect 269606 632898 269648 633134
rect 269328 632866 269648 632898
rect 300048 633454 300368 633486
rect 300048 633218 300090 633454
rect 300326 633218 300368 633454
rect 300048 633134 300368 633218
rect 300048 632898 300090 633134
rect 300326 632898 300368 633134
rect 300048 632866 300368 632898
rect 330768 633454 331088 633486
rect 330768 633218 330810 633454
rect 331046 633218 331088 633454
rect 330768 633134 331088 633218
rect 330768 632898 330810 633134
rect 331046 632898 331088 633134
rect 330768 632866 331088 632898
rect 361488 633454 361808 633486
rect 361488 633218 361530 633454
rect 361766 633218 361808 633454
rect 361488 633134 361808 633218
rect 361488 632898 361530 633134
rect 361766 632898 361808 633134
rect 361488 632866 361808 632898
rect 392208 633454 392528 633486
rect 392208 633218 392250 633454
rect 392486 633218 392528 633454
rect 392208 633134 392528 633218
rect 392208 632898 392250 633134
rect 392486 632898 392528 633134
rect 392208 632866 392528 632898
rect 422928 633454 423248 633486
rect 422928 633218 422970 633454
rect 423206 633218 423248 633454
rect 422928 633134 423248 633218
rect 422928 632898 422970 633134
rect 423206 632898 423248 633134
rect 422928 632866 423248 632898
rect 453648 633454 453968 633486
rect 453648 633218 453690 633454
rect 453926 633218 453968 633454
rect 453648 633134 453968 633218
rect 453648 632898 453690 633134
rect 453926 632898 453968 633134
rect 453648 632866 453968 632898
rect 484368 633454 484688 633486
rect 484368 633218 484410 633454
rect 484646 633218 484688 633454
rect 484368 633134 484688 633218
rect 484368 632898 484410 633134
rect 484646 632898 484688 633134
rect 484368 632866 484688 632898
rect 515088 633454 515408 633486
rect 515088 633218 515130 633454
rect 515366 633218 515408 633454
rect 515088 633134 515408 633218
rect 515088 632898 515130 633134
rect 515366 632898 515408 633134
rect 515088 632866 515408 632898
rect 545808 633454 546128 633486
rect 545808 633218 545850 633454
rect 546086 633218 546128 633454
rect 545808 633134 546128 633218
rect 545808 632898 545850 633134
rect 546086 632898 546128 633134
rect 545808 632866 546128 632898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect 8208 615454 8528 615486
rect 8208 615218 8250 615454
rect 8486 615218 8528 615454
rect 8208 615134 8528 615218
rect 8208 614898 8250 615134
rect 8486 614898 8528 615134
rect 8208 614866 8528 614898
rect 38928 615454 39248 615486
rect 38928 615218 38970 615454
rect 39206 615218 39248 615454
rect 38928 615134 39248 615218
rect 38928 614898 38970 615134
rect 39206 614898 39248 615134
rect 38928 614866 39248 614898
rect 69648 615454 69968 615486
rect 69648 615218 69690 615454
rect 69926 615218 69968 615454
rect 69648 615134 69968 615218
rect 69648 614898 69690 615134
rect 69926 614898 69968 615134
rect 69648 614866 69968 614898
rect 100368 615454 100688 615486
rect 100368 615218 100410 615454
rect 100646 615218 100688 615454
rect 100368 615134 100688 615218
rect 100368 614898 100410 615134
rect 100646 614898 100688 615134
rect 100368 614866 100688 614898
rect 131088 615454 131408 615486
rect 131088 615218 131130 615454
rect 131366 615218 131408 615454
rect 131088 615134 131408 615218
rect 131088 614898 131130 615134
rect 131366 614898 131408 615134
rect 131088 614866 131408 614898
rect 161808 615454 162128 615486
rect 161808 615218 161850 615454
rect 162086 615218 162128 615454
rect 161808 615134 162128 615218
rect 161808 614898 161850 615134
rect 162086 614898 162128 615134
rect 161808 614866 162128 614898
rect 192528 615454 192848 615486
rect 192528 615218 192570 615454
rect 192806 615218 192848 615454
rect 192528 615134 192848 615218
rect 192528 614898 192570 615134
rect 192806 614898 192848 615134
rect 192528 614866 192848 614898
rect 223248 615454 223568 615486
rect 223248 615218 223290 615454
rect 223526 615218 223568 615454
rect 223248 615134 223568 615218
rect 223248 614898 223290 615134
rect 223526 614898 223568 615134
rect 223248 614866 223568 614898
rect 253968 615454 254288 615486
rect 253968 615218 254010 615454
rect 254246 615218 254288 615454
rect 253968 615134 254288 615218
rect 253968 614898 254010 615134
rect 254246 614898 254288 615134
rect 253968 614866 254288 614898
rect 284688 615454 285008 615486
rect 284688 615218 284730 615454
rect 284966 615218 285008 615454
rect 284688 615134 285008 615218
rect 284688 614898 284730 615134
rect 284966 614898 285008 615134
rect 284688 614866 285008 614898
rect 315408 615454 315728 615486
rect 315408 615218 315450 615454
rect 315686 615218 315728 615454
rect 315408 615134 315728 615218
rect 315408 614898 315450 615134
rect 315686 614898 315728 615134
rect 315408 614866 315728 614898
rect 346128 615454 346448 615486
rect 346128 615218 346170 615454
rect 346406 615218 346448 615454
rect 346128 615134 346448 615218
rect 346128 614898 346170 615134
rect 346406 614898 346448 615134
rect 346128 614866 346448 614898
rect 376848 615454 377168 615486
rect 376848 615218 376890 615454
rect 377126 615218 377168 615454
rect 376848 615134 377168 615218
rect 376848 614898 376890 615134
rect 377126 614898 377168 615134
rect 376848 614866 377168 614898
rect 407568 615454 407888 615486
rect 407568 615218 407610 615454
rect 407846 615218 407888 615454
rect 407568 615134 407888 615218
rect 407568 614898 407610 615134
rect 407846 614898 407888 615134
rect 407568 614866 407888 614898
rect 438288 615454 438608 615486
rect 438288 615218 438330 615454
rect 438566 615218 438608 615454
rect 438288 615134 438608 615218
rect 438288 614898 438330 615134
rect 438566 614898 438608 615134
rect 438288 614866 438608 614898
rect 469008 615454 469328 615486
rect 469008 615218 469050 615454
rect 469286 615218 469328 615454
rect 469008 615134 469328 615218
rect 469008 614898 469050 615134
rect 469286 614898 469328 615134
rect 469008 614866 469328 614898
rect 499728 615454 500048 615486
rect 499728 615218 499770 615454
rect 500006 615218 500048 615454
rect 499728 615134 500048 615218
rect 499728 614898 499770 615134
rect 500006 614898 500048 615134
rect 499728 614866 500048 614898
rect 530448 615454 530768 615486
rect 530448 615218 530490 615454
rect 530726 615218 530768 615454
rect 530448 615134 530768 615218
rect 530448 614898 530490 615134
rect 530726 614898 530768 615134
rect 530448 614866 530768 614898
rect 561168 615454 561488 615486
rect 561168 615218 561210 615454
rect 561446 615218 561488 615454
rect 561168 615134 561488 615218
rect 561168 614898 561210 615134
rect 561446 614898 561488 615134
rect 561168 614866 561488 614898
rect 567234 604894 567854 640338
rect 567234 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 567854 604894
rect 567234 604574 567854 604658
rect 567234 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 567854 604574
rect 23568 597454 23888 597486
rect 23568 597218 23610 597454
rect 23846 597218 23888 597454
rect 23568 597134 23888 597218
rect 23568 596898 23610 597134
rect 23846 596898 23888 597134
rect 23568 596866 23888 596898
rect 54288 597454 54608 597486
rect 54288 597218 54330 597454
rect 54566 597218 54608 597454
rect 54288 597134 54608 597218
rect 54288 596898 54330 597134
rect 54566 596898 54608 597134
rect 54288 596866 54608 596898
rect 85008 597454 85328 597486
rect 85008 597218 85050 597454
rect 85286 597218 85328 597454
rect 85008 597134 85328 597218
rect 85008 596898 85050 597134
rect 85286 596898 85328 597134
rect 85008 596866 85328 596898
rect 115728 597454 116048 597486
rect 115728 597218 115770 597454
rect 116006 597218 116048 597454
rect 115728 597134 116048 597218
rect 115728 596898 115770 597134
rect 116006 596898 116048 597134
rect 115728 596866 116048 596898
rect 146448 597454 146768 597486
rect 146448 597218 146490 597454
rect 146726 597218 146768 597454
rect 146448 597134 146768 597218
rect 146448 596898 146490 597134
rect 146726 596898 146768 597134
rect 146448 596866 146768 596898
rect 177168 597454 177488 597486
rect 177168 597218 177210 597454
rect 177446 597218 177488 597454
rect 177168 597134 177488 597218
rect 177168 596898 177210 597134
rect 177446 596898 177488 597134
rect 177168 596866 177488 596898
rect 207888 597454 208208 597486
rect 207888 597218 207930 597454
rect 208166 597218 208208 597454
rect 207888 597134 208208 597218
rect 207888 596898 207930 597134
rect 208166 596898 208208 597134
rect 207888 596866 208208 596898
rect 238608 597454 238928 597486
rect 238608 597218 238650 597454
rect 238886 597218 238928 597454
rect 238608 597134 238928 597218
rect 238608 596898 238650 597134
rect 238886 596898 238928 597134
rect 238608 596866 238928 596898
rect 269328 597454 269648 597486
rect 269328 597218 269370 597454
rect 269606 597218 269648 597454
rect 269328 597134 269648 597218
rect 269328 596898 269370 597134
rect 269606 596898 269648 597134
rect 269328 596866 269648 596898
rect 300048 597454 300368 597486
rect 300048 597218 300090 597454
rect 300326 597218 300368 597454
rect 300048 597134 300368 597218
rect 300048 596898 300090 597134
rect 300326 596898 300368 597134
rect 300048 596866 300368 596898
rect 330768 597454 331088 597486
rect 330768 597218 330810 597454
rect 331046 597218 331088 597454
rect 330768 597134 331088 597218
rect 330768 596898 330810 597134
rect 331046 596898 331088 597134
rect 330768 596866 331088 596898
rect 361488 597454 361808 597486
rect 361488 597218 361530 597454
rect 361766 597218 361808 597454
rect 361488 597134 361808 597218
rect 361488 596898 361530 597134
rect 361766 596898 361808 597134
rect 361488 596866 361808 596898
rect 392208 597454 392528 597486
rect 392208 597218 392250 597454
rect 392486 597218 392528 597454
rect 392208 597134 392528 597218
rect 392208 596898 392250 597134
rect 392486 596898 392528 597134
rect 392208 596866 392528 596898
rect 422928 597454 423248 597486
rect 422928 597218 422970 597454
rect 423206 597218 423248 597454
rect 422928 597134 423248 597218
rect 422928 596898 422970 597134
rect 423206 596898 423248 597134
rect 422928 596866 423248 596898
rect 453648 597454 453968 597486
rect 453648 597218 453690 597454
rect 453926 597218 453968 597454
rect 453648 597134 453968 597218
rect 453648 596898 453690 597134
rect 453926 596898 453968 597134
rect 453648 596866 453968 596898
rect 484368 597454 484688 597486
rect 484368 597218 484410 597454
rect 484646 597218 484688 597454
rect 484368 597134 484688 597218
rect 484368 596898 484410 597134
rect 484646 596898 484688 597134
rect 484368 596866 484688 596898
rect 515088 597454 515408 597486
rect 515088 597218 515130 597454
rect 515366 597218 515408 597454
rect 515088 597134 515408 597218
rect 515088 596898 515130 597134
rect 515366 596898 515408 597134
rect 515088 596866 515408 596898
rect 545808 597454 546128 597486
rect 545808 597218 545850 597454
rect 546086 597218 546128 597454
rect 545808 597134 546128 597218
rect 545808 596898 545850 597134
rect 546086 596898 546128 597134
rect 545808 596866 546128 596898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect 8208 579454 8528 579486
rect 8208 579218 8250 579454
rect 8486 579218 8528 579454
rect 8208 579134 8528 579218
rect 8208 578898 8250 579134
rect 8486 578898 8528 579134
rect 8208 578866 8528 578898
rect 38928 579454 39248 579486
rect 38928 579218 38970 579454
rect 39206 579218 39248 579454
rect 38928 579134 39248 579218
rect 38928 578898 38970 579134
rect 39206 578898 39248 579134
rect 38928 578866 39248 578898
rect 69648 579454 69968 579486
rect 69648 579218 69690 579454
rect 69926 579218 69968 579454
rect 69648 579134 69968 579218
rect 69648 578898 69690 579134
rect 69926 578898 69968 579134
rect 69648 578866 69968 578898
rect 100368 579454 100688 579486
rect 100368 579218 100410 579454
rect 100646 579218 100688 579454
rect 100368 579134 100688 579218
rect 100368 578898 100410 579134
rect 100646 578898 100688 579134
rect 100368 578866 100688 578898
rect 131088 579454 131408 579486
rect 131088 579218 131130 579454
rect 131366 579218 131408 579454
rect 131088 579134 131408 579218
rect 131088 578898 131130 579134
rect 131366 578898 131408 579134
rect 131088 578866 131408 578898
rect 161808 579454 162128 579486
rect 161808 579218 161850 579454
rect 162086 579218 162128 579454
rect 161808 579134 162128 579218
rect 161808 578898 161850 579134
rect 162086 578898 162128 579134
rect 161808 578866 162128 578898
rect 192528 579454 192848 579486
rect 192528 579218 192570 579454
rect 192806 579218 192848 579454
rect 192528 579134 192848 579218
rect 192528 578898 192570 579134
rect 192806 578898 192848 579134
rect 192528 578866 192848 578898
rect 223248 579454 223568 579486
rect 223248 579218 223290 579454
rect 223526 579218 223568 579454
rect 223248 579134 223568 579218
rect 223248 578898 223290 579134
rect 223526 578898 223568 579134
rect 223248 578866 223568 578898
rect 253968 579454 254288 579486
rect 253968 579218 254010 579454
rect 254246 579218 254288 579454
rect 253968 579134 254288 579218
rect 253968 578898 254010 579134
rect 254246 578898 254288 579134
rect 253968 578866 254288 578898
rect 284688 579454 285008 579486
rect 284688 579218 284730 579454
rect 284966 579218 285008 579454
rect 284688 579134 285008 579218
rect 284688 578898 284730 579134
rect 284966 578898 285008 579134
rect 284688 578866 285008 578898
rect 315408 579454 315728 579486
rect 315408 579218 315450 579454
rect 315686 579218 315728 579454
rect 315408 579134 315728 579218
rect 315408 578898 315450 579134
rect 315686 578898 315728 579134
rect 315408 578866 315728 578898
rect 346128 579454 346448 579486
rect 346128 579218 346170 579454
rect 346406 579218 346448 579454
rect 346128 579134 346448 579218
rect 346128 578898 346170 579134
rect 346406 578898 346448 579134
rect 346128 578866 346448 578898
rect 376848 579454 377168 579486
rect 376848 579218 376890 579454
rect 377126 579218 377168 579454
rect 376848 579134 377168 579218
rect 376848 578898 376890 579134
rect 377126 578898 377168 579134
rect 376848 578866 377168 578898
rect 407568 579454 407888 579486
rect 407568 579218 407610 579454
rect 407846 579218 407888 579454
rect 407568 579134 407888 579218
rect 407568 578898 407610 579134
rect 407846 578898 407888 579134
rect 407568 578866 407888 578898
rect 438288 579454 438608 579486
rect 438288 579218 438330 579454
rect 438566 579218 438608 579454
rect 438288 579134 438608 579218
rect 438288 578898 438330 579134
rect 438566 578898 438608 579134
rect 438288 578866 438608 578898
rect 469008 579454 469328 579486
rect 469008 579218 469050 579454
rect 469286 579218 469328 579454
rect 469008 579134 469328 579218
rect 469008 578898 469050 579134
rect 469286 578898 469328 579134
rect 469008 578866 469328 578898
rect 499728 579454 500048 579486
rect 499728 579218 499770 579454
rect 500006 579218 500048 579454
rect 499728 579134 500048 579218
rect 499728 578898 499770 579134
rect 500006 578898 500048 579134
rect 499728 578866 500048 578898
rect 530448 579454 530768 579486
rect 530448 579218 530490 579454
rect 530726 579218 530768 579454
rect 530448 579134 530768 579218
rect 530448 578898 530490 579134
rect 530726 578898 530768 579134
rect 530448 578866 530768 578898
rect 561168 579454 561488 579486
rect 561168 579218 561210 579454
rect 561446 579218 561488 579454
rect 561168 579134 561488 579218
rect 561168 578898 561210 579134
rect 561446 578898 561488 579134
rect 561168 578866 561488 578898
rect 567234 568894 567854 604338
rect 567234 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 567854 568894
rect 567234 568574 567854 568658
rect 567234 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 567854 568574
rect 23568 561454 23888 561486
rect 23568 561218 23610 561454
rect 23846 561218 23888 561454
rect 23568 561134 23888 561218
rect 23568 560898 23610 561134
rect 23846 560898 23888 561134
rect 23568 560866 23888 560898
rect 54288 561454 54608 561486
rect 54288 561218 54330 561454
rect 54566 561218 54608 561454
rect 54288 561134 54608 561218
rect 54288 560898 54330 561134
rect 54566 560898 54608 561134
rect 54288 560866 54608 560898
rect 85008 561454 85328 561486
rect 85008 561218 85050 561454
rect 85286 561218 85328 561454
rect 85008 561134 85328 561218
rect 85008 560898 85050 561134
rect 85286 560898 85328 561134
rect 85008 560866 85328 560898
rect 115728 561454 116048 561486
rect 115728 561218 115770 561454
rect 116006 561218 116048 561454
rect 115728 561134 116048 561218
rect 115728 560898 115770 561134
rect 116006 560898 116048 561134
rect 115728 560866 116048 560898
rect 146448 561454 146768 561486
rect 146448 561218 146490 561454
rect 146726 561218 146768 561454
rect 146448 561134 146768 561218
rect 146448 560898 146490 561134
rect 146726 560898 146768 561134
rect 146448 560866 146768 560898
rect 177168 561454 177488 561486
rect 177168 561218 177210 561454
rect 177446 561218 177488 561454
rect 177168 561134 177488 561218
rect 177168 560898 177210 561134
rect 177446 560898 177488 561134
rect 177168 560866 177488 560898
rect 207888 561454 208208 561486
rect 207888 561218 207930 561454
rect 208166 561218 208208 561454
rect 207888 561134 208208 561218
rect 207888 560898 207930 561134
rect 208166 560898 208208 561134
rect 207888 560866 208208 560898
rect 238608 561454 238928 561486
rect 238608 561218 238650 561454
rect 238886 561218 238928 561454
rect 238608 561134 238928 561218
rect 238608 560898 238650 561134
rect 238886 560898 238928 561134
rect 238608 560866 238928 560898
rect 269328 561454 269648 561486
rect 269328 561218 269370 561454
rect 269606 561218 269648 561454
rect 269328 561134 269648 561218
rect 269328 560898 269370 561134
rect 269606 560898 269648 561134
rect 269328 560866 269648 560898
rect 300048 561454 300368 561486
rect 300048 561218 300090 561454
rect 300326 561218 300368 561454
rect 300048 561134 300368 561218
rect 300048 560898 300090 561134
rect 300326 560898 300368 561134
rect 300048 560866 300368 560898
rect 330768 561454 331088 561486
rect 330768 561218 330810 561454
rect 331046 561218 331088 561454
rect 330768 561134 331088 561218
rect 330768 560898 330810 561134
rect 331046 560898 331088 561134
rect 330768 560866 331088 560898
rect 361488 561454 361808 561486
rect 361488 561218 361530 561454
rect 361766 561218 361808 561454
rect 361488 561134 361808 561218
rect 361488 560898 361530 561134
rect 361766 560898 361808 561134
rect 361488 560866 361808 560898
rect 392208 561454 392528 561486
rect 392208 561218 392250 561454
rect 392486 561218 392528 561454
rect 392208 561134 392528 561218
rect 392208 560898 392250 561134
rect 392486 560898 392528 561134
rect 392208 560866 392528 560898
rect 422928 561454 423248 561486
rect 422928 561218 422970 561454
rect 423206 561218 423248 561454
rect 422928 561134 423248 561218
rect 422928 560898 422970 561134
rect 423206 560898 423248 561134
rect 422928 560866 423248 560898
rect 453648 561454 453968 561486
rect 453648 561218 453690 561454
rect 453926 561218 453968 561454
rect 453648 561134 453968 561218
rect 453648 560898 453690 561134
rect 453926 560898 453968 561134
rect 453648 560866 453968 560898
rect 484368 561454 484688 561486
rect 484368 561218 484410 561454
rect 484646 561218 484688 561454
rect 484368 561134 484688 561218
rect 484368 560898 484410 561134
rect 484646 560898 484688 561134
rect 484368 560866 484688 560898
rect 515088 561454 515408 561486
rect 515088 561218 515130 561454
rect 515366 561218 515408 561454
rect 515088 561134 515408 561218
rect 515088 560898 515130 561134
rect 515366 560898 515408 561134
rect 515088 560866 515408 560898
rect 545808 561454 546128 561486
rect 545808 561218 545850 561454
rect 546086 561218 546128 561454
rect 545808 561134 546128 561218
rect 545808 560898 545850 561134
rect 546086 560898 546128 561134
rect 545808 560866 546128 560898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect 8208 543454 8528 543486
rect 8208 543218 8250 543454
rect 8486 543218 8528 543454
rect 8208 543134 8528 543218
rect 8208 542898 8250 543134
rect 8486 542898 8528 543134
rect 8208 542866 8528 542898
rect 38928 543454 39248 543486
rect 38928 543218 38970 543454
rect 39206 543218 39248 543454
rect 38928 543134 39248 543218
rect 38928 542898 38970 543134
rect 39206 542898 39248 543134
rect 38928 542866 39248 542898
rect 69648 543454 69968 543486
rect 69648 543218 69690 543454
rect 69926 543218 69968 543454
rect 69648 543134 69968 543218
rect 69648 542898 69690 543134
rect 69926 542898 69968 543134
rect 69648 542866 69968 542898
rect 100368 543454 100688 543486
rect 100368 543218 100410 543454
rect 100646 543218 100688 543454
rect 100368 543134 100688 543218
rect 100368 542898 100410 543134
rect 100646 542898 100688 543134
rect 100368 542866 100688 542898
rect 131088 543454 131408 543486
rect 131088 543218 131130 543454
rect 131366 543218 131408 543454
rect 131088 543134 131408 543218
rect 131088 542898 131130 543134
rect 131366 542898 131408 543134
rect 131088 542866 131408 542898
rect 161808 543454 162128 543486
rect 161808 543218 161850 543454
rect 162086 543218 162128 543454
rect 161808 543134 162128 543218
rect 161808 542898 161850 543134
rect 162086 542898 162128 543134
rect 161808 542866 162128 542898
rect 192528 543454 192848 543486
rect 192528 543218 192570 543454
rect 192806 543218 192848 543454
rect 192528 543134 192848 543218
rect 192528 542898 192570 543134
rect 192806 542898 192848 543134
rect 192528 542866 192848 542898
rect 223248 543454 223568 543486
rect 223248 543218 223290 543454
rect 223526 543218 223568 543454
rect 223248 543134 223568 543218
rect 223248 542898 223290 543134
rect 223526 542898 223568 543134
rect 223248 542866 223568 542898
rect 253968 543454 254288 543486
rect 253968 543218 254010 543454
rect 254246 543218 254288 543454
rect 253968 543134 254288 543218
rect 253968 542898 254010 543134
rect 254246 542898 254288 543134
rect 253968 542866 254288 542898
rect 284688 543454 285008 543486
rect 284688 543218 284730 543454
rect 284966 543218 285008 543454
rect 284688 543134 285008 543218
rect 284688 542898 284730 543134
rect 284966 542898 285008 543134
rect 284688 542866 285008 542898
rect 315408 543454 315728 543486
rect 315408 543218 315450 543454
rect 315686 543218 315728 543454
rect 315408 543134 315728 543218
rect 315408 542898 315450 543134
rect 315686 542898 315728 543134
rect 315408 542866 315728 542898
rect 346128 543454 346448 543486
rect 346128 543218 346170 543454
rect 346406 543218 346448 543454
rect 346128 543134 346448 543218
rect 346128 542898 346170 543134
rect 346406 542898 346448 543134
rect 346128 542866 346448 542898
rect 376848 543454 377168 543486
rect 376848 543218 376890 543454
rect 377126 543218 377168 543454
rect 376848 543134 377168 543218
rect 376848 542898 376890 543134
rect 377126 542898 377168 543134
rect 376848 542866 377168 542898
rect 407568 543454 407888 543486
rect 407568 543218 407610 543454
rect 407846 543218 407888 543454
rect 407568 543134 407888 543218
rect 407568 542898 407610 543134
rect 407846 542898 407888 543134
rect 407568 542866 407888 542898
rect 438288 543454 438608 543486
rect 438288 543218 438330 543454
rect 438566 543218 438608 543454
rect 438288 543134 438608 543218
rect 438288 542898 438330 543134
rect 438566 542898 438608 543134
rect 438288 542866 438608 542898
rect 469008 543454 469328 543486
rect 469008 543218 469050 543454
rect 469286 543218 469328 543454
rect 469008 543134 469328 543218
rect 469008 542898 469050 543134
rect 469286 542898 469328 543134
rect 469008 542866 469328 542898
rect 499728 543454 500048 543486
rect 499728 543218 499770 543454
rect 500006 543218 500048 543454
rect 499728 543134 500048 543218
rect 499728 542898 499770 543134
rect 500006 542898 500048 543134
rect 499728 542866 500048 542898
rect 530448 543454 530768 543486
rect 530448 543218 530490 543454
rect 530726 543218 530768 543454
rect 530448 543134 530768 543218
rect 530448 542898 530490 543134
rect 530726 542898 530768 543134
rect 530448 542866 530768 542898
rect 561168 543454 561488 543486
rect 561168 543218 561210 543454
rect 561446 543218 561488 543454
rect 561168 543134 561488 543218
rect 561168 542898 561210 543134
rect 561446 542898 561488 543134
rect 561168 542866 561488 542898
rect 567234 532894 567854 568338
rect 567234 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 567854 532894
rect 567234 532574 567854 532658
rect 567234 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 567854 532574
rect 23568 525454 23888 525486
rect 23568 525218 23610 525454
rect 23846 525218 23888 525454
rect 23568 525134 23888 525218
rect 23568 524898 23610 525134
rect 23846 524898 23888 525134
rect 23568 524866 23888 524898
rect 54288 525454 54608 525486
rect 54288 525218 54330 525454
rect 54566 525218 54608 525454
rect 54288 525134 54608 525218
rect 54288 524898 54330 525134
rect 54566 524898 54608 525134
rect 54288 524866 54608 524898
rect 85008 525454 85328 525486
rect 85008 525218 85050 525454
rect 85286 525218 85328 525454
rect 85008 525134 85328 525218
rect 85008 524898 85050 525134
rect 85286 524898 85328 525134
rect 85008 524866 85328 524898
rect 115728 525454 116048 525486
rect 115728 525218 115770 525454
rect 116006 525218 116048 525454
rect 115728 525134 116048 525218
rect 115728 524898 115770 525134
rect 116006 524898 116048 525134
rect 115728 524866 116048 524898
rect 146448 525454 146768 525486
rect 146448 525218 146490 525454
rect 146726 525218 146768 525454
rect 146448 525134 146768 525218
rect 146448 524898 146490 525134
rect 146726 524898 146768 525134
rect 146448 524866 146768 524898
rect 177168 525454 177488 525486
rect 177168 525218 177210 525454
rect 177446 525218 177488 525454
rect 177168 525134 177488 525218
rect 177168 524898 177210 525134
rect 177446 524898 177488 525134
rect 177168 524866 177488 524898
rect 207888 525454 208208 525486
rect 207888 525218 207930 525454
rect 208166 525218 208208 525454
rect 207888 525134 208208 525218
rect 207888 524898 207930 525134
rect 208166 524898 208208 525134
rect 207888 524866 208208 524898
rect 238608 525454 238928 525486
rect 238608 525218 238650 525454
rect 238886 525218 238928 525454
rect 238608 525134 238928 525218
rect 238608 524898 238650 525134
rect 238886 524898 238928 525134
rect 238608 524866 238928 524898
rect 269328 525454 269648 525486
rect 269328 525218 269370 525454
rect 269606 525218 269648 525454
rect 269328 525134 269648 525218
rect 269328 524898 269370 525134
rect 269606 524898 269648 525134
rect 269328 524866 269648 524898
rect 300048 525454 300368 525486
rect 300048 525218 300090 525454
rect 300326 525218 300368 525454
rect 300048 525134 300368 525218
rect 300048 524898 300090 525134
rect 300326 524898 300368 525134
rect 300048 524866 300368 524898
rect 330768 525454 331088 525486
rect 330768 525218 330810 525454
rect 331046 525218 331088 525454
rect 330768 525134 331088 525218
rect 330768 524898 330810 525134
rect 331046 524898 331088 525134
rect 330768 524866 331088 524898
rect 361488 525454 361808 525486
rect 361488 525218 361530 525454
rect 361766 525218 361808 525454
rect 361488 525134 361808 525218
rect 361488 524898 361530 525134
rect 361766 524898 361808 525134
rect 361488 524866 361808 524898
rect 392208 525454 392528 525486
rect 392208 525218 392250 525454
rect 392486 525218 392528 525454
rect 392208 525134 392528 525218
rect 392208 524898 392250 525134
rect 392486 524898 392528 525134
rect 392208 524866 392528 524898
rect 422928 525454 423248 525486
rect 422928 525218 422970 525454
rect 423206 525218 423248 525454
rect 422928 525134 423248 525218
rect 422928 524898 422970 525134
rect 423206 524898 423248 525134
rect 422928 524866 423248 524898
rect 453648 525454 453968 525486
rect 453648 525218 453690 525454
rect 453926 525218 453968 525454
rect 453648 525134 453968 525218
rect 453648 524898 453690 525134
rect 453926 524898 453968 525134
rect 453648 524866 453968 524898
rect 484368 525454 484688 525486
rect 484368 525218 484410 525454
rect 484646 525218 484688 525454
rect 484368 525134 484688 525218
rect 484368 524898 484410 525134
rect 484646 524898 484688 525134
rect 484368 524866 484688 524898
rect 515088 525454 515408 525486
rect 515088 525218 515130 525454
rect 515366 525218 515408 525454
rect 515088 525134 515408 525218
rect 515088 524898 515130 525134
rect 515366 524898 515408 525134
rect 515088 524866 515408 524898
rect 545808 525454 546128 525486
rect 545808 525218 545850 525454
rect 546086 525218 546128 525454
rect 545808 525134 546128 525218
rect 545808 524898 545850 525134
rect 546086 524898 546128 525134
rect 545808 524866 546128 524898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect 8208 507454 8528 507486
rect 8208 507218 8250 507454
rect 8486 507218 8528 507454
rect 8208 507134 8528 507218
rect 8208 506898 8250 507134
rect 8486 506898 8528 507134
rect 8208 506866 8528 506898
rect 38928 507454 39248 507486
rect 38928 507218 38970 507454
rect 39206 507218 39248 507454
rect 38928 507134 39248 507218
rect 38928 506898 38970 507134
rect 39206 506898 39248 507134
rect 38928 506866 39248 506898
rect 69648 507454 69968 507486
rect 69648 507218 69690 507454
rect 69926 507218 69968 507454
rect 69648 507134 69968 507218
rect 69648 506898 69690 507134
rect 69926 506898 69968 507134
rect 69648 506866 69968 506898
rect 100368 507454 100688 507486
rect 100368 507218 100410 507454
rect 100646 507218 100688 507454
rect 100368 507134 100688 507218
rect 100368 506898 100410 507134
rect 100646 506898 100688 507134
rect 100368 506866 100688 506898
rect 131088 507454 131408 507486
rect 131088 507218 131130 507454
rect 131366 507218 131408 507454
rect 131088 507134 131408 507218
rect 131088 506898 131130 507134
rect 131366 506898 131408 507134
rect 131088 506866 131408 506898
rect 161808 507454 162128 507486
rect 161808 507218 161850 507454
rect 162086 507218 162128 507454
rect 161808 507134 162128 507218
rect 161808 506898 161850 507134
rect 162086 506898 162128 507134
rect 161808 506866 162128 506898
rect 192528 507454 192848 507486
rect 192528 507218 192570 507454
rect 192806 507218 192848 507454
rect 192528 507134 192848 507218
rect 192528 506898 192570 507134
rect 192806 506898 192848 507134
rect 192528 506866 192848 506898
rect 223248 507454 223568 507486
rect 223248 507218 223290 507454
rect 223526 507218 223568 507454
rect 223248 507134 223568 507218
rect 223248 506898 223290 507134
rect 223526 506898 223568 507134
rect 223248 506866 223568 506898
rect 253968 507454 254288 507486
rect 253968 507218 254010 507454
rect 254246 507218 254288 507454
rect 253968 507134 254288 507218
rect 253968 506898 254010 507134
rect 254246 506898 254288 507134
rect 253968 506866 254288 506898
rect 284688 507454 285008 507486
rect 284688 507218 284730 507454
rect 284966 507218 285008 507454
rect 284688 507134 285008 507218
rect 284688 506898 284730 507134
rect 284966 506898 285008 507134
rect 284688 506866 285008 506898
rect 315408 507454 315728 507486
rect 315408 507218 315450 507454
rect 315686 507218 315728 507454
rect 315408 507134 315728 507218
rect 315408 506898 315450 507134
rect 315686 506898 315728 507134
rect 315408 506866 315728 506898
rect 346128 507454 346448 507486
rect 346128 507218 346170 507454
rect 346406 507218 346448 507454
rect 346128 507134 346448 507218
rect 346128 506898 346170 507134
rect 346406 506898 346448 507134
rect 346128 506866 346448 506898
rect 376848 507454 377168 507486
rect 376848 507218 376890 507454
rect 377126 507218 377168 507454
rect 376848 507134 377168 507218
rect 376848 506898 376890 507134
rect 377126 506898 377168 507134
rect 376848 506866 377168 506898
rect 407568 507454 407888 507486
rect 407568 507218 407610 507454
rect 407846 507218 407888 507454
rect 407568 507134 407888 507218
rect 407568 506898 407610 507134
rect 407846 506898 407888 507134
rect 407568 506866 407888 506898
rect 438288 507454 438608 507486
rect 438288 507218 438330 507454
rect 438566 507218 438608 507454
rect 438288 507134 438608 507218
rect 438288 506898 438330 507134
rect 438566 506898 438608 507134
rect 438288 506866 438608 506898
rect 469008 507454 469328 507486
rect 469008 507218 469050 507454
rect 469286 507218 469328 507454
rect 469008 507134 469328 507218
rect 469008 506898 469050 507134
rect 469286 506898 469328 507134
rect 469008 506866 469328 506898
rect 499728 507454 500048 507486
rect 499728 507218 499770 507454
rect 500006 507218 500048 507454
rect 499728 507134 500048 507218
rect 499728 506898 499770 507134
rect 500006 506898 500048 507134
rect 499728 506866 500048 506898
rect 530448 507454 530768 507486
rect 530448 507218 530490 507454
rect 530726 507218 530768 507454
rect 530448 507134 530768 507218
rect 530448 506898 530490 507134
rect 530726 506898 530768 507134
rect 530448 506866 530768 506898
rect 561168 507454 561488 507486
rect 561168 507218 561210 507454
rect 561446 507218 561488 507454
rect 561168 507134 561488 507218
rect 561168 506898 561210 507134
rect 561446 506898 561488 507134
rect 561168 506866 561488 506898
rect 567234 496894 567854 532338
rect 567234 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 567854 496894
rect 567234 496574 567854 496658
rect 567234 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 567854 496574
rect 23568 489454 23888 489486
rect 23568 489218 23610 489454
rect 23846 489218 23888 489454
rect 23568 489134 23888 489218
rect 23568 488898 23610 489134
rect 23846 488898 23888 489134
rect 23568 488866 23888 488898
rect 54288 489454 54608 489486
rect 54288 489218 54330 489454
rect 54566 489218 54608 489454
rect 54288 489134 54608 489218
rect 54288 488898 54330 489134
rect 54566 488898 54608 489134
rect 54288 488866 54608 488898
rect 85008 489454 85328 489486
rect 85008 489218 85050 489454
rect 85286 489218 85328 489454
rect 85008 489134 85328 489218
rect 85008 488898 85050 489134
rect 85286 488898 85328 489134
rect 85008 488866 85328 488898
rect 115728 489454 116048 489486
rect 115728 489218 115770 489454
rect 116006 489218 116048 489454
rect 115728 489134 116048 489218
rect 115728 488898 115770 489134
rect 116006 488898 116048 489134
rect 115728 488866 116048 488898
rect 146448 489454 146768 489486
rect 146448 489218 146490 489454
rect 146726 489218 146768 489454
rect 146448 489134 146768 489218
rect 146448 488898 146490 489134
rect 146726 488898 146768 489134
rect 146448 488866 146768 488898
rect 177168 489454 177488 489486
rect 177168 489218 177210 489454
rect 177446 489218 177488 489454
rect 177168 489134 177488 489218
rect 177168 488898 177210 489134
rect 177446 488898 177488 489134
rect 177168 488866 177488 488898
rect 207888 489454 208208 489486
rect 207888 489218 207930 489454
rect 208166 489218 208208 489454
rect 207888 489134 208208 489218
rect 207888 488898 207930 489134
rect 208166 488898 208208 489134
rect 207888 488866 208208 488898
rect 238608 489454 238928 489486
rect 238608 489218 238650 489454
rect 238886 489218 238928 489454
rect 238608 489134 238928 489218
rect 238608 488898 238650 489134
rect 238886 488898 238928 489134
rect 238608 488866 238928 488898
rect 269328 489454 269648 489486
rect 269328 489218 269370 489454
rect 269606 489218 269648 489454
rect 269328 489134 269648 489218
rect 269328 488898 269370 489134
rect 269606 488898 269648 489134
rect 269328 488866 269648 488898
rect 300048 489454 300368 489486
rect 300048 489218 300090 489454
rect 300326 489218 300368 489454
rect 300048 489134 300368 489218
rect 300048 488898 300090 489134
rect 300326 488898 300368 489134
rect 300048 488866 300368 488898
rect 330768 489454 331088 489486
rect 330768 489218 330810 489454
rect 331046 489218 331088 489454
rect 330768 489134 331088 489218
rect 330768 488898 330810 489134
rect 331046 488898 331088 489134
rect 330768 488866 331088 488898
rect 361488 489454 361808 489486
rect 361488 489218 361530 489454
rect 361766 489218 361808 489454
rect 361488 489134 361808 489218
rect 361488 488898 361530 489134
rect 361766 488898 361808 489134
rect 361488 488866 361808 488898
rect 392208 489454 392528 489486
rect 392208 489218 392250 489454
rect 392486 489218 392528 489454
rect 392208 489134 392528 489218
rect 392208 488898 392250 489134
rect 392486 488898 392528 489134
rect 392208 488866 392528 488898
rect 422928 489454 423248 489486
rect 422928 489218 422970 489454
rect 423206 489218 423248 489454
rect 422928 489134 423248 489218
rect 422928 488898 422970 489134
rect 423206 488898 423248 489134
rect 422928 488866 423248 488898
rect 453648 489454 453968 489486
rect 453648 489218 453690 489454
rect 453926 489218 453968 489454
rect 453648 489134 453968 489218
rect 453648 488898 453690 489134
rect 453926 488898 453968 489134
rect 453648 488866 453968 488898
rect 484368 489454 484688 489486
rect 484368 489218 484410 489454
rect 484646 489218 484688 489454
rect 484368 489134 484688 489218
rect 484368 488898 484410 489134
rect 484646 488898 484688 489134
rect 484368 488866 484688 488898
rect 515088 489454 515408 489486
rect 515088 489218 515130 489454
rect 515366 489218 515408 489454
rect 515088 489134 515408 489218
rect 515088 488898 515130 489134
rect 515366 488898 515408 489134
rect 515088 488866 515408 488898
rect 545808 489454 546128 489486
rect 545808 489218 545850 489454
rect 546086 489218 546128 489454
rect 545808 489134 546128 489218
rect 545808 488898 545850 489134
rect 546086 488898 546128 489134
rect 545808 488866 546128 488898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect 8208 471454 8528 471486
rect 8208 471218 8250 471454
rect 8486 471218 8528 471454
rect 8208 471134 8528 471218
rect 8208 470898 8250 471134
rect 8486 470898 8528 471134
rect 8208 470866 8528 470898
rect 38928 471454 39248 471486
rect 38928 471218 38970 471454
rect 39206 471218 39248 471454
rect 38928 471134 39248 471218
rect 38928 470898 38970 471134
rect 39206 470898 39248 471134
rect 38928 470866 39248 470898
rect 69648 471454 69968 471486
rect 69648 471218 69690 471454
rect 69926 471218 69968 471454
rect 69648 471134 69968 471218
rect 69648 470898 69690 471134
rect 69926 470898 69968 471134
rect 69648 470866 69968 470898
rect 100368 471454 100688 471486
rect 100368 471218 100410 471454
rect 100646 471218 100688 471454
rect 100368 471134 100688 471218
rect 100368 470898 100410 471134
rect 100646 470898 100688 471134
rect 100368 470866 100688 470898
rect 131088 471454 131408 471486
rect 131088 471218 131130 471454
rect 131366 471218 131408 471454
rect 131088 471134 131408 471218
rect 131088 470898 131130 471134
rect 131366 470898 131408 471134
rect 131088 470866 131408 470898
rect 161808 471454 162128 471486
rect 161808 471218 161850 471454
rect 162086 471218 162128 471454
rect 161808 471134 162128 471218
rect 161808 470898 161850 471134
rect 162086 470898 162128 471134
rect 161808 470866 162128 470898
rect 192528 471454 192848 471486
rect 192528 471218 192570 471454
rect 192806 471218 192848 471454
rect 192528 471134 192848 471218
rect 192528 470898 192570 471134
rect 192806 470898 192848 471134
rect 192528 470866 192848 470898
rect 223248 471454 223568 471486
rect 223248 471218 223290 471454
rect 223526 471218 223568 471454
rect 223248 471134 223568 471218
rect 223248 470898 223290 471134
rect 223526 470898 223568 471134
rect 223248 470866 223568 470898
rect 253968 471454 254288 471486
rect 253968 471218 254010 471454
rect 254246 471218 254288 471454
rect 253968 471134 254288 471218
rect 253968 470898 254010 471134
rect 254246 470898 254288 471134
rect 253968 470866 254288 470898
rect 284688 471454 285008 471486
rect 284688 471218 284730 471454
rect 284966 471218 285008 471454
rect 284688 471134 285008 471218
rect 284688 470898 284730 471134
rect 284966 470898 285008 471134
rect 284688 470866 285008 470898
rect 315408 471454 315728 471486
rect 315408 471218 315450 471454
rect 315686 471218 315728 471454
rect 315408 471134 315728 471218
rect 315408 470898 315450 471134
rect 315686 470898 315728 471134
rect 315408 470866 315728 470898
rect 346128 471454 346448 471486
rect 346128 471218 346170 471454
rect 346406 471218 346448 471454
rect 346128 471134 346448 471218
rect 346128 470898 346170 471134
rect 346406 470898 346448 471134
rect 346128 470866 346448 470898
rect 376848 471454 377168 471486
rect 376848 471218 376890 471454
rect 377126 471218 377168 471454
rect 376848 471134 377168 471218
rect 376848 470898 376890 471134
rect 377126 470898 377168 471134
rect 376848 470866 377168 470898
rect 407568 471454 407888 471486
rect 407568 471218 407610 471454
rect 407846 471218 407888 471454
rect 407568 471134 407888 471218
rect 407568 470898 407610 471134
rect 407846 470898 407888 471134
rect 407568 470866 407888 470898
rect 438288 471454 438608 471486
rect 438288 471218 438330 471454
rect 438566 471218 438608 471454
rect 438288 471134 438608 471218
rect 438288 470898 438330 471134
rect 438566 470898 438608 471134
rect 438288 470866 438608 470898
rect 469008 471454 469328 471486
rect 469008 471218 469050 471454
rect 469286 471218 469328 471454
rect 469008 471134 469328 471218
rect 469008 470898 469050 471134
rect 469286 470898 469328 471134
rect 469008 470866 469328 470898
rect 499728 471454 500048 471486
rect 499728 471218 499770 471454
rect 500006 471218 500048 471454
rect 499728 471134 500048 471218
rect 499728 470898 499770 471134
rect 500006 470898 500048 471134
rect 499728 470866 500048 470898
rect 530448 471454 530768 471486
rect 530448 471218 530490 471454
rect 530726 471218 530768 471454
rect 530448 471134 530768 471218
rect 530448 470898 530490 471134
rect 530726 470898 530768 471134
rect 530448 470866 530768 470898
rect 561168 471454 561488 471486
rect 561168 471218 561210 471454
rect 561446 471218 561488 471454
rect 561168 471134 561488 471218
rect 561168 470898 561210 471134
rect 561446 470898 561488 471134
rect 561168 470866 561488 470898
rect 567234 460894 567854 496338
rect 567234 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 567854 460894
rect 567234 460574 567854 460658
rect 567234 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 567854 460574
rect 23568 453454 23888 453486
rect 23568 453218 23610 453454
rect 23846 453218 23888 453454
rect 23568 453134 23888 453218
rect 23568 452898 23610 453134
rect 23846 452898 23888 453134
rect 23568 452866 23888 452898
rect 54288 453454 54608 453486
rect 54288 453218 54330 453454
rect 54566 453218 54608 453454
rect 54288 453134 54608 453218
rect 54288 452898 54330 453134
rect 54566 452898 54608 453134
rect 54288 452866 54608 452898
rect 85008 453454 85328 453486
rect 85008 453218 85050 453454
rect 85286 453218 85328 453454
rect 85008 453134 85328 453218
rect 85008 452898 85050 453134
rect 85286 452898 85328 453134
rect 85008 452866 85328 452898
rect 115728 453454 116048 453486
rect 115728 453218 115770 453454
rect 116006 453218 116048 453454
rect 115728 453134 116048 453218
rect 115728 452898 115770 453134
rect 116006 452898 116048 453134
rect 115728 452866 116048 452898
rect 146448 453454 146768 453486
rect 146448 453218 146490 453454
rect 146726 453218 146768 453454
rect 146448 453134 146768 453218
rect 146448 452898 146490 453134
rect 146726 452898 146768 453134
rect 146448 452866 146768 452898
rect 177168 453454 177488 453486
rect 177168 453218 177210 453454
rect 177446 453218 177488 453454
rect 177168 453134 177488 453218
rect 177168 452898 177210 453134
rect 177446 452898 177488 453134
rect 177168 452866 177488 452898
rect 207888 453454 208208 453486
rect 207888 453218 207930 453454
rect 208166 453218 208208 453454
rect 207888 453134 208208 453218
rect 207888 452898 207930 453134
rect 208166 452898 208208 453134
rect 207888 452866 208208 452898
rect 238608 453454 238928 453486
rect 238608 453218 238650 453454
rect 238886 453218 238928 453454
rect 238608 453134 238928 453218
rect 238608 452898 238650 453134
rect 238886 452898 238928 453134
rect 238608 452866 238928 452898
rect 269328 453454 269648 453486
rect 269328 453218 269370 453454
rect 269606 453218 269648 453454
rect 269328 453134 269648 453218
rect 269328 452898 269370 453134
rect 269606 452898 269648 453134
rect 269328 452866 269648 452898
rect 300048 453454 300368 453486
rect 300048 453218 300090 453454
rect 300326 453218 300368 453454
rect 300048 453134 300368 453218
rect 300048 452898 300090 453134
rect 300326 452898 300368 453134
rect 300048 452866 300368 452898
rect 330768 453454 331088 453486
rect 330768 453218 330810 453454
rect 331046 453218 331088 453454
rect 330768 453134 331088 453218
rect 330768 452898 330810 453134
rect 331046 452898 331088 453134
rect 330768 452866 331088 452898
rect 361488 453454 361808 453486
rect 361488 453218 361530 453454
rect 361766 453218 361808 453454
rect 361488 453134 361808 453218
rect 361488 452898 361530 453134
rect 361766 452898 361808 453134
rect 361488 452866 361808 452898
rect 392208 453454 392528 453486
rect 392208 453218 392250 453454
rect 392486 453218 392528 453454
rect 392208 453134 392528 453218
rect 392208 452898 392250 453134
rect 392486 452898 392528 453134
rect 392208 452866 392528 452898
rect 422928 453454 423248 453486
rect 422928 453218 422970 453454
rect 423206 453218 423248 453454
rect 422928 453134 423248 453218
rect 422928 452898 422970 453134
rect 423206 452898 423248 453134
rect 422928 452866 423248 452898
rect 453648 453454 453968 453486
rect 453648 453218 453690 453454
rect 453926 453218 453968 453454
rect 453648 453134 453968 453218
rect 453648 452898 453690 453134
rect 453926 452898 453968 453134
rect 453648 452866 453968 452898
rect 484368 453454 484688 453486
rect 484368 453218 484410 453454
rect 484646 453218 484688 453454
rect 484368 453134 484688 453218
rect 484368 452898 484410 453134
rect 484646 452898 484688 453134
rect 484368 452866 484688 452898
rect 515088 453454 515408 453486
rect 515088 453218 515130 453454
rect 515366 453218 515408 453454
rect 515088 453134 515408 453218
rect 515088 452898 515130 453134
rect 515366 452898 515408 453134
rect 515088 452866 515408 452898
rect 545808 453454 546128 453486
rect 545808 453218 545850 453454
rect 546086 453218 546128 453454
rect 545808 453134 546128 453218
rect 545808 452898 545850 453134
rect 546086 452898 546128 453134
rect 545808 452866 546128 452898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect 8208 435454 8528 435486
rect 8208 435218 8250 435454
rect 8486 435218 8528 435454
rect 8208 435134 8528 435218
rect 8208 434898 8250 435134
rect 8486 434898 8528 435134
rect 8208 434866 8528 434898
rect 38928 435454 39248 435486
rect 38928 435218 38970 435454
rect 39206 435218 39248 435454
rect 38928 435134 39248 435218
rect 38928 434898 38970 435134
rect 39206 434898 39248 435134
rect 38928 434866 39248 434898
rect 69648 435454 69968 435486
rect 69648 435218 69690 435454
rect 69926 435218 69968 435454
rect 69648 435134 69968 435218
rect 69648 434898 69690 435134
rect 69926 434898 69968 435134
rect 69648 434866 69968 434898
rect 100368 435454 100688 435486
rect 100368 435218 100410 435454
rect 100646 435218 100688 435454
rect 100368 435134 100688 435218
rect 100368 434898 100410 435134
rect 100646 434898 100688 435134
rect 100368 434866 100688 434898
rect 131088 435454 131408 435486
rect 131088 435218 131130 435454
rect 131366 435218 131408 435454
rect 131088 435134 131408 435218
rect 131088 434898 131130 435134
rect 131366 434898 131408 435134
rect 131088 434866 131408 434898
rect 161808 435454 162128 435486
rect 161808 435218 161850 435454
rect 162086 435218 162128 435454
rect 161808 435134 162128 435218
rect 161808 434898 161850 435134
rect 162086 434898 162128 435134
rect 161808 434866 162128 434898
rect 192528 435454 192848 435486
rect 192528 435218 192570 435454
rect 192806 435218 192848 435454
rect 192528 435134 192848 435218
rect 192528 434898 192570 435134
rect 192806 434898 192848 435134
rect 192528 434866 192848 434898
rect 223248 435454 223568 435486
rect 223248 435218 223290 435454
rect 223526 435218 223568 435454
rect 223248 435134 223568 435218
rect 223248 434898 223290 435134
rect 223526 434898 223568 435134
rect 223248 434866 223568 434898
rect 253968 435454 254288 435486
rect 253968 435218 254010 435454
rect 254246 435218 254288 435454
rect 253968 435134 254288 435218
rect 253968 434898 254010 435134
rect 254246 434898 254288 435134
rect 253968 434866 254288 434898
rect 284688 435454 285008 435486
rect 284688 435218 284730 435454
rect 284966 435218 285008 435454
rect 284688 435134 285008 435218
rect 284688 434898 284730 435134
rect 284966 434898 285008 435134
rect 284688 434866 285008 434898
rect 315408 435454 315728 435486
rect 315408 435218 315450 435454
rect 315686 435218 315728 435454
rect 315408 435134 315728 435218
rect 315408 434898 315450 435134
rect 315686 434898 315728 435134
rect 315408 434866 315728 434898
rect 346128 435454 346448 435486
rect 346128 435218 346170 435454
rect 346406 435218 346448 435454
rect 346128 435134 346448 435218
rect 346128 434898 346170 435134
rect 346406 434898 346448 435134
rect 346128 434866 346448 434898
rect 376848 435454 377168 435486
rect 376848 435218 376890 435454
rect 377126 435218 377168 435454
rect 376848 435134 377168 435218
rect 376848 434898 376890 435134
rect 377126 434898 377168 435134
rect 376848 434866 377168 434898
rect 407568 435454 407888 435486
rect 407568 435218 407610 435454
rect 407846 435218 407888 435454
rect 407568 435134 407888 435218
rect 407568 434898 407610 435134
rect 407846 434898 407888 435134
rect 407568 434866 407888 434898
rect 438288 435454 438608 435486
rect 438288 435218 438330 435454
rect 438566 435218 438608 435454
rect 438288 435134 438608 435218
rect 438288 434898 438330 435134
rect 438566 434898 438608 435134
rect 438288 434866 438608 434898
rect 469008 435454 469328 435486
rect 469008 435218 469050 435454
rect 469286 435218 469328 435454
rect 469008 435134 469328 435218
rect 469008 434898 469050 435134
rect 469286 434898 469328 435134
rect 469008 434866 469328 434898
rect 499728 435454 500048 435486
rect 499728 435218 499770 435454
rect 500006 435218 500048 435454
rect 499728 435134 500048 435218
rect 499728 434898 499770 435134
rect 500006 434898 500048 435134
rect 499728 434866 500048 434898
rect 530448 435454 530768 435486
rect 530448 435218 530490 435454
rect 530726 435218 530768 435454
rect 530448 435134 530768 435218
rect 530448 434898 530490 435134
rect 530726 434898 530768 435134
rect 530448 434866 530768 434898
rect 561168 435454 561488 435486
rect 561168 435218 561210 435454
rect 561446 435218 561488 435454
rect 561168 435134 561488 435218
rect 561168 434898 561210 435134
rect 561446 434898 561488 435134
rect 561168 434866 561488 434898
rect 567234 424894 567854 460338
rect 567234 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 567854 424894
rect 567234 424574 567854 424658
rect 567234 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 567854 424574
rect 23568 417454 23888 417486
rect 23568 417218 23610 417454
rect 23846 417218 23888 417454
rect 23568 417134 23888 417218
rect 23568 416898 23610 417134
rect 23846 416898 23888 417134
rect 23568 416866 23888 416898
rect 54288 417454 54608 417486
rect 54288 417218 54330 417454
rect 54566 417218 54608 417454
rect 54288 417134 54608 417218
rect 54288 416898 54330 417134
rect 54566 416898 54608 417134
rect 54288 416866 54608 416898
rect 85008 417454 85328 417486
rect 85008 417218 85050 417454
rect 85286 417218 85328 417454
rect 85008 417134 85328 417218
rect 85008 416898 85050 417134
rect 85286 416898 85328 417134
rect 85008 416866 85328 416898
rect 115728 417454 116048 417486
rect 115728 417218 115770 417454
rect 116006 417218 116048 417454
rect 115728 417134 116048 417218
rect 115728 416898 115770 417134
rect 116006 416898 116048 417134
rect 115728 416866 116048 416898
rect 146448 417454 146768 417486
rect 146448 417218 146490 417454
rect 146726 417218 146768 417454
rect 146448 417134 146768 417218
rect 146448 416898 146490 417134
rect 146726 416898 146768 417134
rect 146448 416866 146768 416898
rect 177168 417454 177488 417486
rect 177168 417218 177210 417454
rect 177446 417218 177488 417454
rect 177168 417134 177488 417218
rect 177168 416898 177210 417134
rect 177446 416898 177488 417134
rect 177168 416866 177488 416898
rect 207888 417454 208208 417486
rect 207888 417218 207930 417454
rect 208166 417218 208208 417454
rect 207888 417134 208208 417218
rect 207888 416898 207930 417134
rect 208166 416898 208208 417134
rect 207888 416866 208208 416898
rect 238608 417454 238928 417486
rect 238608 417218 238650 417454
rect 238886 417218 238928 417454
rect 238608 417134 238928 417218
rect 238608 416898 238650 417134
rect 238886 416898 238928 417134
rect 238608 416866 238928 416898
rect 269328 417454 269648 417486
rect 269328 417218 269370 417454
rect 269606 417218 269648 417454
rect 269328 417134 269648 417218
rect 269328 416898 269370 417134
rect 269606 416898 269648 417134
rect 269328 416866 269648 416898
rect 300048 417454 300368 417486
rect 300048 417218 300090 417454
rect 300326 417218 300368 417454
rect 300048 417134 300368 417218
rect 300048 416898 300090 417134
rect 300326 416898 300368 417134
rect 300048 416866 300368 416898
rect 330768 417454 331088 417486
rect 330768 417218 330810 417454
rect 331046 417218 331088 417454
rect 330768 417134 331088 417218
rect 330768 416898 330810 417134
rect 331046 416898 331088 417134
rect 330768 416866 331088 416898
rect 361488 417454 361808 417486
rect 361488 417218 361530 417454
rect 361766 417218 361808 417454
rect 361488 417134 361808 417218
rect 361488 416898 361530 417134
rect 361766 416898 361808 417134
rect 361488 416866 361808 416898
rect 392208 417454 392528 417486
rect 392208 417218 392250 417454
rect 392486 417218 392528 417454
rect 392208 417134 392528 417218
rect 392208 416898 392250 417134
rect 392486 416898 392528 417134
rect 392208 416866 392528 416898
rect 422928 417454 423248 417486
rect 422928 417218 422970 417454
rect 423206 417218 423248 417454
rect 422928 417134 423248 417218
rect 422928 416898 422970 417134
rect 423206 416898 423248 417134
rect 422928 416866 423248 416898
rect 453648 417454 453968 417486
rect 453648 417218 453690 417454
rect 453926 417218 453968 417454
rect 453648 417134 453968 417218
rect 453648 416898 453690 417134
rect 453926 416898 453968 417134
rect 453648 416866 453968 416898
rect 484368 417454 484688 417486
rect 484368 417218 484410 417454
rect 484646 417218 484688 417454
rect 484368 417134 484688 417218
rect 484368 416898 484410 417134
rect 484646 416898 484688 417134
rect 484368 416866 484688 416898
rect 515088 417454 515408 417486
rect 515088 417218 515130 417454
rect 515366 417218 515408 417454
rect 515088 417134 515408 417218
rect 515088 416898 515130 417134
rect 515366 416898 515408 417134
rect 515088 416866 515408 416898
rect 545808 417454 546128 417486
rect 545808 417218 545850 417454
rect 546086 417218 546128 417454
rect 545808 417134 546128 417218
rect 545808 416898 545850 417134
rect 546086 416898 546128 417134
rect 545808 416866 546128 416898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect 8208 399454 8528 399486
rect 8208 399218 8250 399454
rect 8486 399218 8528 399454
rect 8208 399134 8528 399218
rect 8208 398898 8250 399134
rect 8486 398898 8528 399134
rect 8208 398866 8528 398898
rect 38928 399454 39248 399486
rect 38928 399218 38970 399454
rect 39206 399218 39248 399454
rect 38928 399134 39248 399218
rect 38928 398898 38970 399134
rect 39206 398898 39248 399134
rect 38928 398866 39248 398898
rect 69648 399454 69968 399486
rect 69648 399218 69690 399454
rect 69926 399218 69968 399454
rect 69648 399134 69968 399218
rect 69648 398898 69690 399134
rect 69926 398898 69968 399134
rect 69648 398866 69968 398898
rect 100368 399454 100688 399486
rect 100368 399218 100410 399454
rect 100646 399218 100688 399454
rect 100368 399134 100688 399218
rect 100368 398898 100410 399134
rect 100646 398898 100688 399134
rect 100368 398866 100688 398898
rect 131088 399454 131408 399486
rect 131088 399218 131130 399454
rect 131366 399218 131408 399454
rect 131088 399134 131408 399218
rect 131088 398898 131130 399134
rect 131366 398898 131408 399134
rect 131088 398866 131408 398898
rect 161808 399454 162128 399486
rect 161808 399218 161850 399454
rect 162086 399218 162128 399454
rect 161808 399134 162128 399218
rect 161808 398898 161850 399134
rect 162086 398898 162128 399134
rect 161808 398866 162128 398898
rect 192528 399454 192848 399486
rect 192528 399218 192570 399454
rect 192806 399218 192848 399454
rect 192528 399134 192848 399218
rect 192528 398898 192570 399134
rect 192806 398898 192848 399134
rect 192528 398866 192848 398898
rect 223248 399454 223568 399486
rect 223248 399218 223290 399454
rect 223526 399218 223568 399454
rect 223248 399134 223568 399218
rect 223248 398898 223290 399134
rect 223526 398898 223568 399134
rect 223248 398866 223568 398898
rect 253968 399454 254288 399486
rect 253968 399218 254010 399454
rect 254246 399218 254288 399454
rect 253968 399134 254288 399218
rect 253968 398898 254010 399134
rect 254246 398898 254288 399134
rect 253968 398866 254288 398898
rect 284688 399454 285008 399486
rect 284688 399218 284730 399454
rect 284966 399218 285008 399454
rect 284688 399134 285008 399218
rect 284688 398898 284730 399134
rect 284966 398898 285008 399134
rect 284688 398866 285008 398898
rect 315408 399454 315728 399486
rect 315408 399218 315450 399454
rect 315686 399218 315728 399454
rect 315408 399134 315728 399218
rect 315408 398898 315450 399134
rect 315686 398898 315728 399134
rect 315408 398866 315728 398898
rect 346128 399454 346448 399486
rect 346128 399218 346170 399454
rect 346406 399218 346448 399454
rect 346128 399134 346448 399218
rect 346128 398898 346170 399134
rect 346406 398898 346448 399134
rect 346128 398866 346448 398898
rect 376848 399454 377168 399486
rect 376848 399218 376890 399454
rect 377126 399218 377168 399454
rect 376848 399134 377168 399218
rect 376848 398898 376890 399134
rect 377126 398898 377168 399134
rect 376848 398866 377168 398898
rect 407568 399454 407888 399486
rect 407568 399218 407610 399454
rect 407846 399218 407888 399454
rect 407568 399134 407888 399218
rect 407568 398898 407610 399134
rect 407846 398898 407888 399134
rect 407568 398866 407888 398898
rect 438288 399454 438608 399486
rect 438288 399218 438330 399454
rect 438566 399218 438608 399454
rect 438288 399134 438608 399218
rect 438288 398898 438330 399134
rect 438566 398898 438608 399134
rect 438288 398866 438608 398898
rect 469008 399454 469328 399486
rect 469008 399218 469050 399454
rect 469286 399218 469328 399454
rect 469008 399134 469328 399218
rect 469008 398898 469050 399134
rect 469286 398898 469328 399134
rect 469008 398866 469328 398898
rect 499728 399454 500048 399486
rect 499728 399218 499770 399454
rect 500006 399218 500048 399454
rect 499728 399134 500048 399218
rect 499728 398898 499770 399134
rect 500006 398898 500048 399134
rect 499728 398866 500048 398898
rect 530448 399454 530768 399486
rect 530448 399218 530490 399454
rect 530726 399218 530768 399454
rect 530448 399134 530768 399218
rect 530448 398898 530490 399134
rect 530726 398898 530768 399134
rect 530448 398866 530768 398898
rect 561168 399454 561488 399486
rect 561168 399218 561210 399454
rect 561446 399218 561488 399454
rect 561168 399134 561488 399218
rect 561168 398898 561210 399134
rect 561446 398898 561488 399134
rect 561168 398866 561488 398898
rect 567234 388894 567854 424338
rect 567234 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 567854 388894
rect 567234 388574 567854 388658
rect 567234 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 567854 388574
rect 23568 381454 23888 381486
rect 23568 381218 23610 381454
rect 23846 381218 23888 381454
rect 23568 381134 23888 381218
rect 23568 380898 23610 381134
rect 23846 380898 23888 381134
rect 23568 380866 23888 380898
rect 54288 381454 54608 381486
rect 54288 381218 54330 381454
rect 54566 381218 54608 381454
rect 54288 381134 54608 381218
rect 54288 380898 54330 381134
rect 54566 380898 54608 381134
rect 54288 380866 54608 380898
rect 85008 381454 85328 381486
rect 85008 381218 85050 381454
rect 85286 381218 85328 381454
rect 85008 381134 85328 381218
rect 85008 380898 85050 381134
rect 85286 380898 85328 381134
rect 85008 380866 85328 380898
rect 115728 381454 116048 381486
rect 115728 381218 115770 381454
rect 116006 381218 116048 381454
rect 115728 381134 116048 381218
rect 115728 380898 115770 381134
rect 116006 380898 116048 381134
rect 115728 380866 116048 380898
rect 146448 381454 146768 381486
rect 146448 381218 146490 381454
rect 146726 381218 146768 381454
rect 146448 381134 146768 381218
rect 146448 380898 146490 381134
rect 146726 380898 146768 381134
rect 146448 380866 146768 380898
rect 177168 381454 177488 381486
rect 177168 381218 177210 381454
rect 177446 381218 177488 381454
rect 177168 381134 177488 381218
rect 177168 380898 177210 381134
rect 177446 380898 177488 381134
rect 177168 380866 177488 380898
rect 207888 381454 208208 381486
rect 207888 381218 207930 381454
rect 208166 381218 208208 381454
rect 207888 381134 208208 381218
rect 207888 380898 207930 381134
rect 208166 380898 208208 381134
rect 207888 380866 208208 380898
rect 238608 381454 238928 381486
rect 238608 381218 238650 381454
rect 238886 381218 238928 381454
rect 238608 381134 238928 381218
rect 238608 380898 238650 381134
rect 238886 380898 238928 381134
rect 238608 380866 238928 380898
rect 269328 381454 269648 381486
rect 269328 381218 269370 381454
rect 269606 381218 269648 381454
rect 269328 381134 269648 381218
rect 269328 380898 269370 381134
rect 269606 380898 269648 381134
rect 269328 380866 269648 380898
rect 300048 381454 300368 381486
rect 300048 381218 300090 381454
rect 300326 381218 300368 381454
rect 300048 381134 300368 381218
rect 300048 380898 300090 381134
rect 300326 380898 300368 381134
rect 300048 380866 300368 380898
rect 330768 381454 331088 381486
rect 330768 381218 330810 381454
rect 331046 381218 331088 381454
rect 330768 381134 331088 381218
rect 330768 380898 330810 381134
rect 331046 380898 331088 381134
rect 330768 380866 331088 380898
rect 361488 381454 361808 381486
rect 361488 381218 361530 381454
rect 361766 381218 361808 381454
rect 361488 381134 361808 381218
rect 361488 380898 361530 381134
rect 361766 380898 361808 381134
rect 361488 380866 361808 380898
rect 392208 381454 392528 381486
rect 392208 381218 392250 381454
rect 392486 381218 392528 381454
rect 392208 381134 392528 381218
rect 392208 380898 392250 381134
rect 392486 380898 392528 381134
rect 392208 380866 392528 380898
rect 422928 381454 423248 381486
rect 422928 381218 422970 381454
rect 423206 381218 423248 381454
rect 422928 381134 423248 381218
rect 422928 380898 422970 381134
rect 423206 380898 423248 381134
rect 422928 380866 423248 380898
rect 453648 381454 453968 381486
rect 453648 381218 453690 381454
rect 453926 381218 453968 381454
rect 453648 381134 453968 381218
rect 453648 380898 453690 381134
rect 453926 380898 453968 381134
rect 453648 380866 453968 380898
rect 484368 381454 484688 381486
rect 484368 381218 484410 381454
rect 484646 381218 484688 381454
rect 484368 381134 484688 381218
rect 484368 380898 484410 381134
rect 484646 380898 484688 381134
rect 484368 380866 484688 380898
rect 515088 381454 515408 381486
rect 515088 381218 515130 381454
rect 515366 381218 515408 381454
rect 515088 381134 515408 381218
rect 515088 380898 515130 381134
rect 515366 380898 515408 381134
rect 515088 380866 515408 380898
rect 545808 381454 546128 381486
rect 545808 381218 545850 381454
rect 546086 381218 546128 381454
rect 545808 381134 546128 381218
rect 545808 380898 545850 381134
rect 546086 380898 546128 381134
rect 545808 380866 546128 380898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect 8208 363454 8528 363486
rect 8208 363218 8250 363454
rect 8486 363218 8528 363454
rect 8208 363134 8528 363218
rect 8208 362898 8250 363134
rect 8486 362898 8528 363134
rect 8208 362866 8528 362898
rect 38928 363454 39248 363486
rect 38928 363218 38970 363454
rect 39206 363218 39248 363454
rect 38928 363134 39248 363218
rect 38928 362898 38970 363134
rect 39206 362898 39248 363134
rect 38928 362866 39248 362898
rect 69648 363454 69968 363486
rect 69648 363218 69690 363454
rect 69926 363218 69968 363454
rect 69648 363134 69968 363218
rect 69648 362898 69690 363134
rect 69926 362898 69968 363134
rect 69648 362866 69968 362898
rect 100368 363454 100688 363486
rect 100368 363218 100410 363454
rect 100646 363218 100688 363454
rect 100368 363134 100688 363218
rect 100368 362898 100410 363134
rect 100646 362898 100688 363134
rect 100368 362866 100688 362898
rect 131088 363454 131408 363486
rect 131088 363218 131130 363454
rect 131366 363218 131408 363454
rect 131088 363134 131408 363218
rect 131088 362898 131130 363134
rect 131366 362898 131408 363134
rect 131088 362866 131408 362898
rect 161808 363454 162128 363486
rect 161808 363218 161850 363454
rect 162086 363218 162128 363454
rect 161808 363134 162128 363218
rect 161808 362898 161850 363134
rect 162086 362898 162128 363134
rect 161808 362866 162128 362898
rect 192528 363454 192848 363486
rect 192528 363218 192570 363454
rect 192806 363218 192848 363454
rect 192528 363134 192848 363218
rect 192528 362898 192570 363134
rect 192806 362898 192848 363134
rect 192528 362866 192848 362898
rect 223248 363454 223568 363486
rect 223248 363218 223290 363454
rect 223526 363218 223568 363454
rect 223248 363134 223568 363218
rect 223248 362898 223290 363134
rect 223526 362898 223568 363134
rect 223248 362866 223568 362898
rect 253968 363454 254288 363486
rect 253968 363218 254010 363454
rect 254246 363218 254288 363454
rect 253968 363134 254288 363218
rect 253968 362898 254010 363134
rect 254246 362898 254288 363134
rect 253968 362866 254288 362898
rect 284688 363454 285008 363486
rect 284688 363218 284730 363454
rect 284966 363218 285008 363454
rect 284688 363134 285008 363218
rect 284688 362898 284730 363134
rect 284966 362898 285008 363134
rect 284688 362866 285008 362898
rect 315408 363454 315728 363486
rect 315408 363218 315450 363454
rect 315686 363218 315728 363454
rect 315408 363134 315728 363218
rect 315408 362898 315450 363134
rect 315686 362898 315728 363134
rect 315408 362866 315728 362898
rect 346128 363454 346448 363486
rect 346128 363218 346170 363454
rect 346406 363218 346448 363454
rect 346128 363134 346448 363218
rect 346128 362898 346170 363134
rect 346406 362898 346448 363134
rect 346128 362866 346448 362898
rect 376848 363454 377168 363486
rect 376848 363218 376890 363454
rect 377126 363218 377168 363454
rect 376848 363134 377168 363218
rect 376848 362898 376890 363134
rect 377126 362898 377168 363134
rect 376848 362866 377168 362898
rect 407568 363454 407888 363486
rect 407568 363218 407610 363454
rect 407846 363218 407888 363454
rect 407568 363134 407888 363218
rect 407568 362898 407610 363134
rect 407846 362898 407888 363134
rect 407568 362866 407888 362898
rect 438288 363454 438608 363486
rect 438288 363218 438330 363454
rect 438566 363218 438608 363454
rect 438288 363134 438608 363218
rect 438288 362898 438330 363134
rect 438566 362898 438608 363134
rect 438288 362866 438608 362898
rect 469008 363454 469328 363486
rect 469008 363218 469050 363454
rect 469286 363218 469328 363454
rect 469008 363134 469328 363218
rect 469008 362898 469050 363134
rect 469286 362898 469328 363134
rect 469008 362866 469328 362898
rect 499728 363454 500048 363486
rect 499728 363218 499770 363454
rect 500006 363218 500048 363454
rect 499728 363134 500048 363218
rect 499728 362898 499770 363134
rect 500006 362898 500048 363134
rect 499728 362866 500048 362898
rect 530448 363454 530768 363486
rect 530448 363218 530490 363454
rect 530726 363218 530768 363454
rect 530448 363134 530768 363218
rect 530448 362898 530490 363134
rect 530726 362898 530768 363134
rect 530448 362866 530768 362898
rect 561168 363454 561488 363486
rect 561168 363218 561210 363454
rect 561446 363218 561488 363454
rect 561168 363134 561488 363218
rect 561168 362898 561210 363134
rect 561446 362898 561488 363134
rect 561168 362866 561488 362898
rect 567234 352894 567854 388338
rect 567234 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 567854 352894
rect 567234 352574 567854 352658
rect 567234 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 567854 352574
rect 23568 345454 23888 345486
rect 23568 345218 23610 345454
rect 23846 345218 23888 345454
rect 23568 345134 23888 345218
rect 23568 344898 23610 345134
rect 23846 344898 23888 345134
rect 23568 344866 23888 344898
rect 54288 345454 54608 345486
rect 54288 345218 54330 345454
rect 54566 345218 54608 345454
rect 54288 345134 54608 345218
rect 54288 344898 54330 345134
rect 54566 344898 54608 345134
rect 54288 344866 54608 344898
rect 85008 345454 85328 345486
rect 85008 345218 85050 345454
rect 85286 345218 85328 345454
rect 85008 345134 85328 345218
rect 85008 344898 85050 345134
rect 85286 344898 85328 345134
rect 85008 344866 85328 344898
rect 115728 345454 116048 345486
rect 115728 345218 115770 345454
rect 116006 345218 116048 345454
rect 115728 345134 116048 345218
rect 115728 344898 115770 345134
rect 116006 344898 116048 345134
rect 115728 344866 116048 344898
rect 146448 345454 146768 345486
rect 146448 345218 146490 345454
rect 146726 345218 146768 345454
rect 146448 345134 146768 345218
rect 146448 344898 146490 345134
rect 146726 344898 146768 345134
rect 146448 344866 146768 344898
rect 177168 345454 177488 345486
rect 177168 345218 177210 345454
rect 177446 345218 177488 345454
rect 177168 345134 177488 345218
rect 177168 344898 177210 345134
rect 177446 344898 177488 345134
rect 177168 344866 177488 344898
rect 207888 345454 208208 345486
rect 207888 345218 207930 345454
rect 208166 345218 208208 345454
rect 207888 345134 208208 345218
rect 207888 344898 207930 345134
rect 208166 344898 208208 345134
rect 207888 344866 208208 344898
rect 238608 345454 238928 345486
rect 238608 345218 238650 345454
rect 238886 345218 238928 345454
rect 238608 345134 238928 345218
rect 238608 344898 238650 345134
rect 238886 344898 238928 345134
rect 238608 344866 238928 344898
rect 269328 345454 269648 345486
rect 269328 345218 269370 345454
rect 269606 345218 269648 345454
rect 269328 345134 269648 345218
rect 269328 344898 269370 345134
rect 269606 344898 269648 345134
rect 269328 344866 269648 344898
rect 300048 345454 300368 345486
rect 300048 345218 300090 345454
rect 300326 345218 300368 345454
rect 300048 345134 300368 345218
rect 300048 344898 300090 345134
rect 300326 344898 300368 345134
rect 300048 344866 300368 344898
rect 330768 345454 331088 345486
rect 330768 345218 330810 345454
rect 331046 345218 331088 345454
rect 330768 345134 331088 345218
rect 330768 344898 330810 345134
rect 331046 344898 331088 345134
rect 330768 344866 331088 344898
rect 361488 345454 361808 345486
rect 361488 345218 361530 345454
rect 361766 345218 361808 345454
rect 361488 345134 361808 345218
rect 361488 344898 361530 345134
rect 361766 344898 361808 345134
rect 361488 344866 361808 344898
rect 392208 345454 392528 345486
rect 392208 345218 392250 345454
rect 392486 345218 392528 345454
rect 392208 345134 392528 345218
rect 392208 344898 392250 345134
rect 392486 344898 392528 345134
rect 392208 344866 392528 344898
rect 422928 345454 423248 345486
rect 422928 345218 422970 345454
rect 423206 345218 423248 345454
rect 422928 345134 423248 345218
rect 422928 344898 422970 345134
rect 423206 344898 423248 345134
rect 422928 344866 423248 344898
rect 453648 345454 453968 345486
rect 453648 345218 453690 345454
rect 453926 345218 453968 345454
rect 453648 345134 453968 345218
rect 453648 344898 453690 345134
rect 453926 344898 453968 345134
rect 453648 344866 453968 344898
rect 484368 345454 484688 345486
rect 484368 345218 484410 345454
rect 484646 345218 484688 345454
rect 484368 345134 484688 345218
rect 484368 344898 484410 345134
rect 484646 344898 484688 345134
rect 484368 344866 484688 344898
rect 515088 345454 515408 345486
rect 515088 345218 515130 345454
rect 515366 345218 515408 345454
rect 515088 345134 515408 345218
rect 515088 344898 515130 345134
rect 515366 344898 515408 345134
rect 515088 344866 515408 344898
rect 545808 345454 546128 345486
rect 545808 345218 545850 345454
rect 546086 345218 546128 345454
rect 545808 345134 546128 345218
rect 545808 344898 545850 345134
rect 546086 344898 546128 345134
rect 545808 344866 546128 344898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect 8208 327454 8528 327486
rect 8208 327218 8250 327454
rect 8486 327218 8528 327454
rect 8208 327134 8528 327218
rect 8208 326898 8250 327134
rect 8486 326898 8528 327134
rect 8208 326866 8528 326898
rect 38928 327454 39248 327486
rect 38928 327218 38970 327454
rect 39206 327218 39248 327454
rect 38928 327134 39248 327218
rect 38928 326898 38970 327134
rect 39206 326898 39248 327134
rect 38928 326866 39248 326898
rect 69648 327454 69968 327486
rect 69648 327218 69690 327454
rect 69926 327218 69968 327454
rect 69648 327134 69968 327218
rect 69648 326898 69690 327134
rect 69926 326898 69968 327134
rect 69648 326866 69968 326898
rect 100368 327454 100688 327486
rect 100368 327218 100410 327454
rect 100646 327218 100688 327454
rect 100368 327134 100688 327218
rect 100368 326898 100410 327134
rect 100646 326898 100688 327134
rect 100368 326866 100688 326898
rect 131088 327454 131408 327486
rect 131088 327218 131130 327454
rect 131366 327218 131408 327454
rect 131088 327134 131408 327218
rect 131088 326898 131130 327134
rect 131366 326898 131408 327134
rect 131088 326866 131408 326898
rect 161808 327454 162128 327486
rect 161808 327218 161850 327454
rect 162086 327218 162128 327454
rect 161808 327134 162128 327218
rect 161808 326898 161850 327134
rect 162086 326898 162128 327134
rect 161808 326866 162128 326898
rect 192528 327454 192848 327486
rect 192528 327218 192570 327454
rect 192806 327218 192848 327454
rect 192528 327134 192848 327218
rect 192528 326898 192570 327134
rect 192806 326898 192848 327134
rect 192528 326866 192848 326898
rect 223248 327454 223568 327486
rect 223248 327218 223290 327454
rect 223526 327218 223568 327454
rect 223248 327134 223568 327218
rect 223248 326898 223290 327134
rect 223526 326898 223568 327134
rect 223248 326866 223568 326898
rect 253968 327454 254288 327486
rect 253968 327218 254010 327454
rect 254246 327218 254288 327454
rect 253968 327134 254288 327218
rect 253968 326898 254010 327134
rect 254246 326898 254288 327134
rect 253968 326866 254288 326898
rect 284688 327454 285008 327486
rect 284688 327218 284730 327454
rect 284966 327218 285008 327454
rect 284688 327134 285008 327218
rect 284688 326898 284730 327134
rect 284966 326898 285008 327134
rect 284688 326866 285008 326898
rect 315408 327454 315728 327486
rect 315408 327218 315450 327454
rect 315686 327218 315728 327454
rect 315408 327134 315728 327218
rect 315408 326898 315450 327134
rect 315686 326898 315728 327134
rect 315408 326866 315728 326898
rect 346128 327454 346448 327486
rect 346128 327218 346170 327454
rect 346406 327218 346448 327454
rect 346128 327134 346448 327218
rect 346128 326898 346170 327134
rect 346406 326898 346448 327134
rect 346128 326866 346448 326898
rect 376848 327454 377168 327486
rect 376848 327218 376890 327454
rect 377126 327218 377168 327454
rect 376848 327134 377168 327218
rect 376848 326898 376890 327134
rect 377126 326898 377168 327134
rect 376848 326866 377168 326898
rect 407568 327454 407888 327486
rect 407568 327218 407610 327454
rect 407846 327218 407888 327454
rect 407568 327134 407888 327218
rect 407568 326898 407610 327134
rect 407846 326898 407888 327134
rect 407568 326866 407888 326898
rect 438288 327454 438608 327486
rect 438288 327218 438330 327454
rect 438566 327218 438608 327454
rect 438288 327134 438608 327218
rect 438288 326898 438330 327134
rect 438566 326898 438608 327134
rect 438288 326866 438608 326898
rect 469008 327454 469328 327486
rect 469008 327218 469050 327454
rect 469286 327218 469328 327454
rect 469008 327134 469328 327218
rect 469008 326898 469050 327134
rect 469286 326898 469328 327134
rect 469008 326866 469328 326898
rect 499728 327454 500048 327486
rect 499728 327218 499770 327454
rect 500006 327218 500048 327454
rect 499728 327134 500048 327218
rect 499728 326898 499770 327134
rect 500006 326898 500048 327134
rect 499728 326866 500048 326898
rect 530448 327454 530768 327486
rect 530448 327218 530490 327454
rect 530726 327218 530768 327454
rect 530448 327134 530768 327218
rect 530448 326898 530490 327134
rect 530726 326898 530768 327134
rect 530448 326866 530768 326898
rect 561168 327454 561488 327486
rect 561168 327218 561210 327454
rect 561446 327218 561488 327454
rect 561168 327134 561488 327218
rect 561168 326898 561210 327134
rect 561446 326898 561488 327134
rect 561168 326866 561488 326898
rect 567234 316894 567854 352338
rect 567234 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 567854 316894
rect 567234 316574 567854 316658
rect 567234 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 567854 316574
rect 23568 309454 23888 309486
rect 23568 309218 23610 309454
rect 23846 309218 23888 309454
rect 23568 309134 23888 309218
rect 23568 308898 23610 309134
rect 23846 308898 23888 309134
rect 23568 308866 23888 308898
rect 54288 309454 54608 309486
rect 54288 309218 54330 309454
rect 54566 309218 54608 309454
rect 54288 309134 54608 309218
rect 54288 308898 54330 309134
rect 54566 308898 54608 309134
rect 54288 308866 54608 308898
rect 85008 309454 85328 309486
rect 85008 309218 85050 309454
rect 85286 309218 85328 309454
rect 85008 309134 85328 309218
rect 85008 308898 85050 309134
rect 85286 308898 85328 309134
rect 85008 308866 85328 308898
rect 115728 309454 116048 309486
rect 115728 309218 115770 309454
rect 116006 309218 116048 309454
rect 115728 309134 116048 309218
rect 115728 308898 115770 309134
rect 116006 308898 116048 309134
rect 115728 308866 116048 308898
rect 146448 309454 146768 309486
rect 146448 309218 146490 309454
rect 146726 309218 146768 309454
rect 146448 309134 146768 309218
rect 146448 308898 146490 309134
rect 146726 308898 146768 309134
rect 146448 308866 146768 308898
rect 177168 309454 177488 309486
rect 177168 309218 177210 309454
rect 177446 309218 177488 309454
rect 177168 309134 177488 309218
rect 177168 308898 177210 309134
rect 177446 308898 177488 309134
rect 177168 308866 177488 308898
rect 207888 309454 208208 309486
rect 207888 309218 207930 309454
rect 208166 309218 208208 309454
rect 207888 309134 208208 309218
rect 207888 308898 207930 309134
rect 208166 308898 208208 309134
rect 207888 308866 208208 308898
rect 238608 309454 238928 309486
rect 238608 309218 238650 309454
rect 238886 309218 238928 309454
rect 238608 309134 238928 309218
rect 238608 308898 238650 309134
rect 238886 308898 238928 309134
rect 238608 308866 238928 308898
rect 269328 309454 269648 309486
rect 269328 309218 269370 309454
rect 269606 309218 269648 309454
rect 269328 309134 269648 309218
rect 269328 308898 269370 309134
rect 269606 308898 269648 309134
rect 269328 308866 269648 308898
rect 300048 309454 300368 309486
rect 300048 309218 300090 309454
rect 300326 309218 300368 309454
rect 300048 309134 300368 309218
rect 300048 308898 300090 309134
rect 300326 308898 300368 309134
rect 300048 308866 300368 308898
rect 330768 309454 331088 309486
rect 330768 309218 330810 309454
rect 331046 309218 331088 309454
rect 330768 309134 331088 309218
rect 330768 308898 330810 309134
rect 331046 308898 331088 309134
rect 330768 308866 331088 308898
rect 361488 309454 361808 309486
rect 361488 309218 361530 309454
rect 361766 309218 361808 309454
rect 361488 309134 361808 309218
rect 361488 308898 361530 309134
rect 361766 308898 361808 309134
rect 361488 308866 361808 308898
rect 392208 309454 392528 309486
rect 392208 309218 392250 309454
rect 392486 309218 392528 309454
rect 392208 309134 392528 309218
rect 392208 308898 392250 309134
rect 392486 308898 392528 309134
rect 392208 308866 392528 308898
rect 422928 309454 423248 309486
rect 422928 309218 422970 309454
rect 423206 309218 423248 309454
rect 422928 309134 423248 309218
rect 422928 308898 422970 309134
rect 423206 308898 423248 309134
rect 422928 308866 423248 308898
rect 453648 309454 453968 309486
rect 453648 309218 453690 309454
rect 453926 309218 453968 309454
rect 453648 309134 453968 309218
rect 453648 308898 453690 309134
rect 453926 308898 453968 309134
rect 453648 308866 453968 308898
rect 484368 309454 484688 309486
rect 484368 309218 484410 309454
rect 484646 309218 484688 309454
rect 484368 309134 484688 309218
rect 484368 308898 484410 309134
rect 484646 308898 484688 309134
rect 484368 308866 484688 308898
rect 515088 309454 515408 309486
rect 515088 309218 515130 309454
rect 515366 309218 515408 309454
rect 515088 309134 515408 309218
rect 515088 308898 515130 309134
rect 515366 308898 515408 309134
rect 515088 308866 515408 308898
rect 545808 309454 546128 309486
rect 545808 309218 545850 309454
rect 546086 309218 546128 309454
rect 545808 309134 546128 309218
rect 545808 308898 545850 309134
rect 546086 308898 546128 309134
rect 545808 308866 546128 308898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect 8208 291454 8528 291486
rect 8208 291218 8250 291454
rect 8486 291218 8528 291454
rect 8208 291134 8528 291218
rect 8208 290898 8250 291134
rect 8486 290898 8528 291134
rect 8208 290866 8528 290898
rect 38928 291454 39248 291486
rect 38928 291218 38970 291454
rect 39206 291218 39248 291454
rect 38928 291134 39248 291218
rect 38928 290898 38970 291134
rect 39206 290898 39248 291134
rect 38928 290866 39248 290898
rect 69648 291454 69968 291486
rect 69648 291218 69690 291454
rect 69926 291218 69968 291454
rect 69648 291134 69968 291218
rect 69648 290898 69690 291134
rect 69926 290898 69968 291134
rect 69648 290866 69968 290898
rect 100368 291454 100688 291486
rect 100368 291218 100410 291454
rect 100646 291218 100688 291454
rect 100368 291134 100688 291218
rect 100368 290898 100410 291134
rect 100646 290898 100688 291134
rect 100368 290866 100688 290898
rect 131088 291454 131408 291486
rect 131088 291218 131130 291454
rect 131366 291218 131408 291454
rect 131088 291134 131408 291218
rect 131088 290898 131130 291134
rect 131366 290898 131408 291134
rect 131088 290866 131408 290898
rect 161808 291454 162128 291486
rect 161808 291218 161850 291454
rect 162086 291218 162128 291454
rect 161808 291134 162128 291218
rect 161808 290898 161850 291134
rect 162086 290898 162128 291134
rect 161808 290866 162128 290898
rect 192528 291454 192848 291486
rect 192528 291218 192570 291454
rect 192806 291218 192848 291454
rect 192528 291134 192848 291218
rect 192528 290898 192570 291134
rect 192806 290898 192848 291134
rect 192528 290866 192848 290898
rect 223248 291454 223568 291486
rect 223248 291218 223290 291454
rect 223526 291218 223568 291454
rect 223248 291134 223568 291218
rect 223248 290898 223290 291134
rect 223526 290898 223568 291134
rect 223248 290866 223568 290898
rect 253968 291454 254288 291486
rect 253968 291218 254010 291454
rect 254246 291218 254288 291454
rect 253968 291134 254288 291218
rect 253968 290898 254010 291134
rect 254246 290898 254288 291134
rect 253968 290866 254288 290898
rect 284688 291454 285008 291486
rect 284688 291218 284730 291454
rect 284966 291218 285008 291454
rect 284688 291134 285008 291218
rect 284688 290898 284730 291134
rect 284966 290898 285008 291134
rect 284688 290866 285008 290898
rect 315408 291454 315728 291486
rect 315408 291218 315450 291454
rect 315686 291218 315728 291454
rect 315408 291134 315728 291218
rect 315408 290898 315450 291134
rect 315686 290898 315728 291134
rect 315408 290866 315728 290898
rect 346128 291454 346448 291486
rect 346128 291218 346170 291454
rect 346406 291218 346448 291454
rect 346128 291134 346448 291218
rect 346128 290898 346170 291134
rect 346406 290898 346448 291134
rect 346128 290866 346448 290898
rect 376848 291454 377168 291486
rect 376848 291218 376890 291454
rect 377126 291218 377168 291454
rect 376848 291134 377168 291218
rect 376848 290898 376890 291134
rect 377126 290898 377168 291134
rect 376848 290866 377168 290898
rect 407568 291454 407888 291486
rect 407568 291218 407610 291454
rect 407846 291218 407888 291454
rect 407568 291134 407888 291218
rect 407568 290898 407610 291134
rect 407846 290898 407888 291134
rect 407568 290866 407888 290898
rect 438288 291454 438608 291486
rect 438288 291218 438330 291454
rect 438566 291218 438608 291454
rect 438288 291134 438608 291218
rect 438288 290898 438330 291134
rect 438566 290898 438608 291134
rect 438288 290866 438608 290898
rect 469008 291454 469328 291486
rect 469008 291218 469050 291454
rect 469286 291218 469328 291454
rect 469008 291134 469328 291218
rect 469008 290898 469050 291134
rect 469286 290898 469328 291134
rect 469008 290866 469328 290898
rect 499728 291454 500048 291486
rect 499728 291218 499770 291454
rect 500006 291218 500048 291454
rect 499728 291134 500048 291218
rect 499728 290898 499770 291134
rect 500006 290898 500048 291134
rect 499728 290866 500048 290898
rect 530448 291454 530768 291486
rect 530448 291218 530490 291454
rect 530726 291218 530768 291454
rect 530448 291134 530768 291218
rect 530448 290898 530490 291134
rect 530726 290898 530768 291134
rect 530448 290866 530768 290898
rect 561168 291454 561488 291486
rect 561168 291218 561210 291454
rect 561446 291218 561488 291454
rect 561168 291134 561488 291218
rect 561168 290898 561210 291134
rect 561446 290898 561488 291134
rect 561168 290866 561488 290898
rect 567234 280894 567854 316338
rect 567234 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 567854 280894
rect 567234 280574 567854 280658
rect 567234 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 567854 280574
rect 23568 273454 23888 273486
rect 23568 273218 23610 273454
rect 23846 273218 23888 273454
rect 23568 273134 23888 273218
rect 23568 272898 23610 273134
rect 23846 272898 23888 273134
rect 23568 272866 23888 272898
rect 54288 273454 54608 273486
rect 54288 273218 54330 273454
rect 54566 273218 54608 273454
rect 54288 273134 54608 273218
rect 54288 272898 54330 273134
rect 54566 272898 54608 273134
rect 54288 272866 54608 272898
rect 85008 273454 85328 273486
rect 85008 273218 85050 273454
rect 85286 273218 85328 273454
rect 85008 273134 85328 273218
rect 85008 272898 85050 273134
rect 85286 272898 85328 273134
rect 85008 272866 85328 272898
rect 115728 273454 116048 273486
rect 115728 273218 115770 273454
rect 116006 273218 116048 273454
rect 115728 273134 116048 273218
rect 115728 272898 115770 273134
rect 116006 272898 116048 273134
rect 115728 272866 116048 272898
rect 146448 273454 146768 273486
rect 146448 273218 146490 273454
rect 146726 273218 146768 273454
rect 146448 273134 146768 273218
rect 146448 272898 146490 273134
rect 146726 272898 146768 273134
rect 146448 272866 146768 272898
rect 177168 273454 177488 273486
rect 177168 273218 177210 273454
rect 177446 273218 177488 273454
rect 177168 273134 177488 273218
rect 177168 272898 177210 273134
rect 177446 272898 177488 273134
rect 177168 272866 177488 272898
rect 207888 273454 208208 273486
rect 207888 273218 207930 273454
rect 208166 273218 208208 273454
rect 207888 273134 208208 273218
rect 207888 272898 207930 273134
rect 208166 272898 208208 273134
rect 207888 272866 208208 272898
rect 238608 273454 238928 273486
rect 238608 273218 238650 273454
rect 238886 273218 238928 273454
rect 238608 273134 238928 273218
rect 238608 272898 238650 273134
rect 238886 272898 238928 273134
rect 238608 272866 238928 272898
rect 269328 273454 269648 273486
rect 269328 273218 269370 273454
rect 269606 273218 269648 273454
rect 269328 273134 269648 273218
rect 269328 272898 269370 273134
rect 269606 272898 269648 273134
rect 269328 272866 269648 272898
rect 300048 273454 300368 273486
rect 300048 273218 300090 273454
rect 300326 273218 300368 273454
rect 300048 273134 300368 273218
rect 300048 272898 300090 273134
rect 300326 272898 300368 273134
rect 300048 272866 300368 272898
rect 330768 273454 331088 273486
rect 330768 273218 330810 273454
rect 331046 273218 331088 273454
rect 330768 273134 331088 273218
rect 330768 272898 330810 273134
rect 331046 272898 331088 273134
rect 330768 272866 331088 272898
rect 361488 273454 361808 273486
rect 361488 273218 361530 273454
rect 361766 273218 361808 273454
rect 361488 273134 361808 273218
rect 361488 272898 361530 273134
rect 361766 272898 361808 273134
rect 361488 272866 361808 272898
rect 392208 273454 392528 273486
rect 392208 273218 392250 273454
rect 392486 273218 392528 273454
rect 392208 273134 392528 273218
rect 392208 272898 392250 273134
rect 392486 272898 392528 273134
rect 392208 272866 392528 272898
rect 422928 273454 423248 273486
rect 422928 273218 422970 273454
rect 423206 273218 423248 273454
rect 422928 273134 423248 273218
rect 422928 272898 422970 273134
rect 423206 272898 423248 273134
rect 422928 272866 423248 272898
rect 453648 273454 453968 273486
rect 453648 273218 453690 273454
rect 453926 273218 453968 273454
rect 453648 273134 453968 273218
rect 453648 272898 453690 273134
rect 453926 272898 453968 273134
rect 453648 272866 453968 272898
rect 484368 273454 484688 273486
rect 484368 273218 484410 273454
rect 484646 273218 484688 273454
rect 484368 273134 484688 273218
rect 484368 272898 484410 273134
rect 484646 272898 484688 273134
rect 484368 272866 484688 272898
rect 515088 273454 515408 273486
rect 515088 273218 515130 273454
rect 515366 273218 515408 273454
rect 515088 273134 515408 273218
rect 515088 272898 515130 273134
rect 515366 272898 515408 273134
rect 515088 272866 515408 272898
rect 545808 273454 546128 273486
rect 545808 273218 545850 273454
rect 546086 273218 546128 273454
rect 545808 273134 546128 273218
rect 545808 272898 545850 273134
rect 546086 272898 546128 273134
rect 545808 272866 546128 272898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect 8208 255454 8528 255486
rect 8208 255218 8250 255454
rect 8486 255218 8528 255454
rect 8208 255134 8528 255218
rect 8208 254898 8250 255134
rect 8486 254898 8528 255134
rect 8208 254866 8528 254898
rect 38928 255454 39248 255486
rect 38928 255218 38970 255454
rect 39206 255218 39248 255454
rect 38928 255134 39248 255218
rect 38928 254898 38970 255134
rect 39206 254898 39248 255134
rect 38928 254866 39248 254898
rect 69648 255454 69968 255486
rect 69648 255218 69690 255454
rect 69926 255218 69968 255454
rect 69648 255134 69968 255218
rect 69648 254898 69690 255134
rect 69926 254898 69968 255134
rect 69648 254866 69968 254898
rect 100368 255454 100688 255486
rect 100368 255218 100410 255454
rect 100646 255218 100688 255454
rect 100368 255134 100688 255218
rect 100368 254898 100410 255134
rect 100646 254898 100688 255134
rect 100368 254866 100688 254898
rect 131088 255454 131408 255486
rect 131088 255218 131130 255454
rect 131366 255218 131408 255454
rect 131088 255134 131408 255218
rect 131088 254898 131130 255134
rect 131366 254898 131408 255134
rect 131088 254866 131408 254898
rect 161808 255454 162128 255486
rect 161808 255218 161850 255454
rect 162086 255218 162128 255454
rect 161808 255134 162128 255218
rect 161808 254898 161850 255134
rect 162086 254898 162128 255134
rect 161808 254866 162128 254898
rect 192528 255454 192848 255486
rect 192528 255218 192570 255454
rect 192806 255218 192848 255454
rect 192528 255134 192848 255218
rect 192528 254898 192570 255134
rect 192806 254898 192848 255134
rect 192528 254866 192848 254898
rect 223248 255454 223568 255486
rect 223248 255218 223290 255454
rect 223526 255218 223568 255454
rect 223248 255134 223568 255218
rect 223248 254898 223290 255134
rect 223526 254898 223568 255134
rect 223248 254866 223568 254898
rect 253968 255454 254288 255486
rect 253968 255218 254010 255454
rect 254246 255218 254288 255454
rect 253968 255134 254288 255218
rect 253968 254898 254010 255134
rect 254246 254898 254288 255134
rect 253968 254866 254288 254898
rect 284688 255454 285008 255486
rect 284688 255218 284730 255454
rect 284966 255218 285008 255454
rect 284688 255134 285008 255218
rect 284688 254898 284730 255134
rect 284966 254898 285008 255134
rect 284688 254866 285008 254898
rect 315408 255454 315728 255486
rect 315408 255218 315450 255454
rect 315686 255218 315728 255454
rect 315408 255134 315728 255218
rect 315408 254898 315450 255134
rect 315686 254898 315728 255134
rect 315408 254866 315728 254898
rect 346128 255454 346448 255486
rect 346128 255218 346170 255454
rect 346406 255218 346448 255454
rect 346128 255134 346448 255218
rect 346128 254898 346170 255134
rect 346406 254898 346448 255134
rect 346128 254866 346448 254898
rect 376848 255454 377168 255486
rect 376848 255218 376890 255454
rect 377126 255218 377168 255454
rect 376848 255134 377168 255218
rect 376848 254898 376890 255134
rect 377126 254898 377168 255134
rect 376848 254866 377168 254898
rect 407568 255454 407888 255486
rect 407568 255218 407610 255454
rect 407846 255218 407888 255454
rect 407568 255134 407888 255218
rect 407568 254898 407610 255134
rect 407846 254898 407888 255134
rect 407568 254866 407888 254898
rect 438288 255454 438608 255486
rect 438288 255218 438330 255454
rect 438566 255218 438608 255454
rect 438288 255134 438608 255218
rect 438288 254898 438330 255134
rect 438566 254898 438608 255134
rect 438288 254866 438608 254898
rect 469008 255454 469328 255486
rect 469008 255218 469050 255454
rect 469286 255218 469328 255454
rect 469008 255134 469328 255218
rect 469008 254898 469050 255134
rect 469286 254898 469328 255134
rect 469008 254866 469328 254898
rect 499728 255454 500048 255486
rect 499728 255218 499770 255454
rect 500006 255218 500048 255454
rect 499728 255134 500048 255218
rect 499728 254898 499770 255134
rect 500006 254898 500048 255134
rect 499728 254866 500048 254898
rect 530448 255454 530768 255486
rect 530448 255218 530490 255454
rect 530726 255218 530768 255454
rect 530448 255134 530768 255218
rect 530448 254898 530490 255134
rect 530726 254898 530768 255134
rect 530448 254866 530768 254898
rect 561168 255454 561488 255486
rect 561168 255218 561210 255454
rect 561446 255218 561488 255454
rect 561168 255134 561488 255218
rect 561168 254898 561210 255134
rect 561446 254898 561488 255134
rect 561168 254866 561488 254898
rect 567234 244894 567854 280338
rect 567234 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 567854 244894
rect 567234 244574 567854 244658
rect 567234 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 567854 244574
rect 23568 237454 23888 237486
rect 23568 237218 23610 237454
rect 23846 237218 23888 237454
rect 23568 237134 23888 237218
rect 23568 236898 23610 237134
rect 23846 236898 23888 237134
rect 23568 236866 23888 236898
rect 54288 237454 54608 237486
rect 54288 237218 54330 237454
rect 54566 237218 54608 237454
rect 54288 237134 54608 237218
rect 54288 236898 54330 237134
rect 54566 236898 54608 237134
rect 54288 236866 54608 236898
rect 85008 237454 85328 237486
rect 85008 237218 85050 237454
rect 85286 237218 85328 237454
rect 85008 237134 85328 237218
rect 85008 236898 85050 237134
rect 85286 236898 85328 237134
rect 85008 236866 85328 236898
rect 115728 237454 116048 237486
rect 115728 237218 115770 237454
rect 116006 237218 116048 237454
rect 115728 237134 116048 237218
rect 115728 236898 115770 237134
rect 116006 236898 116048 237134
rect 115728 236866 116048 236898
rect 146448 237454 146768 237486
rect 146448 237218 146490 237454
rect 146726 237218 146768 237454
rect 146448 237134 146768 237218
rect 146448 236898 146490 237134
rect 146726 236898 146768 237134
rect 146448 236866 146768 236898
rect 177168 237454 177488 237486
rect 177168 237218 177210 237454
rect 177446 237218 177488 237454
rect 177168 237134 177488 237218
rect 177168 236898 177210 237134
rect 177446 236898 177488 237134
rect 177168 236866 177488 236898
rect 207888 237454 208208 237486
rect 207888 237218 207930 237454
rect 208166 237218 208208 237454
rect 207888 237134 208208 237218
rect 207888 236898 207930 237134
rect 208166 236898 208208 237134
rect 207888 236866 208208 236898
rect 238608 237454 238928 237486
rect 238608 237218 238650 237454
rect 238886 237218 238928 237454
rect 238608 237134 238928 237218
rect 238608 236898 238650 237134
rect 238886 236898 238928 237134
rect 238608 236866 238928 236898
rect 269328 237454 269648 237486
rect 269328 237218 269370 237454
rect 269606 237218 269648 237454
rect 269328 237134 269648 237218
rect 269328 236898 269370 237134
rect 269606 236898 269648 237134
rect 269328 236866 269648 236898
rect 300048 237454 300368 237486
rect 300048 237218 300090 237454
rect 300326 237218 300368 237454
rect 300048 237134 300368 237218
rect 300048 236898 300090 237134
rect 300326 236898 300368 237134
rect 300048 236866 300368 236898
rect 330768 237454 331088 237486
rect 330768 237218 330810 237454
rect 331046 237218 331088 237454
rect 330768 237134 331088 237218
rect 330768 236898 330810 237134
rect 331046 236898 331088 237134
rect 330768 236866 331088 236898
rect 361488 237454 361808 237486
rect 361488 237218 361530 237454
rect 361766 237218 361808 237454
rect 361488 237134 361808 237218
rect 361488 236898 361530 237134
rect 361766 236898 361808 237134
rect 361488 236866 361808 236898
rect 392208 237454 392528 237486
rect 392208 237218 392250 237454
rect 392486 237218 392528 237454
rect 392208 237134 392528 237218
rect 392208 236898 392250 237134
rect 392486 236898 392528 237134
rect 392208 236866 392528 236898
rect 422928 237454 423248 237486
rect 422928 237218 422970 237454
rect 423206 237218 423248 237454
rect 422928 237134 423248 237218
rect 422928 236898 422970 237134
rect 423206 236898 423248 237134
rect 422928 236866 423248 236898
rect 453648 237454 453968 237486
rect 453648 237218 453690 237454
rect 453926 237218 453968 237454
rect 453648 237134 453968 237218
rect 453648 236898 453690 237134
rect 453926 236898 453968 237134
rect 453648 236866 453968 236898
rect 484368 237454 484688 237486
rect 484368 237218 484410 237454
rect 484646 237218 484688 237454
rect 484368 237134 484688 237218
rect 484368 236898 484410 237134
rect 484646 236898 484688 237134
rect 484368 236866 484688 236898
rect 515088 237454 515408 237486
rect 515088 237218 515130 237454
rect 515366 237218 515408 237454
rect 515088 237134 515408 237218
rect 515088 236898 515130 237134
rect 515366 236898 515408 237134
rect 515088 236866 515408 236898
rect 545808 237454 546128 237486
rect 545808 237218 545850 237454
rect 546086 237218 546128 237454
rect 545808 237134 546128 237218
rect 545808 236898 545850 237134
rect 546086 236898 546128 237134
rect 545808 236866 546128 236898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect 8208 219454 8528 219486
rect 8208 219218 8250 219454
rect 8486 219218 8528 219454
rect 8208 219134 8528 219218
rect 8208 218898 8250 219134
rect 8486 218898 8528 219134
rect 8208 218866 8528 218898
rect 38928 219454 39248 219486
rect 38928 219218 38970 219454
rect 39206 219218 39248 219454
rect 38928 219134 39248 219218
rect 38928 218898 38970 219134
rect 39206 218898 39248 219134
rect 38928 218866 39248 218898
rect 69648 219454 69968 219486
rect 69648 219218 69690 219454
rect 69926 219218 69968 219454
rect 69648 219134 69968 219218
rect 69648 218898 69690 219134
rect 69926 218898 69968 219134
rect 69648 218866 69968 218898
rect 100368 219454 100688 219486
rect 100368 219218 100410 219454
rect 100646 219218 100688 219454
rect 100368 219134 100688 219218
rect 100368 218898 100410 219134
rect 100646 218898 100688 219134
rect 100368 218866 100688 218898
rect 131088 219454 131408 219486
rect 131088 219218 131130 219454
rect 131366 219218 131408 219454
rect 131088 219134 131408 219218
rect 131088 218898 131130 219134
rect 131366 218898 131408 219134
rect 131088 218866 131408 218898
rect 161808 219454 162128 219486
rect 161808 219218 161850 219454
rect 162086 219218 162128 219454
rect 161808 219134 162128 219218
rect 161808 218898 161850 219134
rect 162086 218898 162128 219134
rect 161808 218866 162128 218898
rect 192528 219454 192848 219486
rect 192528 219218 192570 219454
rect 192806 219218 192848 219454
rect 192528 219134 192848 219218
rect 192528 218898 192570 219134
rect 192806 218898 192848 219134
rect 192528 218866 192848 218898
rect 223248 219454 223568 219486
rect 223248 219218 223290 219454
rect 223526 219218 223568 219454
rect 223248 219134 223568 219218
rect 223248 218898 223290 219134
rect 223526 218898 223568 219134
rect 223248 218866 223568 218898
rect 253968 219454 254288 219486
rect 253968 219218 254010 219454
rect 254246 219218 254288 219454
rect 253968 219134 254288 219218
rect 253968 218898 254010 219134
rect 254246 218898 254288 219134
rect 253968 218866 254288 218898
rect 284688 219454 285008 219486
rect 284688 219218 284730 219454
rect 284966 219218 285008 219454
rect 284688 219134 285008 219218
rect 284688 218898 284730 219134
rect 284966 218898 285008 219134
rect 284688 218866 285008 218898
rect 315408 219454 315728 219486
rect 315408 219218 315450 219454
rect 315686 219218 315728 219454
rect 315408 219134 315728 219218
rect 315408 218898 315450 219134
rect 315686 218898 315728 219134
rect 315408 218866 315728 218898
rect 346128 219454 346448 219486
rect 346128 219218 346170 219454
rect 346406 219218 346448 219454
rect 346128 219134 346448 219218
rect 346128 218898 346170 219134
rect 346406 218898 346448 219134
rect 346128 218866 346448 218898
rect 376848 219454 377168 219486
rect 376848 219218 376890 219454
rect 377126 219218 377168 219454
rect 376848 219134 377168 219218
rect 376848 218898 376890 219134
rect 377126 218898 377168 219134
rect 376848 218866 377168 218898
rect 407568 219454 407888 219486
rect 407568 219218 407610 219454
rect 407846 219218 407888 219454
rect 407568 219134 407888 219218
rect 407568 218898 407610 219134
rect 407846 218898 407888 219134
rect 407568 218866 407888 218898
rect 438288 219454 438608 219486
rect 438288 219218 438330 219454
rect 438566 219218 438608 219454
rect 438288 219134 438608 219218
rect 438288 218898 438330 219134
rect 438566 218898 438608 219134
rect 438288 218866 438608 218898
rect 469008 219454 469328 219486
rect 469008 219218 469050 219454
rect 469286 219218 469328 219454
rect 469008 219134 469328 219218
rect 469008 218898 469050 219134
rect 469286 218898 469328 219134
rect 469008 218866 469328 218898
rect 499728 219454 500048 219486
rect 499728 219218 499770 219454
rect 500006 219218 500048 219454
rect 499728 219134 500048 219218
rect 499728 218898 499770 219134
rect 500006 218898 500048 219134
rect 499728 218866 500048 218898
rect 530448 219454 530768 219486
rect 530448 219218 530490 219454
rect 530726 219218 530768 219454
rect 530448 219134 530768 219218
rect 530448 218898 530490 219134
rect 530726 218898 530768 219134
rect 530448 218866 530768 218898
rect 561168 219454 561488 219486
rect 561168 219218 561210 219454
rect 561446 219218 561488 219454
rect 561168 219134 561488 219218
rect 561168 218898 561210 219134
rect 561446 218898 561488 219134
rect 561168 218866 561488 218898
rect 567234 208894 567854 244338
rect 567234 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 567854 208894
rect 567234 208574 567854 208658
rect 567234 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 567854 208574
rect 23568 201454 23888 201486
rect 23568 201218 23610 201454
rect 23846 201218 23888 201454
rect 23568 201134 23888 201218
rect 23568 200898 23610 201134
rect 23846 200898 23888 201134
rect 23568 200866 23888 200898
rect 54288 201454 54608 201486
rect 54288 201218 54330 201454
rect 54566 201218 54608 201454
rect 54288 201134 54608 201218
rect 54288 200898 54330 201134
rect 54566 200898 54608 201134
rect 54288 200866 54608 200898
rect 85008 201454 85328 201486
rect 85008 201218 85050 201454
rect 85286 201218 85328 201454
rect 85008 201134 85328 201218
rect 85008 200898 85050 201134
rect 85286 200898 85328 201134
rect 85008 200866 85328 200898
rect 115728 201454 116048 201486
rect 115728 201218 115770 201454
rect 116006 201218 116048 201454
rect 115728 201134 116048 201218
rect 115728 200898 115770 201134
rect 116006 200898 116048 201134
rect 115728 200866 116048 200898
rect 146448 201454 146768 201486
rect 146448 201218 146490 201454
rect 146726 201218 146768 201454
rect 146448 201134 146768 201218
rect 146448 200898 146490 201134
rect 146726 200898 146768 201134
rect 146448 200866 146768 200898
rect 177168 201454 177488 201486
rect 177168 201218 177210 201454
rect 177446 201218 177488 201454
rect 177168 201134 177488 201218
rect 177168 200898 177210 201134
rect 177446 200898 177488 201134
rect 177168 200866 177488 200898
rect 207888 201454 208208 201486
rect 207888 201218 207930 201454
rect 208166 201218 208208 201454
rect 207888 201134 208208 201218
rect 207888 200898 207930 201134
rect 208166 200898 208208 201134
rect 207888 200866 208208 200898
rect 238608 201454 238928 201486
rect 238608 201218 238650 201454
rect 238886 201218 238928 201454
rect 238608 201134 238928 201218
rect 238608 200898 238650 201134
rect 238886 200898 238928 201134
rect 238608 200866 238928 200898
rect 269328 201454 269648 201486
rect 269328 201218 269370 201454
rect 269606 201218 269648 201454
rect 269328 201134 269648 201218
rect 269328 200898 269370 201134
rect 269606 200898 269648 201134
rect 269328 200866 269648 200898
rect 300048 201454 300368 201486
rect 300048 201218 300090 201454
rect 300326 201218 300368 201454
rect 300048 201134 300368 201218
rect 300048 200898 300090 201134
rect 300326 200898 300368 201134
rect 300048 200866 300368 200898
rect 330768 201454 331088 201486
rect 330768 201218 330810 201454
rect 331046 201218 331088 201454
rect 330768 201134 331088 201218
rect 330768 200898 330810 201134
rect 331046 200898 331088 201134
rect 330768 200866 331088 200898
rect 361488 201454 361808 201486
rect 361488 201218 361530 201454
rect 361766 201218 361808 201454
rect 361488 201134 361808 201218
rect 361488 200898 361530 201134
rect 361766 200898 361808 201134
rect 361488 200866 361808 200898
rect 392208 201454 392528 201486
rect 392208 201218 392250 201454
rect 392486 201218 392528 201454
rect 392208 201134 392528 201218
rect 392208 200898 392250 201134
rect 392486 200898 392528 201134
rect 392208 200866 392528 200898
rect 422928 201454 423248 201486
rect 422928 201218 422970 201454
rect 423206 201218 423248 201454
rect 422928 201134 423248 201218
rect 422928 200898 422970 201134
rect 423206 200898 423248 201134
rect 422928 200866 423248 200898
rect 453648 201454 453968 201486
rect 453648 201218 453690 201454
rect 453926 201218 453968 201454
rect 453648 201134 453968 201218
rect 453648 200898 453690 201134
rect 453926 200898 453968 201134
rect 453648 200866 453968 200898
rect 484368 201454 484688 201486
rect 484368 201218 484410 201454
rect 484646 201218 484688 201454
rect 484368 201134 484688 201218
rect 484368 200898 484410 201134
rect 484646 200898 484688 201134
rect 484368 200866 484688 200898
rect 515088 201454 515408 201486
rect 515088 201218 515130 201454
rect 515366 201218 515408 201454
rect 515088 201134 515408 201218
rect 515088 200898 515130 201134
rect 515366 200898 515408 201134
rect 515088 200866 515408 200898
rect 545808 201454 546128 201486
rect 545808 201218 545850 201454
rect 546086 201218 546128 201454
rect 545808 201134 546128 201218
rect 545808 200898 545850 201134
rect 546086 200898 546128 201134
rect 545808 200866 546128 200898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect 8208 183454 8528 183486
rect 8208 183218 8250 183454
rect 8486 183218 8528 183454
rect 8208 183134 8528 183218
rect 8208 182898 8250 183134
rect 8486 182898 8528 183134
rect 8208 182866 8528 182898
rect 38928 183454 39248 183486
rect 38928 183218 38970 183454
rect 39206 183218 39248 183454
rect 38928 183134 39248 183218
rect 38928 182898 38970 183134
rect 39206 182898 39248 183134
rect 38928 182866 39248 182898
rect 69648 183454 69968 183486
rect 69648 183218 69690 183454
rect 69926 183218 69968 183454
rect 69648 183134 69968 183218
rect 69648 182898 69690 183134
rect 69926 182898 69968 183134
rect 69648 182866 69968 182898
rect 100368 183454 100688 183486
rect 100368 183218 100410 183454
rect 100646 183218 100688 183454
rect 100368 183134 100688 183218
rect 100368 182898 100410 183134
rect 100646 182898 100688 183134
rect 100368 182866 100688 182898
rect 131088 183454 131408 183486
rect 131088 183218 131130 183454
rect 131366 183218 131408 183454
rect 131088 183134 131408 183218
rect 131088 182898 131130 183134
rect 131366 182898 131408 183134
rect 131088 182866 131408 182898
rect 161808 183454 162128 183486
rect 161808 183218 161850 183454
rect 162086 183218 162128 183454
rect 161808 183134 162128 183218
rect 161808 182898 161850 183134
rect 162086 182898 162128 183134
rect 161808 182866 162128 182898
rect 192528 183454 192848 183486
rect 192528 183218 192570 183454
rect 192806 183218 192848 183454
rect 192528 183134 192848 183218
rect 192528 182898 192570 183134
rect 192806 182898 192848 183134
rect 192528 182866 192848 182898
rect 223248 183454 223568 183486
rect 223248 183218 223290 183454
rect 223526 183218 223568 183454
rect 223248 183134 223568 183218
rect 223248 182898 223290 183134
rect 223526 182898 223568 183134
rect 223248 182866 223568 182898
rect 253968 183454 254288 183486
rect 253968 183218 254010 183454
rect 254246 183218 254288 183454
rect 253968 183134 254288 183218
rect 253968 182898 254010 183134
rect 254246 182898 254288 183134
rect 253968 182866 254288 182898
rect 284688 183454 285008 183486
rect 284688 183218 284730 183454
rect 284966 183218 285008 183454
rect 284688 183134 285008 183218
rect 284688 182898 284730 183134
rect 284966 182898 285008 183134
rect 284688 182866 285008 182898
rect 315408 183454 315728 183486
rect 315408 183218 315450 183454
rect 315686 183218 315728 183454
rect 315408 183134 315728 183218
rect 315408 182898 315450 183134
rect 315686 182898 315728 183134
rect 315408 182866 315728 182898
rect 346128 183454 346448 183486
rect 346128 183218 346170 183454
rect 346406 183218 346448 183454
rect 346128 183134 346448 183218
rect 346128 182898 346170 183134
rect 346406 182898 346448 183134
rect 346128 182866 346448 182898
rect 376848 183454 377168 183486
rect 376848 183218 376890 183454
rect 377126 183218 377168 183454
rect 376848 183134 377168 183218
rect 376848 182898 376890 183134
rect 377126 182898 377168 183134
rect 376848 182866 377168 182898
rect 407568 183454 407888 183486
rect 407568 183218 407610 183454
rect 407846 183218 407888 183454
rect 407568 183134 407888 183218
rect 407568 182898 407610 183134
rect 407846 182898 407888 183134
rect 407568 182866 407888 182898
rect 438288 183454 438608 183486
rect 438288 183218 438330 183454
rect 438566 183218 438608 183454
rect 438288 183134 438608 183218
rect 438288 182898 438330 183134
rect 438566 182898 438608 183134
rect 438288 182866 438608 182898
rect 469008 183454 469328 183486
rect 469008 183218 469050 183454
rect 469286 183218 469328 183454
rect 469008 183134 469328 183218
rect 469008 182898 469050 183134
rect 469286 182898 469328 183134
rect 469008 182866 469328 182898
rect 499728 183454 500048 183486
rect 499728 183218 499770 183454
rect 500006 183218 500048 183454
rect 499728 183134 500048 183218
rect 499728 182898 499770 183134
rect 500006 182898 500048 183134
rect 499728 182866 500048 182898
rect 530448 183454 530768 183486
rect 530448 183218 530490 183454
rect 530726 183218 530768 183454
rect 530448 183134 530768 183218
rect 530448 182898 530490 183134
rect 530726 182898 530768 183134
rect 530448 182866 530768 182898
rect 561168 183454 561488 183486
rect 561168 183218 561210 183454
rect 561446 183218 561488 183454
rect 561168 183134 561488 183218
rect 561168 182898 561210 183134
rect 561446 182898 561488 183134
rect 561168 182866 561488 182898
rect 567234 172894 567854 208338
rect 567234 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 567854 172894
rect 567234 172574 567854 172658
rect 567234 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 567854 172574
rect 23568 165454 23888 165486
rect 23568 165218 23610 165454
rect 23846 165218 23888 165454
rect 23568 165134 23888 165218
rect 23568 164898 23610 165134
rect 23846 164898 23888 165134
rect 23568 164866 23888 164898
rect 54288 165454 54608 165486
rect 54288 165218 54330 165454
rect 54566 165218 54608 165454
rect 54288 165134 54608 165218
rect 54288 164898 54330 165134
rect 54566 164898 54608 165134
rect 54288 164866 54608 164898
rect 85008 165454 85328 165486
rect 85008 165218 85050 165454
rect 85286 165218 85328 165454
rect 85008 165134 85328 165218
rect 85008 164898 85050 165134
rect 85286 164898 85328 165134
rect 85008 164866 85328 164898
rect 115728 165454 116048 165486
rect 115728 165218 115770 165454
rect 116006 165218 116048 165454
rect 115728 165134 116048 165218
rect 115728 164898 115770 165134
rect 116006 164898 116048 165134
rect 115728 164866 116048 164898
rect 146448 165454 146768 165486
rect 146448 165218 146490 165454
rect 146726 165218 146768 165454
rect 146448 165134 146768 165218
rect 146448 164898 146490 165134
rect 146726 164898 146768 165134
rect 146448 164866 146768 164898
rect 177168 165454 177488 165486
rect 177168 165218 177210 165454
rect 177446 165218 177488 165454
rect 177168 165134 177488 165218
rect 177168 164898 177210 165134
rect 177446 164898 177488 165134
rect 177168 164866 177488 164898
rect 207888 165454 208208 165486
rect 207888 165218 207930 165454
rect 208166 165218 208208 165454
rect 207888 165134 208208 165218
rect 207888 164898 207930 165134
rect 208166 164898 208208 165134
rect 207888 164866 208208 164898
rect 238608 165454 238928 165486
rect 238608 165218 238650 165454
rect 238886 165218 238928 165454
rect 238608 165134 238928 165218
rect 238608 164898 238650 165134
rect 238886 164898 238928 165134
rect 238608 164866 238928 164898
rect 269328 165454 269648 165486
rect 269328 165218 269370 165454
rect 269606 165218 269648 165454
rect 269328 165134 269648 165218
rect 269328 164898 269370 165134
rect 269606 164898 269648 165134
rect 269328 164866 269648 164898
rect 300048 165454 300368 165486
rect 300048 165218 300090 165454
rect 300326 165218 300368 165454
rect 300048 165134 300368 165218
rect 300048 164898 300090 165134
rect 300326 164898 300368 165134
rect 300048 164866 300368 164898
rect 330768 165454 331088 165486
rect 330768 165218 330810 165454
rect 331046 165218 331088 165454
rect 330768 165134 331088 165218
rect 330768 164898 330810 165134
rect 331046 164898 331088 165134
rect 330768 164866 331088 164898
rect 361488 165454 361808 165486
rect 361488 165218 361530 165454
rect 361766 165218 361808 165454
rect 361488 165134 361808 165218
rect 361488 164898 361530 165134
rect 361766 164898 361808 165134
rect 361488 164866 361808 164898
rect 392208 165454 392528 165486
rect 392208 165218 392250 165454
rect 392486 165218 392528 165454
rect 392208 165134 392528 165218
rect 392208 164898 392250 165134
rect 392486 164898 392528 165134
rect 392208 164866 392528 164898
rect 422928 165454 423248 165486
rect 422928 165218 422970 165454
rect 423206 165218 423248 165454
rect 422928 165134 423248 165218
rect 422928 164898 422970 165134
rect 423206 164898 423248 165134
rect 422928 164866 423248 164898
rect 453648 165454 453968 165486
rect 453648 165218 453690 165454
rect 453926 165218 453968 165454
rect 453648 165134 453968 165218
rect 453648 164898 453690 165134
rect 453926 164898 453968 165134
rect 453648 164866 453968 164898
rect 484368 165454 484688 165486
rect 484368 165218 484410 165454
rect 484646 165218 484688 165454
rect 484368 165134 484688 165218
rect 484368 164898 484410 165134
rect 484646 164898 484688 165134
rect 484368 164866 484688 164898
rect 515088 165454 515408 165486
rect 515088 165218 515130 165454
rect 515366 165218 515408 165454
rect 515088 165134 515408 165218
rect 515088 164898 515130 165134
rect 515366 164898 515408 165134
rect 515088 164866 515408 164898
rect 545808 165454 546128 165486
rect 545808 165218 545850 165454
rect 546086 165218 546128 165454
rect 545808 165134 546128 165218
rect 545808 164898 545850 165134
rect 546086 164898 546128 165134
rect 545808 164866 546128 164898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect 8208 147454 8528 147486
rect 8208 147218 8250 147454
rect 8486 147218 8528 147454
rect 8208 147134 8528 147218
rect 8208 146898 8250 147134
rect 8486 146898 8528 147134
rect 8208 146866 8528 146898
rect 38928 147454 39248 147486
rect 38928 147218 38970 147454
rect 39206 147218 39248 147454
rect 38928 147134 39248 147218
rect 38928 146898 38970 147134
rect 39206 146898 39248 147134
rect 38928 146866 39248 146898
rect 69648 147454 69968 147486
rect 69648 147218 69690 147454
rect 69926 147218 69968 147454
rect 69648 147134 69968 147218
rect 69648 146898 69690 147134
rect 69926 146898 69968 147134
rect 69648 146866 69968 146898
rect 100368 147454 100688 147486
rect 100368 147218 100410 147454
rect 100646 147218 100688 147454
rect 100368 147134 100688 147218
rect 100368 146898 100410 147134
rect 100646 146898 100688 147134
rect 100368 146866 100688 146898
rect 131088 147454 131408 147486
rect 131088 147218 131130 147454
rect 131366 147218 131408 147454
rect 131088 147134 131408 147218
rect 131088 146898 131130 147134
rect 131366 146898 131408 147134
rect 131088 146866 131408 146898
rect 161808 147454 162128 147486
rect 161808 147218 161850 147454
rect 162086 147218 162128 147454
rect 161808 147134 162128 147218
rect 161808 146898 161850 147134
rect 162086 146898 162128 147134
rect 161808 146866 162128 146898
rect 192528 147454 192848 147486
rect 192528 147218 192570 147454
rect 192806 147218 192848 147454
rect 192528 147134 192848 147218
rect 192528 146898 192570 147134
rect 192806 146898 192848 147134
rect 192528 146866 192848 146898
rect 223248 147454 223568 147486
rect 223248 147218 223290 147454
rect 223526 147218 223568 147454
rect 223248 147134 223568 147218
rect 223248 146898 223290 147134
rect 223526 146898 223568 147134
rect 223248 146866 223568 146898
rect 253968 147454 254288 147486
rect 253968 147218 254010 147454
rect 254246 147218 254288 147454
rect 253968 147134 254288 147218
rect 253968 146898 254010 147134
rect 254246 146898 254288 147134
rect 253968 146866 254288 146898
rect 284688 147454 285008 147486
rect 284688 147218 284730 147454
rect 284966 147218 285008 147454
rect 284688 147134 285008 147218
rect 284688 146898 284730 147134
rect 284966 146898 285008 147134
rect 284688 146866 285008 146898
rect 315408 147454 315728 147486
rect 315408 147218 315450 147454
rect 315686 147218 315728 147454
rect 315408 147134 315728 147218
rect 315408 146898 315450 147134
rect 315686 146898 315728 147134
rect 315408 146866 315728 146898
rect 346128 147454 346448 147486
rect 346128 147218 346170 147454
rect 346406 147218 346448 147454
rect 346128 147134 346448 147218
rect 346128 146898 346170 147134
rect 346406 146898 346448 147134
rect 346128 146866 346448 146898
rect 376848 147454 377168 147486
rect 376848 147218 376890 147454
rect 377126 147218 377168 147454
rect 376848 147134 377168 147218
rect 376848 146898 376890 147134
rect 377126 146898 377168 147134
rect 376848 146866 377168 146898
rect 407568 147454 407888 147486
rect 407568 147218 407610 147454
rect 407846 147218 407888 147454
rect 407568 147134 407888 147218
rect 407568 146898 407610 147134
rect 407846 146898 407888 147134
rect 407568 146866 407888 146898
rect 438288 147454 438608 147486
rect 438288 147218 438330 147454
rect 438566 147218 438608 147454
rect 438288 147134 438608 147218
rect 438288 146898 438330 147134
rect 438566 146898 438608 147134
rect 438288 146866 438608 146898
rect 469008 147454 469328 147486
rect 469008 147218 469050 147454
rect 469286 147218 469328 147454
rect 469008 147134 469328 147218
rect 469008 146898 469050 147134
rect 469286 146898 469328 147134
rect 469008 146866 469328 146898
rect 499728 147454 500048 147486
rect 499728 147218 499770 147454
rect 500006 147218 500048 147454
rect 499728 147134 500048 147218
rect 499728 146898 499770 147134
rect 500006 146898 500048 147134
rect 499728 146866 500048 146898
rect 530448 147454 530768 147486
rect 530448 147218 530490 147454
rect 530726 147218 530768 147454
rect 530448 147134 530768 147218
rect 530448 146898 530490 147134
rect 530726 146898 530768 147134
rect 530448 146866 530768 146898
rect 561168 147454 561488 147486
rect 561168 147218 561210 147454
rect 561446 147218 561488 147454
rect 561168 147134 561488 147218
rect 561168 146898 561210 147134
rect 561446 146898 561488 147134
rect 561168 146866 561488 146898
rect 567234 136894 567854 172338
rect 567234 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 567854 136894
rect 567234 136574 567854 136658
rect 567234 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 567854 136574
rect 23568 129454 23888 129486
rect 23568 129218 23610 129454
rect 23846 129218 23888 129454
rect 23568 129134 23888 129218
rect 23568 128898 23610 129134
rect 23846 128898 23888 129134
rect 23568 128866 23888 128898
rect 54288 129454 54608 129486
rect 54288 129218 54330 129454
rect 54566 129218 54608 129454
rect 54288 129134 54608 129218
rect 54288 128898 54330 129134
rect 54566 128898 54608 129134
rect 54288 128866 54608 128898
rect 85008 129454 85328 129486
rect 85008 129218 85050 129454
rect 85286 129218 85328 129454
rect 85008 129134 85328 129218
rect 85008 128898 85050 129134
rect 85286 128898 85328 129134
rect 85008 128866 85328 128898
rect 115728 129454 116048 129486
rect 115728 129218 115770 129454
rect 116006 129218 116048 129454
rect 115728 129134 116048 129218
rect 115728 128898 115770 129134
rect 116006 128898 116048 129134
rect 115728 128866 116048 128898
rect 146448 129454 146768 129486
rect 146448 129218 146490 129454
rect 146726 129218 146768 129454
rect 146448 129134 146768 129218
rect 146448 128898 146490 129134
rect 146726 128898 146768 129134
rect 146448 128866 146768 128898
rect 177168 129454 177488 129486
rect 177168 129218 177210 129454
rect 177446 129218 177488 129454
rect 177168 129134 177488 129218
rect 177168 128898 177210 129134
rect 177446 128898 177488 129134
rect 177168 128866 177488 128898
rect 207888 129454 208208 129486
rect 207888 129218 207930 129454
rect 208166 129218 208208 129454
rect 207888 129134 208208 129218
rect 207888 128898 207930 129134
rect 208166 128898 208208 129134
rect 207888 128866 208208 128898
rect 238608 129454 238928 129486
rect 238608 129218 238650 129454
rect 238886 129218 238928 129454
rect 238608 129134 238928 129218
rect 238608 128898 238650 129134
rect 238886 128898 238928 129134
rect 238608 128866 238928 128898
rect 269328 129454 269648 129486
rect 269328 129218 269370 129454
rect 269606 129218 269648 129454
rect 269328 129134 269648 129218
rect 269328 128898 269370 129134
rect 269606 128898 269648 129134
rect 269328 128866 269648 128898
rect 300048 129454 300368 129486
rect 300048 129218 300090 129454
rect 300326 129218 300368 129454
rect 300048 129134 300368 129218
rect 300048 128898 300090 129134
rect 300326 128898 300368 129134
rect 300048 128866 300368 128898
rect 330768 129454 331088 129486
rect 330768 129218 330810 129454
rect 331046 129218 331088 129454
rect 330768 129134 331088 129218
rect 330768 128898 330810 129134
rect 331046 128898 331088 129134
rect 330768 128866 331088 128898
rect 361488 129454 361808 129486
rect 361488 129218 361530 129454
rect 361766 129218 361808 129454
rect 361488 129134 361808 129218
rect 361488 128898 361530 129134
rect 361766 128898 361808 129134
rect 361488 128866 361808 128898
rect 392208 129454 392528 129486
rect 392208 129218 392250 129454
rect 392486 129218 392528 129454
rect 392208 129134 392528 129218
rect 392208 128898 392250 129134
rect 392486 128898 392528 129134
rect 392208 128866 392528 128898
rect 422928 129454 423248 129486
rect 422928 129218 422970 129454
rect 423206 129218 423248 129454
rect 422928 129134 423248 129218
rect 422928 128898 422970 129134
rect 423206 128898 423248 129134
rect 422928 128866 423248 128898
rect 453648 129454 453968 129486
rect 453648 129218 453690 129454
rect 453926 129218 453968 129454
rect 453648 129134 453968 129218
rect 453648 128898 453690 129134
rect 453926 128898 453968 129134
rect 453648 128866 453968 128898
rect 484368 129454 484688 129486
rect 484368 129218 484410 129454
rect 484646 129218 484688 129454
rect 484368 129134 484688 129218
rect 484368 128898 484410 129134
rect 484646 128898 484688 129134
rect 484368 128866 484688 128898
rect 515088 129454 515408 129486
rect 515088 129218 515130 129454
rect 515366 129218 515408 129454
rect 515088 129134 515408 129218
rect 515088 128898 515130 129134
rect 515366 128898 515408 129134
rect 515088 128866 515408 128898
rect 545808 129454 546128 129486
rect 545808 129218 545850 129454
rect 546086 129218 546128 129454
rect 545808 129134 546128 129218
rect 545808 128898 545850 129134
rect 546086 128898 546128 129134
rect 545808 128866 546128 128898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect 8208 111454 8528 111486
rect 8208 111218 8250 111454
rect 8486 111218 8528 111454
rect 8208 111134 8528 111218
rect 8208 110898 8250 111134
rect 8486 110898 8528 111134
rect 8208 110866 8528 110898
rect 38928 111454 39248 111486
rect 38928 111218 38970 111454
rect 39206 111218 39248 111454
rect 38928 111134 39248 111218
rect 38928 110898 38970 111134
rect 39206 110898 39248 111134
rect 38928 110866 39248 110898
rect 69648 111454 69968 111486
rect 69648 111218 69690 111454
rect 69926 111218 69968 111454
rect 69648 111134 69968 111218
rect 69648 110898 69690 111134
rect 69926 110898 69968 111134
rect 69648 110866 69968 110898
rect 100368 111454 100688 111486
rect 100368 111218 100410 111454
rect 100646 111218 100688 111454
rect 100368 111134 100688 111218
rect 100368 110898 100410 111134
rect 100646 110898 100688 111134
rect 100368 110866 100688 110898
rect 131088 111454 131408 111486
rect 131088 111218 131130 111454
rect 131366 111218 131408 111454
rect 131088 111134 131408 111218
rect 131088 110898 131130 111134
rect 131366 110898 131408 111134
rect 131088 110866 131408 110898
rect 161808 111454 162128 111486
rect 161808 111218 161850 111454
rect 162086 111218 162128 111454
rect 161808 111134 162128 111218
rect 161808 110898 161850 111134
rect 162086 110898 162128 111134
rect 161808 110866 162128 110898
rect 192528 111454 192848 111486
rect 192528 111218 192570 111454
rect 192806 111218 192848 111454
rect 192528 111134 192848 111218
rect 192528 110898 192570 111134
rect 192806 110898 192848 111134
rect 192528 110866 192848 110898
rect 223248 111454 223568 111486
rect 223248 111218 223290 111454
rect 223526 111218 223568 111454
rect 223248 111134 223568 111218
rect 223248 110898 223290 111134
rect 223526 110898 223568 111134
rect 223248 110866 223568 110898
rect 253968 111454 254288 111486
rect 253968 111218 254010 111454
rect 254246 111218 254288 111454
rect 253968 111134 254288 111218
rect 253968 110898 254010 111134
rect 254246 110898 254288 111134
rect 253968 110866 254288 110898
rect 284688 111454 285008 111486
rect 284688 111218 284730 111454
rect 284966 111218 285008 111454
rect 284688 111134 285008 111218
rect 284688 110898 284730 111134
rect 284966 110898 285008 111134
rect 284688 110866 285008 110898
rect 315408 111454 315728 111486
rect 315408 111218 315450 111454
rect 315686 111218 315728 111454
rect 315408 111134 315728 111218
rect 315408 110898 315450 111134
rect 315686 110898 315728 111134
rect 315408 110866 315728 110898
rect 346128 111454 346448 111486
rect 346128 111218 346170 111454
rect 346406 111218 346448 111454
rect 346128 111134 346448 111218
rect 346128 110898 346170 111134
rect 346406 110898 346448 111134
rect 346128 110866 346448 110898
rect 376848 111454 377168 111486
rect 376848 111218 376890 111454
rect 377126 111218 377168 111454
rect 376848 111134 377168 111218
rect 376848 110898 376890 111134
rect 377126 110898 377168 111134
rect 376848 110866 377168 110898
rect 407568 111454 407888 111486
rect 407568 111218 407610 111454
rect 407846 111218 407888 111454
rect 407568 111134 407888 111218
rect 407568 110898 407610 111134
rect 407846 110898 407888 111134
rect 407568 110866 407888 110898
rect 438288 111454 438608 111486
rect 438288 111218 438330 111454
rect 438566 111218 438608 111454
rect 438288 111134 438608 111218
rect 438288 110898 438330 111134
rect 438566 110898 438608 111134
rect 438288 110866 438608 110898
rect 469008 111454 469328 111486
rect 469008 111218 469050 111454
rect 469286 111218 469328 111454
rect 469008 111134 469328 111218
rect 469008 110898 469050 111134
rect 469286 110898 469328 111134
rect 469008 110866 469328 110898
rect 499728 111454 500048 111486
rect 499728 111218 499770 111454
rect 500006 111218 500048 111454
rect 499728 111134 500048 111218
rect 499728 110898 499770 111134
rect 500006 110898 500048 111134
rect 499728 110866 500048 110898
rect 530448 111454 530768 111486
rect 530448 111218 530490 111454
rect 530726 111218 530768 111454
rect 530448 111134 530768 111218
rect 530448 110898 530490 111134
rect 530726 110898 530768 111134
rect 530448 110866 530768 110898
rect 561168 111454 561488 111486
rect 561168 111218 561210 111454
rect 561446 111218 561488 111454
rect 561168 111134 561488 111218
rect 561168 110898 561210 111134
rect 561446 110898 561488 111134
rect 561168 110866 561488 110898
rect 567234 100894 567854 136338
rect 567234 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 567854 100894
rect 567234 100574 567854 100658
rect 567234 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 567854 100574
rect 23568 93454 23888 93486
rect 23568 93218 23610 93454
rect 23846 93218 23888 93454
rect 23568 93134 23888 93218
rect 23568 92898 23610 93134
rect 23846 92898 23888 93134
rect 23568 92866 23888 92898
rect 54288 93454 54608 93486
rect 54288 93218 54330 93454
rect 54566 93218 54608 93454
rect 54288 93134 54608 93218
rect 54288 92898 54330 93134
rect 54566 92898 54608 93134
rect 54288 92866 54608 92898
rect 85008 93454 85328 93486
rect 85008 93218 85050 93454
rect 85286 93218 85328 93454
rect 85008 93134 85328 93218
rect 85008 92898 85050 93134
rect 85286 92898 85328 93134
rect 85008 92866 85328 92898
rect 115728 93454 116048 93486
rect 115728 93218 115770 93454
rect 116006 93218 116048 93454
rect 115728 93134 116048 93218
rect 115728 92898 115770 93134
rect 116006 92898 116048 93134
rect 115728 92866 116048 92898
rect 146448 93454 146768 93486
rect 146448 93218 146490 93454
rect 146726 93218 146768 93454
rect 146448 93134 146768 93218
rect 146448 92898 146490 93134
rect 146726 92898 146768 93134
rect 146448 92866 146768 92898
rect 177168 93454 177488 93486
rect 177168 93218 177210 93454
rect 177446 93218 177488 93454
rect 177168 93134 177488 93218
rect 177168 92898 177210 93134
rect 177446 92898 177488 93134
rect 177168 92866 177488 92898
rect 207888 93454 208208 93486
rect 207888 93218 207930 93454
rect 208166 93218 208208 93454
rect 207888 93134 208208 93218
rect 207888 92898 207930 93134
rect 208166 92898 208208 93134
rect 207888 92866 208208 92898
rect 238608 93454 238928 93486
rect 238608 93218 238650 93454
rect 238886 93218 238928 93454
rect 238608 93134 238928 93218
rect 238608 92898 238650 93134
rect 238886 92898 238928 93134
rect 238608 92866 238928 92898
rect 269328 93454 269648 93486
rect 269328 93218 269370 93454
rect 269606 93218 269648 93454
rect 269328 93134 269648 93218
rect 269328 92898 269370 93134
rect 269606 92898 269648 93134
rect 269328 92866 269648 92898
rect 300048 93454 300368 93486
rect 300048 93218 300090 93454
rect 300326 93218 300368 93454
rect 300048 93134 300368 93218
rect 300048 92898 300090 93134
rect 300326 92898 300368 93134
rect 300048 92866 300368 92898
rect 330768 93454 331088 93486
rect 330768 93218 330810 93454
rect 331046 93218 331088 93454
rect 330768 93134 331088 93218
rect 330768 92898 330810 93134
rect 331046 92898 331088 93134
rect 330768 92866 331088 92898
rect 361488 93454 361808 93486
rect 361488 93218 361530 93454
rect 361766 93218 361808 93454
rect 361488 93134 361808 93218
rect 361488 92898 361530 93134
rect 361766 92898 361808 93134
rect 361488 92866 361808 92898
rect 392208 93454 392528 93486
rect 392208 93218 392250 93454
rect 392486 93218 392528 93454
rect 392208 93134 392528 93218
rect 392208 92898 392250 93134
rect 392486 92898 392528 93134
rect 392208 92866 392528 92898
rect 422928 93454 423248 93486
rect 422928 93218 422970 93454
rect 423206 93218 423248 93454
rect 422928 93134 423248 93218
rect 422928 92898 422970 93134
rect 423206 92898 423248 93134
rect 422928 92866 423248 92898
rect 453648 93454 453968 93486
rect 453648 93218 453690 93454
rect 453926 93218 453968 93454
rect 453648 93134 453968 93218
rect 453648 92898 453690 93134
rect 453926 92898 453968 93134
rect 453648 92866 453968 92898
rect 484368 93454 484688 93486
rect 484368 93218 484410 93454
rect 484646 93218 484688 93454
rect 484368 93134 484688 93218
rect 484368 92898 484410 93134
rect 484646 92898 484688 93134
rect 484368 92866 484688 92898
rect 515088 93454 515408 93486
rect 515088 93218 515130 93454
rect 515366 93218 515408 93454
rect 515088 93134 515408 93218
rect 515088 92898 515130 93134
rect 515366 92898 515408 93134
rect 515088 92866 515408 92898
rect 545808 93454 546128 93486
rect 545808 93218 545850 93454
rect 546086 93218 546128 93454
rect 545808 93134 546128 93218
rect 545808 92898 545850 93134
rect 546086 92898 546128 93134
rect 545808 92866 546128 92898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect 8208 75454 8528 75486
rect 8208 75218 8250 75454
rect 8486 75218 8528 75454
rect 8208 75134 8528 75218
rect 8208 74898 8250 75134
rect 8486 74898 8528 75134
rect 8208 74866 8528 74898
rect 38928 75454 39248 75486
rect 38928 75218 38970 75454
rect 39206 75218 39248 75454
rect 38928 75134 39248 75218
rect 38928 74898 38970 75134
rect 39206 74898 39248 75134
rect 38928 74866 39248 74898
rect 69648 75454 69968 75486
rect 69648 75218 69690 75454
rect 69926 75218 69968 75454
rect 69648 75134 69968 75218
rect 69648 74898 69690 75134
rect 69926 74898 69968 75134
rect 69648 74866 69968 74898
rect 100368 75454 100688 75486
rect 100368 75218 100410 75454
rect 100646 75218 100688 75454
rect 100368 75134 100688 75218
rect 100368 74898 100410 75134
rect 100646 74898 100688 75134
rect 100368 74866 100688 74898
rect 131088 75454 131408 75486
rect 131088 75218 131130 75454
rect 131366 75218 131408 75454
rect 131088 75134 131408 75218
rect 131088 74898 131130 75134
rect 131366 74898 131408 75134
rect 131088 74866 131408 74898
rect 161808 75454 162128 75486
rect 161808 75218 161850 75454
rect 162086 75218 162128 75454
rect 161808 75134 162128 75218
rect 161808 74898 161850 75134
rect 162086 74898 162128 75134
rect 161808 74866 162128 74898
rect 192528 75454 192848 75486
rect 192528 75218 192570 75454
rect 192806 75218 192848 75454
rect 192528 75134 192848 75218
rect 192528 74898 192570 75134
rect 192806 74898 192848 75134
rect 192528 74866 192848 74898
rect 223248 75454 223568 75486
rect 223248 75218 223290 75454
rect 223526 75218 223568 75454
rect 223248 75134 223568 75218
rect 223248 74898 223290 75134
rect 223526 74898 223568 75134
rect 223248 74866 223568 74898
rect 253968 75454 254288 75486
rect 253968 75218 254010 75454
rect 254246 75218 254288 75454
rect 253968 75134 254288 75218
rect 253968 74898 254010 75134
rect 254246 74898 254288 75134
rect 253968 74866 254288 74898
rect 284688 75454 285008 75486
rect 284688 75218 284730 75454
rect 284966 75218 285008 75454
rect 284688 75134 285008 75218
rect 284688 74898 284730 75134
rect 284966 74898 285008 75134
rect 284688 74866 285008 74898
rect 315408 75454 315728 75486
rect 315408 75218 315450 75454
rect 315686 75218 315728 75454
rect 315408 75134 315728 75218
rect 315408 74898 315450 75134
rect 315686 74898 315728 75134
rect 315408 74866 315728 74898
rect 346128 75454 346448 75486
rect 346128 75218 346170 75454
rect 346406 75218 346448 75454
rect 346128 75134 346448 75218
rect 346128 74898 346170 75134
rect 346406 74898 346448 75134
rect 346128 74866 346448 74898
rect 376848 75454 377168 75486
rect 376848 75218 376890 75454
rect 377126 75218 377168 75454
rect 376848 75134 377168 75218
rect 376848 74898 376890 75134
rect 377126 74898 377168 75134
rect 376848 74866 377168 74898
rect 407568 75454 407888 75486
rect 407568 75218 407610 75454
rect 407846 75218 407888 75454
rect 407568 75134 407888 75218
rect 407568 74898 407610 75134
rect 407846 74898 407888 75134
rect 407568 74866 407888 74898
rect 438288 75454 438608 75486
rect 438288 75218 438330 75454
rect 438566 75218 438608 75454
rect 438288 75134 438608 75218
rect 438288 74898 438330 75134
rect 438566 74898 438608 75134
rect 438288 74866 438608 74898
rect 469008 75454 469328 75486
rect 469008 75218 469050 75454
rect 469286 75218 469328 75454
rect 469008 75134 469328 75218
rect 469008 74898 469050 75134
rect 469286 74898 469328 75134
rect 469008 74866 469328 74898
rect 499728 75454 500048 75486
rect 499728 75218 499770 75454
rect 500006 75218 500048 75454
rect 499728 75134 500048 75218
rect 499728 74898 499770 75134
rect 500006 74898 500048 75134
rect 499728 74866 500048 74898
rect 530448 75454 530768 75486
rect 530448 75218 530490 75454
rect 530726 75218 530768 75454
rect 530448 75134 530768 75218
rect 530448 74898 530490 75134
rect 530726 74898 530768 75134
rect 530448 74866 530768 74898
rect 561168 75454 561488 75486
rect 561168 75218 561210 75454
rect 561446 75218 561488 75454
rect 561168 75134 561488 75218
rect 561168 74898 561210 75134
rect 561446 74898 561488 75134
rect 561168 74866 561488 74898
rect 567234 64894 567854 100338
rect 567234 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 567854 64894
rect 567234 64574 567854 64658
rect 567234 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 567854 64574
rect 23568 57454 23888 57486
rect 23568 57218 23610 57454
rect 23846 57218 23888 57454
rect 23568 57134 23888 57218
rect 23568 56898 23610 57134
rect 23846 56898 23888 57134
rect 23568 56866 23888 56898
rect 54288 57454 54608 57486
rect 54288 57218 54330 57454
rect 54566 57218 54608 57454
rect 54288 57134 54608 57218
rect 54288 56898 54330 57134
rect 54566 56898 54608 57134
rect 54288 56866 54608 56898
rect 85008 57454 85328 57486
rect 85008 57218 85050 57454
rect 85286 57218 85328 57454
rect 85008 57134 85328 57218
rect 85008 56898 85050 57134
rect 85286 56898 85328 57134
rect 85008 56866 85328 56898
rect 115728 57454 116048 57486
rect 115728 57218 115770 57454
rect 116006 57218 116048 57454
rect 115728 57134 116048 57218
rect 115728 56898 115770 57134
rect 116006 56898 116048 57134
rect 115728 56866 116048 56898
rect 146448 57454 146768 57486
rect 146448 57218 146490 57454
rect 146726 57218 146768 57454
rect 146448 57134 146768 57218
rect 146448 56898 146490 57134
rect 146726 56898 146768 57134
rect 146448 56866 146768 56898
rect 177168 57454 177488 57486
rect 177168 57218 177210 57454
rect 177446 57218 177488 57454
rect 177168 57134 177488 57218
rect 177168 56898 177210 57134
rect 177446 56898 177488 57134
rect 177168 56866 177488 56898
rect 207888 57454 208208 57486
rect 207888 57218 207930 57454
rect 208166 57218 208208 57454
rect 207888 57134 208208 57218
rect 207888 56898 207930 57134
rect 208166 56898 208208 57134
rect 207888 56866 208208 56898
rect 238608 57454 238928 57486
rect 238608 57218 238650 57454
rect 238886 57218 238928 57454
rect 238608 57134 238928 57218
rect 238608 56898 238650 57134
rect 238886 56898 238928 57134
rect 238608 56866 238928 56898
rect 269328 57454 269648 57486
rect 269328 57218 269370 57454
rect 269606 57218 269648 57454
rect 269328 57134 269648 57218
rect 269328 56898 269370 57134
rect 269606 56898 269648 57134
rect 269328 56866 269648 56898
rect 300048 57454 300368 57486
rect 300048 57218 300090 57454
rect 300326 57218 300368 57454
rect 300048 57134 300368 57218
rect 300048 56898 300090 57134
rect 300326 56898 300368 57134
rect 300048 56866 300368 56898
rect 330768 57454 331088 57486
rect 330768 57218 330810 57454
rect 331046 57218 331088 57454
rect 330768 57134 331088 57218
rect 330768 56898 330810 57134
rect 331046 56898 331088 57134
rect 330768 56866 331088 56898
rect 361488 57454 361808 57486
rect 361488 57218 361530 57454
rect 361766 57218 361808 57454
rect 361488 57134 361808 57218
rect 361488 56898 361530 57134
rect 361766 56898 361808 57134
rect 361488 56866 361808 56898
rect 392208 57454 392528 57486
rect 392208 57218 392250 57454
rect 392486 57218 392528 57454
rect 392208 57134 392528 57218
rect 392208 56898 392250 57134
rect 392486 56898 392528 57134
rect 392208 56866 392528 56898
rect 422928 57454 423248 57486
rect 422928 57218 422970 57454
rect 423206 57218 423248 57454
rect 422928 57134 423248 57218
rect 422928 56898 422970 57134
rect 423206 56898 423248 57134
rect 422928 56866 423248 56898
rect 453648 57454 453968 57486
rect 453648 57218 453690 57454
rect 453926 57218 453968 57454
rect 453648 57134 453968 57218
rect 453648 56898 453690 57134
rect 453926 56898 453968 57134
rect 453648 56866 453968 56898
rect 484368 57454 484688 57486
rect 484368 57218 484410 57454
rect 484646 57218 484688 57454
rect 484368 57134 484688 57218
rect 484368 56898 484410 57134
rect 484646 56898 484688 57134
rect 484368 56866 484688 56898
rect 515088 57454 515408 57486
rect 515088 57218 515130 57454
rect 515366 57218 515408 57454
rect 515088 57134 515408 57218
rect 515088 56898 515130 57134
rect 515366 56898 515408 57134
rect 515088 56866 515408 56898
rect 545808 57454 546128 57486
rect 545808 57218 545850 57454
rect 546086 57218 546128 57454
rect 545808 57134 546128 57218
rect 545808 56898 545850 57134
rect 546086 56898 546128 57134
rect 545808 56866 546128 56898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect 8208 39454 8528 39486
rect 8208 39218 8250 39454
rect 8486 39218 8528 39454
rect 8208 39134 8528 39218
rect 8208 38898 8250 39134
rect 8486 38898 8528 39134
rect 8208 38866 8528 38898
rect 38928 39454 39248 39486
rect 38928 39218 38970 39454
rect 39206 39218 39248 39454
rect 38928 39134 39248 39218
rect 38928 38898 38970 39134
rect 39206 38898 39248 39134
rect 38928 38866 39248 38898
rect 69648 39454 69968 39486
rect 69648 39218 69690 39454
rect 69926 39218 69968 39454
rect 69648 39134 69968 39218
rect 69648 38898 69690 39134
rect 69926 38898 69968 39134
rect 69648 38866 69968 38898
rect 100368 39454 100688 39486
rect 100368 39218 100410 39454
rect 100646 39218 100688 39454
rect 100368 39134 100688 39218
rect 100368 38898 100410 39134
rect 100646 38898 100688 39134
rect 100368 38866 100688 38898
rect 131088 39454 131408 39486
rect 131088 39218 131130 39454
rect 131366 39218 131408 39454
rect 131088 39134 131408 39218
rect 131088 38898 131130 39134
rect 131366 38898 131408 39134
rect 131088 38866 131408 38898
rect 161808 39454 162128 39486
rect 161808 39218 161850 39454
rect 162086 39218 162128 39454
rect 161808 39134 162128 39218
rect 161808 38898 161850 39134
rect 162086 38898 162128 39134
rect 161808 38866 162128 38898
rect 192528 39454 192848 39486
rect 192528 39218 192570 39454
rect 192806 39218 192848 39454
rect 192528 39134 192848 39218
rect 192528 38898 192570 39134
rect 192806 38898 192848 39134
rect 192528 38866 192848 38898
rect 223248 39454 223568 39486
rect 223248 39218 223290 39454
rect 223526 39218 223568 39454
rect 223248 39134 223568 39218
rect 223248 38898 223290 39134
rect 223526 38898 223568 39134
rect 223248 38866 223568 38898
rect 253968 39454 254288 39486
rect 253968 39218 254010 39454
rect 254246 39218 254288 39454
rect 253968 39134 254288 39218
rect 253968 38898 254010 39134
rect 254246 38898 254288 39134
rect 253968 38866 254288 38898
rect 284688 39454 285008 39486
rect 284688 39218 284730 39454
rect 284966 39218 285008 39454
rect 284688 39134 285008 39218
rect 284688 38898 284730 39134
rect 284966 38898 285008 39134
rect 284688 38866 285008 38898
rect 315408 39454 315728 39486
rect 315408 39218 315450 39454
rect 315686 39218 315728 39454
rect 315408 39134 315728 39218
rect 315408 38898 315450 39134
rect 315686 38898 315728 39134
rect 315408 38866 315728 38898
rect 346128 39454 346448 39486
rect 346128 39218 346170 39454
rect 346406 39218 346448 39454
rect 346128 39134 346448 39218
rect 346128 38898 346170 39134
rect 346406 38898 346448 39134
rect 346128 38866 346448 38898
rect 376848 39454 377168 39486
rect 376848 39218 376890 39454
rect 377126 39218 377168 39454
rect 376848 39134 377168 39218
rect 376848 38898 376890 39134
rect 377126 38898 377168 39134
rect 376848 38866 377168 38898
rect 407568 39454 407888 39486
rect 407568 39218 407610 39454
rect 407846 39218 407888 39454
rect 407568 39134 407888 39218
rect 407568 38898 407610 39134
rect 407846 38898 407888 39134
rect 407568 38866 407888 38898
rect 438288 39454 438608 39486
rect 438288 39218 438330 39454
rect 438566 39218 438608 39454
rect 438288 39134 438608 39218
rect 438288 38898 438330 39134
rect 438566 38898 438608 39134
rect 438288 38866 438608 38898
rect 469008 39454 469328 39486
rect 469008 39218 469050 39454
rect 469286 39218 469328 39454
rect 469008 39134 469328 39218
rect 469008 38898 469050 39134
rect 469286 38898 469328 39134
rect 469008 38866 469328 38898
rect 499728 39454 500048 39486
rect 499728 39218 499770 39454
rect 500006 39218 500048 39454
rect 499728 39134 500048 39218
rect 499728 38898 499770 39134
rect 500006 38898 500048 39134
rect 499728 38866 500048 38898
rect 530448 39454 530768 39486
rect 530448 39218 530490 39454
rect 530726 39218 530768 39454
rect 530448 39134 530768 39218
rect 530448 38898 530490 39134
rect 530726 38898 530768 39134
rect 530448 38866 530768 38898
rect 561168 39454 561488 39486
rect 561168 39218 561210 39454
rect 561446 39218 561488 39454
rect 561168 39134 561488 39218
rect 561168 38898 561210 39134
rect 561446 38898 561488 39134
rect 561168 38866 561488 38898
rect 567234 28894 567854 64338
rect 567234 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 567854 28894
rect 567234 28574 567854 28658
rect 567234 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 567854 28574
rect 23568 21454 23888 21486
rect 23568 21218 23610 21454
rect 23846 21218 23888 21454
rect 23568 21134 23888 21218
rect 23568 20898 23610 21134
rect 23846 20898 23888 21134
rect 23568 20866 23888 20898
rect 54288 21454 54608 21486
rect 54288 21218 54330 21454
rect 54566 21218 54608 21454
rect 54288 21134 54608 21218
rect 54288 20898 54330 21134
rect 54566 20898 54608 21134
rect 54288 20866 54608 20898
rect 85008 21454 85328 21486
rect 85008 21218 85050 21454
rect 85286 21218 85328 21454
rect 85008 21134 85328 21218
rect 85008 20898 85050 21134
rect 85286 20898 85328 21134
rect 85008 20866 85328 20898
rect 115728 21454 116048 21486
rect 115728 21218 115770 21454
rect 116006 21218 116048 21454
rect 115728 21134 116048 21218
rect 115728 20898 115770 21134
rect 116006 20898 116048 21134
rect 115728 20866 116048 20898
rect 146448 21454 146768 21486
rect 146448 21218 146490 21454
rect 146726 21218 146768 21454
rect 146448 21134 146768 21218
rect 146448 20898 146490 21134
rect 146726 20898 146768 21134
rect 146448 20866 146768 20898
rect 177168 21454 177488 21486
rect 177168 21218 177210 21454
rect 177446 21218 177488 21454
rect 177168 21134 177488 21218
rect 177168 20898 177210 21134
rect 177446 20898 177488 21134
rect 177168 20866 177488 20898
rect 207888 21454 208208 21486
rect 207888 21218 207930 21454
rect 208166 21218 208208 21454
rect 207888 21134 208208 21218
rect 207888 20898 207930 21134
rect 208166 20898 208208 21134
rect 207888 20866 208208 20898
rect 238608 21454 238928 21486
rect 238608 21218 238650 21454
rect 238886 21218 238928 21454
rect 238608 21134 238928 21218
rect 238608 20898 238650 21134
rect 238886 20898 238928 21134
rect 238608 20866 238928 20898
rect 269328 21454 269648 21486
rect 269328 21218 269370 21454
rect 269606 21218 269648 21454
rect 269328 21134 269648 21218
rect 269328 20898 269370 21134
rect 269606 20898 269648 21134
rect 269328 20866 269648 20898
rect 300048 21454 300368 21486
rect 300048 21218 300090 21454
rect 300326 21218 300368 21454
rect 300048 21134 300368 21218
rect 300048 20898 300090 21134
rect 300326 20898 300368 21134
rect 300048 20866 300368 20898
rect 330768 21454 331088 21486
rect 330768 21218 330810 21454
rect 331046 21218 331088 21454
rect 330768 21134 331088 21218
rect 330768 20898 330810 21134
rect 331046 20898 331088 21134
rect 330768 20866 331088 20898
rect 361488 21454 361808 21486
rect 361488 21218 361530 21454
rect 361766 21218 361808 21454
rect 361488 21134 361808 21218
rect 361488 20898 361530 21134
rect 361766 20898 361808 21134
rect 361488 20866 361808 20898
rect 392208 21454 392528 21486
rect 392208 21218 392250 21454
rect 392486 21218 392528 21454
rect 392208 21134 392528 21218
rect 392208 20898 392250 21134
rect 392486 20898 392528 21134
rect 392208 20866 392528 20898
rect 422928 21454 423248 21486
rect 422928 21218 422970 21454
rect 423206 21218 423248 21454
rect 422928 21134 423248 21218
rect 422928 20898 422970 21134
rect 423206 20898 423248 21134
rect 422928 20866 423248 20898
rect 453648 21454 453968 21486
rect 453648 21218 453690 21454
rect 453926 21218 453968 21454
rect 453648 21134 453968 21218
rect 453648 20898 453690 21134
rect 453926 20898 453968 21134
rect 453648 20866 453968 20898
rect 484368 21454 484688 21486
rect 484368 21218 484410 21454
rect 484646 21218 484688 21454
rect 484368 21134 484688 21218
rect 484368 20898 484410 21134
rect 484646 20898 484688 21134
rect 484368 20866 484688 20898
rect 515088 21454 515408 21486
rect 515088 21218 515130 21454
rect 515366 21218 515408 21454
rect 515088 21134 515408 21218
rect 515088 20898 515130 21134
rect 515366 20898 515408 21134
rect 515088 20866 515408 20898
rect 545808 21454 546128 21486
rect 545808 21218 545850 21454
rect 546086 21218 546128 21454
rect 545808 21134 546128 21218
rect 545808 20898 545850 21134
rect 546086 20898 546128 21134
rect 545808 20866 546128 20898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect 8208 3454 8528 3486
rect 8208 3218 8250 3454
rect 8486 3218 8528 3454
rect 8208 3134 8528 3218
rect 8208 2898 8250 3134
rect 8486 2898 8528 3134
rect 8208 2866 8528 2898
rect 38928 3454 39248 3486
rect 38928 3218 38970 3454
rect 39206 3218 39248 3454
rect 38928 3134 39248 3218
rect 38928 2898 38970 3134
rect 39206 2898 39248 3134
rect 38928 2866 39248 2898
rect 69648 3454 69968 3486
rect 69648 3218 69690 3454
rect 69926 3218 69968 3454
rect 69648 3134 69968 3218
rect 69648 2898 69690 3134
rect 69926 2898 69968 3134
rect 69648 2866 69968 2898
rect 100368 3454 100688 3486
rect 100368 3218 100410 3454
rect 100646 3218 100688 3454
rect 100368 3134 100688 3218
rect 100368 2898 100410 3134
rect 100646 2898 100688 3134
rect 100368 2866 100688 2898
rect 131088 3454 131408 3486
rect 131088 3218 131130 3454
rect 131366 3218 131408 3454
rect 131088 3134 131408 3218
rect 131088 2898 131130 3134
rect 131366 2898 131408 3134
rect 131088 2866 131408 2898
rect 161808 3454 162128 3486
rect 161808 3218 161850 3454
rect 162086 3218 162128 3454
rect 161808 3134 162128 3218
rect 161808 2898 161850 3134
rect 162086 2898 162128 3134
rect 161808 2866 162128 2898
rect 192528 3454 192848 3486
rect 192528 3218 192570 3454
rect 192806 3218 192848 3454
rect 192528 3134 192848 3218
rect 192528 2898 192570 3134
rect 192806 2898 192848 3134
rect 192528 2866 192848 2898
rect 223248 3454 223568 3486
rect 223248 3218 223290 3454
rect 223526 3218 223568 3454
rect 223248 3134 223568 3218
rect 223248 2898 223290 3134
rect 223526 2898 223568 3134
rect 223248 2866 223568 2898
rect 253968 3454 254288 3486
rect 253968 3218 254010 3454
rect 254246 3218 254288 3454
rect 253968 3134 254288 3218
rect 253968 2898 254010 3134
rect 254246 2898 254288 3134
rect 253968 2866 254288 2898
rect 284688 3454 285008 3486
rect 284688 3218 284730 3454
rect 284966 3218 285008 3454
rect 284688 3134 285008 3218
rect 284688 2898 284730 3134
rect 284966 2898 285008 3134
rect 284688 2866 285008 2898
rect 315408 3454 315728 3486
rect 315408 3218 315450 3454
rect 315686 3218 315728 3454
rect 315408 3134 315728 3218
rect 315408 2898 315450 3134
rect 315686 2898 315728 3134
rect 315408 2866 315728 2898
rect 346128 3454 346448 3486
rect 346128 3218 346170 3454
rect 346406 3218 346448 3454
rect 346128 3134 346448 3218
rect 346128 2898 346170 3134
rect 346406 2898 346448 3134
rect 346128 2866 346448 2898
rect 376848 3454 377168 3486
rect 376848 3218 376890 3454
rect 377126 3218 377168 3454
rect 376848 3134 377168 3218
rect 376848 2898 376890 3134
rect 377126 2898 377168 3134
rect 376848 2866 377168 2898
rect 407568 3454 407888 3486
rect 407568 3218 407610 3454
rect 407846 3218 407888 3454
rect 407568 3134 407888 3218
rect 407568 2898 407610 3134
rect 407846 2898 407888 3134
rect 407568 2866 407888 2898
rect 438288 3454 438608 3486
rect 438288 3218 438330 3454
rect 438566 3218 438608 3454
rect 438288 3134 438608 3218
rect 438288 2898 438330 3134
rect 438566 2898 438608 3134
rect 438288 2866 438608 2898
rect 469008 3454 469328 3486
rect 469008 3218 469050 3454
rect 469286 3218 469328 3454
rect 469008 3134 469328 3218
rect 469008 2898 469050 3134
rect 469286 2898 469328 3134
rect 469008 2866 469328 2898
rect 499728 3454 500048 3486
rect 499728 3218 499770 3454
rect 500006 3218 500048 3454
rect 499728 3134 500048 3218
rect 499728 2898 499770 3134
rect 500006 2898 500048 3134
rect 499728 2866 500048 2898
rect 530448 3454 530768 3486
rect 530448 3218 530490 3454
rect 530726 3218 530768 3454
rect 530448 3134 530768 3218
rect 530448 2898 530490 3134
rect 530726 2898 530768 3134
rect 530448 2866 530768 2898
rect 561168 3454 561488 3486
rect 561168 3218 561210 3454
rect 561446 3218 561488 3454
rect 561168 3134 561488 3218
rect 561168 2898 561210 3134
rect 561446 2898 561488 3134
rect 561168 2866 561488 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 -2000
rect 5514 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 6134 -2266
rect 5514 -2586 6134 -2502
rect 5514 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 6134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 -2000
rect 9234 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 9854 -4186
rect 9234 -4506 9854 -4422
rect 9234 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 9854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 -2000
rect 23514 -3226 24134 -2000
rect 23514 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 24134 -3226
rect 23514 -3546 24134 -3462
rect 23514 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 24134 -3546
rect 23514 -3814 24134 -3782
rect 27234 -5146 27854 -2000
rect 27234 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 27854 -5146
rect 27234 -5466 27854 -5382
rect 27234 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 27854 -5466
rect 27234 -5734 27854 -5702
rect 12954 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 13574 -6106
rect 12954 -6426 13574 -6342
rect 12954 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 13574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 -2000
rect 41514 -2266 42134 -2000
rect 41514 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 42134 -2266
rect 41514 -2586 42134 -2502
rect 41514 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 42134 -2586
rect 41514 -3814 42134 -2822
rect 45234 -4186 45854 -2000
rect 45234 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 45854 -4186
rect 45234 -4506 45854 -4422
rect 45234 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 45854 -4506
rect 45234 -5734 45854 -4742
rect 30954 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 31574 -7066
rect 30954 -7386 31574 -7302
rect 30954 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 31574 -7386
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 -2000
rect 59514 -3226 60134 -2000
rect 59514 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 60134 -3226
rect 59514 -3546 60134 -3462
rect 59514 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 60134 -3546
rect 59514 -3814 60134 -3782
rect 63234 -5146 63854 -2000
rect 63234 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 63854 -5146
rect 63234 -5466 63854 -5382
rect 63234 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 63854 -5466
rect 63234 -5734 63854 -5702
rect 48954 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 49574 -6106
rect 48954 -6426 49574 -6342
rect 48954 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 49574 -6426
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 -2000
rect 77514 -2266 78134 -2000
rect 77514 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 78134 -2266
rect 77514 -2586 78134 -2502
rect 77514 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 78134 -2586
rect 77514 -3814 78134 -2822
rect 81234 -4186 81854 -2000
rect 81234 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 81854 -4186
rect 81234 -4506 81854 -4422
rect 81234 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 81854 -4506
rect 81234 -5734 81854 -4742
rect 66954 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 67574 -7066
rect 66954 -7386 67574 -7302
rect 66954 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 67574 -7386
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 -2000
rect 95514 -3226 96134 -2000
rect 95514 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 96134 -3226
rect 95514 -3546 96134 -3462
rect 95514 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 96134 -3546
rect 95514 -3814 96134 -3782
rect 99234 -5146 99854 -2000
rect 99234 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 99854 -5146
rect 99234 -5466 99854 -5382
rect 99234 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 99854 -5466
rect 99234 -5734 99854 -5702
rect 84954 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 85574 -6106
rect 84954 -6426 85574 -6342
rect 84954 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 85574 -6426
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 -2000
rect 113514 -2266 114134 -2000
rect 113514 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 114134 -2266
rect 113514 -2586 114134 -2502
rect 113514 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 114134 -2586
rect 113514 -3814 114134 -2822
rect 117234 -4186 117854 -2000
rect 117234 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 117854 -4186
rect 117234 -4506 117854 -4422
rect 117234 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 117854 -4506
rect 117234 -5734 117854 -4742
rect 102954 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 103574 -7066
rect 102954 -7386 103574 -7302
rect 102954 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 103574 -7386
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 -2000
rect 131514 -3226 132134 -2000
rect 131514 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 132134 -3226
rect 131514 -3546 132134 -3462
rect 131514 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 132134 -3546
rect 131514 -3814 132134 -3782
rect 135234 -5146 135854 -2000
rect 135234 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 135854 -5146
rect 135234 -5466 135854 -5382
rect 135234 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 135854 -5466
rect 135234 -5734 135854 -5702
rect 120954 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 121574 -6106
rect 120954 -6426 121574 -6342
rect 120954 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 121574 -6426
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 -2000
rect 149514 -2266 150134 -2000
rect 149514 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 150134 -2266
rect 149514 -2586 150134 -2502
rect 149514 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 150134 -2586
rect 149514 -3814 150134 -2822
rect 153234 -4186 153854 -2000
rect 153234 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 153854 -4186
rect 153234 -4506 153854 -4422
rect 153234 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 153854 -4506
rect 153234 -5734 153854 -4742
rect 138954 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 139574 -7066
rect 138954 -7386 139574 -7302
rect 138954 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 139574 -7386
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 -2000
rect 167514 -3226 168134 -2000
rect 167514 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 168134 -3226
rect 167514 -3546 168134 -3462
rect 167514 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 168134 -3546
rect 167514 -3814 168134 -3782
rect 171234 -5146 171854 -2000
rect 171234 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 171854 -5146
rect 171234 -5466 171854 -5382
rect 171234 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 171854 -5466
rect 171234 -5734 171854 -5702
rect 156954 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 157574 -6106
rect 156954 -6426 157574 -6342
rect 156954 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 157574 -6426
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 -2000
rect 185514 -2266 186134 -2000
rect 185514 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 186134 -2266
rect 185514 -2586 186134 -2502
rect 185514 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 186134 -2586
rect 185514 -3814 186134 -2822
rect 189234 -4186 189854 -2000
rect 189234 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 189854 -4186
rect 189234 -4506 189854 -4422
rect 189234 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 189854 -4506
rect 189234 -5734 189854 -4742
rect 174954 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 175574 -7066
rect 174954 -7386 175574 -7302
rect 174954 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 175574 -7386
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 -2000
rect 203514 -3226 204134 -2000
rect 203514 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 204134 -3226
rect 203514 -3546 204134 -3462
rect 203514 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 204134 -3546
rect 203514 -3814 204134 -3782
rect 207234 -5146 207854 -2000
rect 207234 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 207854 -5146
rect 207234 -5466 207854 -5382
rect 207234 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 207854 -5466
rect 207234 -5734 207854 -5702
rect 192954 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 193574 -6106
rect 192954 -6426 193574 -6342
rect 192954 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 193574 -6426
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 -2000
rect 221514 -2266 222134 -2000
rect 221514 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 222134 -2266
rect 221514 -2586 222134 -2502
rect 221514 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 222134 -2586
rect 221514 -3814 222134 -2822
rect 225234 -4186 225854 -2000
rect 225234 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 225854 -4186
rect 225234 -4506 225854 -4422
rect 225234 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 225854 -4506
rect 225234 -5734 225854 -4742
rect 210954 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 211574 -7066
rect 210954 -7386 211574 -7302
rect 210954 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 211574 -7386
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 -2000
rect 239514 -3226 240134 -2000
rect 239514 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 240134 -3226
rect 239514 -3546 240134 -3462
rect 239514 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 240134 -3546
rect 239514 -3814 240134 -3782
rect 243234 -5146 243854 -2000
rect 243234 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 243854 -5146
rect 243234 -5466 243854 -5382
rect 243234 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 243854 -5466
rect 243234 -5734 243854 -5702
rect 228954 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 229574 -6106
rect 228954 -6426 229574 -6342
rect 228954 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 229574 -6426
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 -2000
rect 257514 -2266 258134 -2000
rect 257514 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 258134 -2266
rect 257514 -2586 258134 -2502
rect 257514 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 258134 -2586
rect 257514 -3814 258134 -2822
rect 261234 -4186 261854 -2000
rect 261234 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 261854 -4186
rect 261234 -4506 261854 -4422
rect 261234 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 261854 -4506
rect 261234 -5734 261854 -4742
rect 246954 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 247574 -7066
rect 246954 -7386 247574 -7302
rect 246954 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 247574 -7386
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 -2000
rect 275514 -3226 276134 -2000
rect 275514 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 276134 -3226
rect 275514 -3546 276134 -3462
rect 275514 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 276134 -3546
rect 275514 -3814 276134 -3782
rect 279234 -5146 279854 -2000
rect 279234 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 279854 -5146
rect 279234 -5466 279854 -5382
rect 279234 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 279854 -5466
rect 279234 -5734 279854 -5702
rect 264954 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 265574 -6106
rect 264954 -6426 265574 -6342
rect 264954 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 265574 -6426
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 -2000
rect 293514 -2266 294134 -2000
rect 293514 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 294134 -2266
rect 293514 -2586 294134 -2502
rect 293514 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 294134 -2586
rect 293514 -3814 294134 -2822
rect 297234 -4186 297854 -2000
rect 297234 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 297854 -4186
rect 297234 -4506 297854 -4422
rect 297234 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 297854 -4506
rect 297234 -5734 297854 -4742
rect 282954 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 283574 -7066
rect 282954 -7386 283574 -7302
rect 282954 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 283574 -7386
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 -2000
rect 311514 -3226 312134 -2000
rect 311514 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 312134 -3226
rect 311514 -3546 312134 -3462
rect 311514 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 312134 -3546
rect 311514 -3814 312134 -3782
rect 315234 -5146 315854 -2000
rect 315234 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 315854 -5146
rect 315234 -5466 315854 -5382
rect 315234 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 315854 -5466
rect 315234 -5734 315854 -5702
rect 300954 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 301574 -6106
rect 300954 -6426 301574 -6342
rect 300954 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 301574 -6426
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 -2000
rect 329514 -2266 330134 -2000
rect 329514 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 330134 -2266
rect 329514 -2586 330134 -2502
rect 329514 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 330134 -2586
rect 329514 -3814 330134 -2822
rect 333234 -4186 333854 -2000
rect 333234 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 333854 -4186
rect 333234 -4506 333854 -4422
rect 333234 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 333854 -4506
rect 333234 -5734 333854 -4742
rect 318954 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 319574 -7066
rect 318954 -7386 319574 -7302
rect 318954 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 319574 -7386
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 -2000
rect 347514 -3226 348134 -2000
rect 347514 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 348134 -3226
rect 347514 -3546 348134 -3462
rect 347514 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 348134 -3546
rect 347514 -3814 348134 -3782
rect 351234 -5146 351854 -2000
rect 351234 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 351854 -5146
rect 351234 -5466 351854 -5382
rect 351234 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 351854 -5466
rect 351234 -5734 351854 -5702
rect 336954 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 337574 -6106
rect 336954 -6426 337574 -6342
rect 336954 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 337574 -6426
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 -2000
rect 365514 -2266 366134 -2000
rect 365514 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 366134 -2266
rect 365514 -2586 366134 -2502
rect 365514 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 366134 -2586
rect 365514 -3814 366134 -2822
rect 369234 -4186 369854 -2000
rect 369234 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 369854 -4186
rect 369234 -4506 369854 -4422
rect 369234 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 369854 -4506
rect 369234 -5734 369854 -4742
rect 354954 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 355574 -7066
rect 354954 -7386 355574 -7302
rect 354954 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 355574 -7386
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 -2000
rect 383514 -3226 384134 -2000
rect 383514 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 384134 -3226
rect 383514 -3546 384134 -3462
rect 383514 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 384134 -3546
rect 383514 -3814 384134 -3782
rect 387234 -5146 387854 -2000
rect 387234 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 387854 -5146
rect 387234 -5466 387854 -5382
rect 387234 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 387854 -5466
rect 387234 -5734 387854 -5702
rect 372954 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 373574 -6106
rect 372954 -6426 373574 -6342
rect 372954 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 373574 -6426
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 -2000
rect 401514 -2266 402134 -2000
rect 401514 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 402134 -2266
rect 401514 -2586 402134 -2502
rect 401514 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 402134 -2586
rect 401514 -3814 402134 -2822
rect 405234 -4186 405854 -2000
rect 405234 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 405854 -4186
rect 405234 -4506 405854 -4422
rect 405234 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 405854 -4506
rect 405234 -5734 405854 -4742
rect 390954 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 391574 -7066
rect 390954 -7386 391574 -7302
rect 390954 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 391574 -7386
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 -2000
rect 419514 -3226 420134 -2000
rect 419514 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 420134 -3226
rect 419514 -3546 420134 -3462
rect 419514 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 420134 -3546
rect 419514 -3814 420134 -3782
rect 423234 -5146 423854 -2000
rect 423234 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 423854 -5146
rect 423234 -5466 423854 -5382
rect 423234 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 423854 -5466
rect 423234 -5734 423854 -5702
rect 408954 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 409574 -6106
rect 408954 -6426 409574 -6342
rect 408954 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 409574 -6426
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 -2000
rect 437514 -2266 438134 -2000
rect 437514 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 438134 -2266
rect 437514 -2586 438134 -2502
rect 437514 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 438134 -2586
rect 437514 -3814 438134 -2822
rect 441234 -4186 441854 -2000
rect 441234 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 441854 -4186
rect 441234 -4506 441854 -4422
rect 441234 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 441854 -4506
rect 441234 -5734 441854 -4742
rect 426954 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 427574 -7066
rect 426954 -7386 427574 -7302
rect 426954 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 427574 -7386
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 -2000
rect 455514 -3226 456134 -2000
rect 455514 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 456134 -3226
rect 455514 -3546 456134 -3462
rect 455514 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 456134 -3546
rect 455514 -3814 456134 -3782
rect 459234 -5146 459854 -2000
rect 459234 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 459854 -5146
rect 459234 -5466 459854 -5382
rect 459234 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 459854 -5466
rect 459234 -5734 459854 -5702
rect 444954 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 445574 -6106
rect 444954 -6426 445574 -6342
rect 444954 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 445574 -6426
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 -2000
rect 473514 -2266 474134 -2000
rect 473514 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 474134 -2266
rect 473514 -2586 474134 -2502
rect 473514 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 474134 -2586
rect 473514 -3814 474134 -2822
rect 477234 -4186 477854 -2000
rect 477234 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 477854 -4186
rect 477234 -4506 477854 -4422
rect 477234 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 477854 -4506
rect 477234 -5734 477854 -4742
rect 462954 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 463574 -7066
rect 462954 -7386 463574 -7302
rect 462954 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 463574 -7386
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 -2000
rect 491514 -3226 492134 -2000
rect 491514 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 492134 -3226
rect 491514 -3546 492134 -3462
rect 491514 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 492134 -3546
rect 491514 -3814 492134 -3782
rect 495234 -5146 495854 -2000
rect 495234 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 495854 -5146
rect 495234 -5466 495854 -5382
rect 495234 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 495854 -5466
rect 495234 -5734 495854 -5702
rect 480954 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 481574 -6106
rect 480954 -6426 481574 -6342
rect 480954 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 481574 -6426
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 -2000
rect 509514 -2266 510134 -2000
rect 509514 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 510134 -2266
rect 509514 -2586 510134 -2502
rect 509514 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 510134 -2586
rect 509514 -3814 510134 -2822
rect 513234 -4186 513854 -2000
rect 513234 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 513854 -4186
rect 513234 -4506 513854 -4422
rect 513234 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 513854 -4506
rect 513234 -5734 513854 -4742
rect 498954 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 499574 -7066
rect 498954 -7386 499574 -7302
rect 498954 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 499574 -7386
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 -2000
rect 527514 -3226 528134 -2000
rect 527514 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 528134 -3226
rect 527514 -3546 528134 -3462
rect 527514 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 528134 -3546
rect 527514 -3814 528134 -3782
rect 531234 -5146 531854 -2000
rect 531234 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 531854 -5146
rect 531234 -5466 531854 -5382
rect 531234 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 531854 -5466
rect 531234 -5734 531854 -5702
rect 516954 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 517574 -6106
rect 516954 -6426 517574 -6342
rect 516954 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 517574 -6426
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 -2000
rect 545514 -2266 546134 -2000
rect 545514 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 546134 -2266
rect 545514 -2586 546134 -2502
rect 545514 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 546134 -2586
rect 545514 -3814 546134 -2822
rect 549234 -4186 549854 -2000
rect 549234 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 549854 -4186
rect 549234 -4506 549854 -4422
rect 549234 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 549854 -4506
rect 549234 -5734 549854 -4742
rect 534954 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 535574 -7066
rect 534954 -7386 535574 -7302
rect 534954 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 535574 -7386
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 -2000
rect 563514 -3226 564134 -2000
rect 563514 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 564134 -3226
rect 563514 -3546 564134 -3462
rect 563514 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 564134 -3546
rect 563514 -3814 564134 -3782
rect 567234 -5146 567854 28338
rect 567234 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 567854 -5146
rect 567234 -5466 567854 -5382
rect 567234 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 567854 -5466
rect 567234 -5734 567854 -5702
rect 570954 680614 571574 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 581514 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 582134 706758
rect 581514 706438 582134 706522
rect 581514 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 582134 706438
rect 570954 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 571574 680614
rect 570954 680294 571574 680378
rect 570954 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 571574 680294
rect 570954 644614 571574 680058
rect 570954 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 571574 644614
rect 570954 644294 571574 644378
rect 570954 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 571574 644294
rect 570954 608614 571574 644058
rect 570954 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 571574 608614
rect 570954 608294 571574 608378
rect 570954 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 571574 608294
rect 570954 572614 571574 608058
rect 570954 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 571574 572614
rect 570954 572294 571574 572378
rect 570954 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 571574 572294
rect 570954 536614 571574 572058
rect 570954 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 571574 536614
rect 570954 536294 571574 536378
rect 570954 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 571574 536294
rect 570954 500614 571574 536058
rect 570954 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 571574 500614
rect 570954 500294 571574 500378
rect 570954 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 571574 500294
rect 570954 464614 571574 500058
rect 570954 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 571574 464614
rect 570954 464294 571574 464378
rect 570954 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 571574 464294
rect 570954 428614 571574 464058
rect 570954 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 571574 428614
rect 570954 428294 571574 428378
rect 570954 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 571574 428294
rect 570954 392614 571574 428058
rect 570954 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 571574 392614
rect 570954 392294 571574 392378
rect 570954 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 571574 392294
rect 570954 356614 571574 392058
rect 570954 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 571574 356614
rect 570954 356294 571574 356378
rect 570954 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 571574 356294
rect 570954 320614 571574 356058
rect 570954 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 571574 320614
rect 570954 320294 571574 320378
rect 570954 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 571574 320294
rect 570954 284614 571574 320058
rect 570954 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 571574 284614
rect 570954 284294 571574 284378
rect 570954 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 571574 284294
rect 570954 248614 571574 284058
rect 570954 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 571574 248614
rect 570954 248294 571574 248378
rect 570954 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 571574 248294
rect 570954 212614 571574 248058
rect 570954 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 571574 212614
rect 570954 212294 571574 212378
rect 570954 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 571574 212294
rect 570954 176614 571574 212058
rect 570954 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 571574 176614
rect 570954 176294 571574 176378
rect 570954 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 571574 176294
rect 570954 140614 571574 176058
rect 570954 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 571574 140614
rect 570954 140294 571574 140378
rect 570954 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 571574 140294
rect 570954 104614 571574 140058
rect 570954 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 571574 104614
rect 570954 104294 571574 104378
rect 570954 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 571574 104294
rect 570954 68614 571574 104058
rect 570954 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 571574 68614
rect 570954 68294 571574 68378
rect 570954 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 571574 68294
rect 570954 32614 571574 68058
rect 570954 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 571574 32614
rect 570954 32294 571574 32378
rect 570954 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 571574 32294
rect 552954 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 553574 -6106
rect 552954 -6426 553574 -6342
rect 552954 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 553574 -6426
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 32058
rect 577794 704838 578414 705830
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 581514 691174 582134 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -2266 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 587850 691174
rect 587230 690854 587850 690938
rect 587230 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 587850 690854
rect 587230 655174 587850 690618
rect 587230 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 587850 655174
rect 587230 654854 587850 654938
rect 587230 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 587850 654854
rect 587230 619174 587850 654618
rect 587230 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 587850 619174
rect 587230 618854 587850 618938
rect 587230 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 587850 618854
rect 587230 583174 587850 618618
rect 587230 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 587850 583174
rect 587230 582854 587850 582938
rect 587230 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 587850 582854
rect 587230 547174 587850 582618
rect 587230 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 587850 547174
rect 587230 546854 587850 546938
rect 587230 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 587850 546854
rect 587230 511174 587850 546618
rect 587230 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 587850 511174
rect 587230 510854 587850 510938
rect 587230 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 587850 510854
rect 587230 475174 587850 510618
rect 587230 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 587850 475174
rect 587230 474854 587850 474938
rect 587230 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 587850 474854
rect 587230 439174 587850 474618
rect 587230 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 587850 439174
rect 587230 438854 587850 438938
rect 587230 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 587850 438854
rect 587230 403174 587850 438618
rect 587230 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 587850 403174
rect 587230 402854 587850 402938
rect 587230 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 587850 402854
rect 587230 367174 587850 402618
rect 587230 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 587850 367174
rect 587230 366854 587850 366938
rect 587230 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 587850 366854
rect 587230 331174 587850 366618
rect 587230 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 587850 331174
rect 587230 330854 587850 330938
rect 587230 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 587850 330854
rect 587230 295174 587850 330618
rect 587230 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 587850 295174
rect 587230 294854 587850 294938
rect 587230 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 587850 294854
rect 587230 259174 587850 294618
rect 587230 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 587850 259174
rect 587230 258854 587850 258938
rect 587230 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 587850 258854
rect 587230 223174 587850 258618
rect 587230 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 587850 223174
rect 587230 222854 587850 222938
rect 587230 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 587850 222854
rect 587230 187174 587850 222618
rect 587230 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 587850 187174
rect 587230 186854 587850 186938
rect 587230 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 587850 186854
rect 587230 151174 587850 186618
rect 587230 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 587850 151174
rect 587230 150854 587850 150938
rect 587230 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 587850 150854
rect 587230 115174 587850 150618
rect 587230 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 587850 115174
rect 587230 114854 587850 114938
rect 587230 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 587850 114854
rect 587230 79174 587850 114618
rect 587230 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 587850 79174
rect 587230 78854 587850 78938
rect 587230 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 587850 78854
rect 587230 43174 587850 78618
rect 587230 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 587850 43174
rect 587230 42854 587850 42938
rect 587230 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 587850 42854
rect 587230 7174 587850 42618
rect 587230 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 587850 7174
rect 587230 6854 587850 6938
rect 587230 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 587850 6854
rect 581514 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 582134 -2266
rect 581514 -2586 582134 -2502
rect 581514 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 582134 -2586
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect 588190 672854 588810 672938
rect 588190 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect 588190 637174 588810 672618
rect 588190 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect 588190 636854 588810 636938
rect 588190 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect 588190 601174 588810 636618
rect 588190 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect 588190 600854 588810 600938
rect 588190 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect 588190 565174 588810 600618
rect 588190 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect 588190 564854 588810 564938
rect 588190 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect 588190 529174 588810 564618
rect 588190 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect 588190 528854 588810 528938
rect 588190 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect 588190 493174 588810 528618
rect 588190 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect 588190 492854 588810 492938
rect 588190 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect 588190 457174 588810 492618
rect 588190 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect 588190 456854 588810 456938
rect 588190 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect 588190 421174 588810 456618
rect 588190 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 588190 420854 588810 420938
rect 588190 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 588190 385174 588810 420618
rect 588190 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 588190 384854 588810 384938
rect 588190 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 588190 349174 588810 384618
rect 588190 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 588190 348854 588810 348938
rect 588190 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 588190 313174 588810 348618
rect 588190 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 588190 312854 588810 312938
rect 588190 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 588190 277174 588810 312618
rect 588190 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 588190 276854 588810 276938
rect 588190 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 588190 241174 588810 276618
rect 588190 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 588190 240854 588810 240938
rect 588190 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 588190 205174 588810 240618
rect 588190 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 588190 204854 588810 204938
rect 588190 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 588190 169174 588810 204618
rect 588190 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 588190 168854 588810 168938
rect 588190 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 588190 133174 588810 168618
rect 588190 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 588190 132854 588810 132938
rect 588190 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 588190 97174 588810 132618
rect 588190 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 588190 96854 588810 96938
rect 588190 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 588190 61174 588810 96618
rect 588190 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 588190 60854 588810 60938
rect 588190 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 588190 25174 588810 60618
rect 588190 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect 588190 24854 588810 24938
rect 588190 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect 588190 -3226 588810 24618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 589770 694894
rect 589150 694574 589770 694658
rect 589150 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 589770 694574
rect 589150 658894 589770 694338
rect 589150 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 589770 658894
rect 589150 658574 589770 658658
rect 589150 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 589770 658574
rect 589150 622894 589770 658338
rect 589150 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 589770 622894
rect 589150 622574 589770 622658
rect 589150 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 589770 622574
rect 589150 586894 589770 622338
rect 589150 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 589770 586894
rect 589150 586574 589770 586658
rect 589150 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 589770 586574
rect 589150 550894 589770 586338
rect 589150 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 589770 550894
rect 589150 550574 589770 550658
rect 589150 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 589770 550574
rect 589150 514894 589770 550338
rect 589150 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 589770 514894
rect 589150 514574 589770 514658
rect 589150 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 589770 514574
rect 589150 478894 589770 514338
rect 589150 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 589770 478894
rect 589150 478574 589770 478658
rect 589150 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 589770 478574
rect 589150 442894 589770 478338
rect 589150 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 589770 442894
rect 589150 442574 589770 442658
rect 589150 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 589770 442574
rect 589150 406894 589770 442338
rect 589150 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 589770 406894
rect 589150 406574 589770 406658
rect 589150 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 589770 406574
rect 589150 370894 589770 406338
rect 589150 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 589770 370894
rect 589150 370574 589770 370658
rect 589150 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 589770 370574
rect 589150 334894 589770 370338
rect 589150 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 589770 334894
rect 589150 334574 589770 334658
rect 589150 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 589770 334574
rect 589150 298894 589770 334338
rect 589150 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 589770 298894
rect 589150 298574 589770 298658
rect 589150 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 589770 298574
rect 589150 262894 589770 298338
rect 589150 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 589770 262894
rect 589150 262574 589770 262658
rect 589150 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 589770 262574
rect 589150 226894 589770 262338
rect 589150 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 589770 226894
rect 589150 226574 589770 226658
rect 589150 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 589770 226574
rect 589150 190894 589770 226338
rect 589150 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 589770 190894
rect 589150 190574 589770 190658
rect 589150 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 589770 190574
rect 589150 154894 589770 190338
rect 589150 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 589770 154894
rect 589150 154574 589770 154658
rect 589150 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 589770 154574
rect 589150 118894 589770 154338
rect 589150 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 589770 118894
rect 589150 118574 589770 118658
rect 589150 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 589770 118574
rect 589150 82894 589770 118338
rect 589150 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 589770 82894
rect 589150 82574 589770 82658
rect 589150 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 589770 82574
rect 589150 46894 589770 82338
rect 589150 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 589770 46894
rect 589150 46574 589770 46658
rect 589150 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 589770 46574
rect 589150 10894 589770 46338
rect 589150 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 589770 10894
rect 589150 10574 589770 10658
rect 589150 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 589770 10574
rect 589150 -4186 589770 10338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect 590110 676574 590730 676658
rect 590110 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect 590110 640894 590730 676338
rect 590110 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect 590110 640574 590730 640658
rect 590110 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect 590110 604894 590730 640338
rect 590110 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect 590110 604574 590730 604658
rect 590110 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect 590110 568894 590730 604338
rect 590110 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect 590110 568574 590730 568658
rect 590110 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect 590110 532894 590730 568338
rect 590110 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect 590110 532574 590730 532658
rect 590110 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect 590110 496894 590730 532338
rect 590110 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect 590110 496574 590730 496658
rect 590110 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect 590110 460894 590730 496338
rect 590110 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect 590110 460574 590730 460658
rect 590110 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect 590110 424894 590730 460338
rect 590110 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 590110 424574 590730 424658
rect 590110 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 590110 388894 590730 424338
rect 590110 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 590110 388574 590730 388658
rect 590110 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 590110 352894 590730 388338
rect 590110 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 590110 352574 590730 352658
rect 590110 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 590110 316894 590730 352338
rect 590110 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 590110 316574 590730 316658
rect 590110 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 590110 280894 590730 316338
rect 590110 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 590110 280574 590730 280658
rect 590110 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 590110 244894 590730 280338
rect 590110 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 590110 244574 590730 244658
rect 590110 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 590110 208894 590730 244338
rect 590110 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 590110 208574 590730 208658
rect 590110 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 590110 172894 590730 208338
rect 590110 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 590110 172574 590730 172658
rect 590110 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 590110 136894 590730 172338
rect 590110 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 590110 136574 590730 136658
rect 590110 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 590110 100894 590730 136338
rect 590110 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 590110 100574 590730 100658
rect 590110 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 590110 64894 590730 100338
rect 590110 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 590110 64574 590730 64658
rect 590110 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 590110 28894 590730 64338
rect 590110 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect 590110 28574 590730 28658
rect 590110 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect 590110 -5146 590730 28338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 591690 698614
rect 591070 698294 591690 698378
rect 591070 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 591690 698294
rect 591070 662614 591690 698058
rect 591070 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 591690 662614
rect 591070 662294 591690 662378
rect 591070 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 591690 662294
rect 591070 626614 591690 662058
rect 591070 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 591690 626614
rect 591070 626294 591690 626378
rect 591070 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 591690 626294
rect 591070 590614 591690 626058
rect 591070 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 591690 590614
rect 591070 590294 591690 590378
rect 591070 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 591690 590294
rect 591070 554614 591690 590058
rect 591070 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 591690 554614
rect 591070 554294 591690 554378
rect 591070 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 591690 554294
rect 591070 518614 591690 554058
rect 591070 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 591690 518614
rect 591070 518294 591690 518378
rect 591070 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 591690 518294
rect 591070 482614 591690 518058
rect 591070 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 591690 482614
rect 591070 482294 591690 482378
rect 591070 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 591690 482294
rect 591070 446614 591690 482058
rect 591070 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 591690 446614
rect 591070 446294 591690 446378
rect 591070 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 591690 446294
rect 591070 410614 591690 446058
rect 591070 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 591690 410614
rect 591070 410294 591690 410378
rect 591070 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 591690 410294
rect 591070 374614 591690 410058
rect 591070 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 591690 374614
rect 591070 374294 591690 374378
rect 591070 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 591690 374294
rect 591070 338614 591690 374058
rect 591070 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 591690 338614
rect 591070 338294 591690 338378
rect 591070 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 591690 338294
rect 591070 302614 591690 338058
rect 591070 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 591690 302614
rect 591070 302294 591690 302378
rect 591070 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 591690 302294
rect 591070 266614 591690 302058
rect 591070 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 591690 266614
rect 591070 266294 591690 266378
rect 591070 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 591690 266294
rect 591070 230614 591690 266058
rect 591070 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 591690 230614
rect 591070 230294 591690 230378
rect 591070 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 591690 230294
rect 591070 194614 591690 230058
rect 591070 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 591690 194614
rect 591070 194294 591690 194378
rect 591070 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 591690 194294
rect 591070 158614 591690 194058
rect 591070 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 591690 158614
rect 591070 158294 591690 158378
rect 591070 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 591690 158294
rect 591070 122614 591690 158058
rect 591070 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 591690 122614
rect 591070 122294 591690 122378
rect 591070 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 591690 122294
rect 591070 86614 591690 122058
rect 591070 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 591690 86614
rect 591070 86294 591690 86378
rect 591070 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 591690 86294
rect 591070 50614 591690 86058
rect 591070 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 591690 50614
rect 591070 50294 591690 50378
rect 591070 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 591690 50294
rect 591070 14614 591690 50058
rect 591070 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 591690 14614
rect 591070 14294 591690 14378
rect 591070 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 591690 14294
rect 591070 -6106 591690 14058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect 592030 680294 592650 680378
rect 592030 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect 592030 644614 592650 680058
rect 592030 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect 592030 644294 592650 644378
rect 592030 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect 592030 608614 592650 644058
rect 592030 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect 592030 608294 592650 608378
rect 592030 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect 592030 572614 592650 608058
rect 592030 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect 592030 572294 592650 572378
rect 592030 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect 592030 536614 592650 572058
rect 592030 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect 592030 536294 592650 536378
rect 592030 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect 592030 500614 592650 536058
rect 592030 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect 592030 500294 592650 500378
rect 592030 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect 592030 464614 592650 500058
rect 592030 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect 592030 464294 592650 464378
rect 592030 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect 592030 428614 592650 464058
rect 592030 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 592030 428294 592650 428378
rect 592030 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 592030 392614 592650 428058
rect 592030 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 592030 392294 592650 392378
rect 592030 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 592030 356614 592650 392058
rect 592030 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 592030 356294 592650 356378
rect 592030 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 592030 320614 592650 356058
rect 592030 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 592030 320294 592650 320378
rect 592030 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 592030 284614 592650 320058
rect 592030 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 592030 284294 592650 284378
rect 592030 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 592030 248614 592650 284058
rect 592030 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 592030 248294 592650 248378
rect 592030 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 592030 212614 592650 248058
rect 592030 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 592030 212294 592650 212378
rect 592030 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 592030 176614 592650 212058
rect 592030 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 592030 176294 592650 176378
rect 592030 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 592030 140614 592650 176058
rect 592030 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 592030 140294 592650 140378
rect 592030 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 592030 104614 592650 140058
rect 592030 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 592030 104294 592650 104378
rect 592030 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 592030 68614 592650 104058
rect 592030 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 592030 68294 592650 68378
rect 592030 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 592030 32614 592650 68058
rect 592030 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect 592030 32294 592650 32378
rect 592030 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect 570954 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 571574 -7066
rect 570954 -7386 571574 -7302
rect 570954 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 571574 -7386
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 680378 -8458 680614
rect -8374 680378 -8138 680614
rect -8694 680058 -8458 680294
rect -8374 680058 -8138 680294
rect -8694 644378 -8458 644614
rect -8374 644378 -8138 644614
rect -8694 644058 -8458 644294
rect -8374 644058 -8138 644294
rect -8694 608378 -8458 608614
rect -8374 608378 -8138 608614
rect -8694 608058 -8458 608294
rect -8374 608058 -8138 608294
rect -8694 572378 -8458 572614
rect -8374 572378 -8138 572614
rect -8694 572058 -8458 572294
rect -8374 572058 -8138 572294
rect -8694 536378 -8458 536614
rect -8374 536378 -8138 536614
rect -8694 536058 -8458 536294
rect -8374 536058 -8138 536294
rect -8694 500378 -8458 500614
rect -8374 500378 -8138 500614
rect -8694 500058 -8458 500294
rect -8374 500058 -8138 500294
rect -8694 464378 -8458 464614
rect -8374 464378 -8138 464614
rect -8694 464058 -8458 464294
rect -8374 464058 -8138 464294
rect -8694 428378 -8458 428614
rect -8374 428378 -8138 428614
rect -8694 428058 -8458 428294
rect -8374 428058 -8138 428294
rect -8694 392378 -8458 392614
rect -8374 392378 -8138 392614
rect -8694 392058 -8458 392294
rect -8374 392058 -8138 392294
rect -8694 356378 -8458 356614
rect -8374 356378 -8138 356614
rect -8694 356058 -8458 356294
rect -8374 356058 -8138 356294
rect -8694 320378 -8458 320614
rect -8374 320378 -8138 320614
rect -8694 320058 -8458 320294
rect -8374 320058 -8138 320294
rect -8694 284378 -8458 284614
rect -8374 284378 -8138 284614
rect -8694 284058 -8458 284294
rect -8374 284058 -8138 284294
rect -8694 248378 -8458 248614
rect -8374 248378 -8138 248614
rect -8694 248058 -8458 248294
rect -8374 248058 -8138 248294
rect -8694 212378 -8458 212614
rect -8374 212378 -8138 212614
rect -8694 212058 -8458 212294
rect -8374 212058 -8138 212294
rect -8694 176378 -8458 176614
rect -8374 176378 -8138 176614
rect -8694 176058 -8458 176294
rect -8374 176058 -8138 176294
rect -8694 140378 -8458 140614
rect -8374 140378 -8138 140614
rect -8694 140058 -8458 140294
rect -8374 140058 -8138 140294
rect -8694 104378 -8458 104614
rect -8374 104378 -8138 104614
rect -8694 104058 -8458 104294
rect -8374 104058 -8138 104294
rect -8694 68378 -8458 68614
rect -8374 68378 -8138 68614
rect -8694 68058 -8458 68294
rect -8374 68058 -8138 68294
rect -8694 32378 -8458 32614
rect -8374 32378 -8138 32614
rect -8694 32058 -8458 32294
rect -8374 32058 -8138 32294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12986 710362 13222 710598
rect 13306 710362 13542 710598
rect 12986 710042 13222 710278
rect 13306 710042 13542 710278
rect -7734 698378 -7498 698614
rect -7414 698378 -7178 698614
rect -7734 698058 -7498 698294
rect -7414 698058 -7178 698294
rect -7734 662378 -7498 662614
rect -7414 662378 -7178 662614
rect -7734 662058 -7498 662294
rect -7414 662058 -7178 662294
rect -7734 626378 -7498 626614
rect -7414 626378 -7178 626614
rect -7734 626058 -7498 626294
rect -7414 626058 -7178 626294
rect -7734 590378 -7498 590614
rect -7414 590378 -7178 590614
rect -7734 590058 -7498 590294
rect -7414 590058 -7178 590294
rect -7734 554378 -7498 554614
rect -7414 554378 -7178 554614
rect -7734 554058 -7498 554294
rect -7414 554058 -7178 554294
rect -7734 518378 -7498 518614
rect -7414 518378 -7178 518614
rect -7734 518058 -7498 518294
rect -7414 518058 -7178 518294
rect -7734 482378 -7498 482614
rect -7414 482378 -7178 482614
rect -7734 482058 -7498 482294
rect -7414 482058 -7178 482294
rect -7734 446378 -7498 446614
rect -7414 446378 -7178 446614
rect -7734 446058 -7498 446294
rect -7414 446058 -7178 446294
rect -7734 410378 -7498 410614
rect -7414 410378 -7178 410614
rect -7734 410058 -7498 410294
rect -7414 410058 -7178 410294
rect -7734 374378 -7498 374614
rect -7414 374378 -7178 374614
rect -7734 374058 -7498 374294
rect -7414 374058 -7178 374294
rect -7734 338378 -7498 338614
rect -7414 338378 -7178 338614
rect -7734 338058 -7498 338294
rect -7414 338058 -7178 338294
rect -7734 302378 -7498 302614
rect -7414 302378 -7178 302614
rect -7734 302058 -7498 302294
rect -7414 302058 -7178 302294
rect -7734 266378 -7498 266614
rect -7414 266378 -7178 266614
rect -7734 266058 -7498 266294
rect -7414 266058 -7178 266294
rect -7734 230378 -7498 230614
rect -7414 230378 -7178 230614
rect -7734 230058 -7498 230294
rect -7414 230058 -7178 230294
rect -7734 194378 -7498 194614
rect -7414 194378 -7178 194614
rect -7734 194058 -7498 194294
rect -7414 194058 -7178 194294
rect -7734 158378 -7498 158614
rect -7414 158378 -7178 158614
rect -7734 158058 -7498 158294
rect -7414 158058 -7178 158294
rect -7734 122378 -7498 122614
rect -7414 122378 -7178 122614
rect -7734 122058 -7498 122294
rect -7414 122058 -7178 122294
rect -7734 86378 -7498 86614
rect -7414 86378 -7178 86614
rect -7734 86058 -7498 86294
rect -7414 86058 -7178 86294
rect -7734 50378 -7498 50614
rect -7414 50378 -7178 50614
rect -7734 50058 -7498 50294
rect -7414 50058 -7178 50294
rect -7734 14378 -7498 14614
rect -7414 14378 -7178 14614
rect -7734 14058 -7498 14294
rect -7414 14058 -7178 14294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 676658 -6538 676894
rect -6454 676658 -6218 676894
rect -6774 676338 -6538 676574
rect -6454 676338 -6218 676574
rect -6774 640658 -6538 640894
rect -6454 640658 -6218 640894
rect -6774 640338 -6538 640574
rect -6454 640338 -6218 640574
rect -6774 604658 -6538 604894
rect -6454 604658 -6218 604894
rect -6774 604338 -6538 604574
rect -6454 604338 -6218 604574
rect -6774 568658 -6538 568894
rect -6454 568658 -6218 568894
rect -6774 568338 -6538 568574
rect -6454 568338 -6218 568574
rect -6774 532658 -6538 532894
rect -6454 532658 -6218 532894
rect -6774 532338 -6538 532574
rect -6454 532338 -6218 532574
rect -6774 496658 -6538 496894
rect -6454 496658 -6218 496894
rect -6774 496338 -6538 496574
rect -6454 496338 -6218 496574
rect -6774 460658 -6538 460894
rect -6454 460658 -6218 460894
rect -6774 460338 -6538 460574
rect -6454 460338 -6218 460574
rect -6774 424658 -6538 424894
rect -6454 424658 -6218 424894
rect -6774 424338 -6538 424574
rect -6454 424338 -6218 424574
rect -6774 388658 -6538 388894
rect -6454 388658 -6218 388894
rect -6774 388338 -6538 388574
rect -6454 388338 -6218 388574
rect -6774 352658 -6538 352894
rect -6454 352658 -6218 352894
rect -6774 352338 -6538 352574
rect -6454 352338 -6218 352574
rect -6774 316658 -6538 316894
rect -6454 316658 -6218 316894
rect -6774 316338 -6538 316574
rect -6454 316338 -6218 316574
rect -6774 280658 -6538 280894
rect -6454 280658 -6218 280894
rect -6774 280338 -6538 280574
rect -6454 280338 -6218 280574
rect -6774 244658 -6538 244894
rect -6454 244658 -6218 244894
rect -6774 244338 -6538 244574
rect -6454 244338 -6218 244574
rect -6774 208658 -6538 208894
rect -6454 208658 -6218 208894
rect -6774 208338 -6538 208574
rect -6454 208338 -6218 208574
rect -6774 172658 -6538 172894
rect -6454 172658 -6218 172894
rect -6774 172338 -6538 172574
rect -6454 172338 -6218 172574
rect -6774 136658 -6538 136894
rect -6454 136658 -6218 136894
rect -6774 136338 -6538 136574
rect -6454 136338 -6218 136574
rect -6774 100658 -6538 100894
rect -6454 100658 -6218 100894
rect -6774 100338 -6538 100574
rect -6454 100338 -6218 100574
rect -6774 64658 -6538 64894
rect -6454 64658 -6218 64894
rect -6774 64338 -6538 64574
rect -6454 64338 -6218 64574
rect -6774 28658 -6538 28894
rect -6454 28658 -6218 28894
rect -6774 28338 -6538 28574
rect -6454 28338 -6218 28574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 9266 708442 9502 708678
rect 9586 708442 9822 708678
rect 9266 708122 9502 708358
rect 9586 708122 9822 708358
rect -5814 694658 -5578 694894
rect -5494 694658 -5258 694894
rect -5814 694338 -5578 694574
rect -5494 694338 -5258 694574
rect -5814 658658 -5578 658894
rect -5494 658658 -5258 658894
rect -5814 658338 -5578 658574
rect -5494 658338 -5258 658574
rect -5814 622658 -5578 622894
rect -5494 622658 -5258 622894
rect -5814 622338 -5578 622574
rect -5494 622338 -5258 622574
rect -5814 586658 -5578 586894
rect -5494 586658 -5258 586894
rect -5814 586338 -5578 586574
rect -5494 586338 -5258 586574
rect -5814 550658 -5578 550894
rect -5494 550658 -5258 550894
rect -5814 550338 -5578 550574
rect -5494 550338 -5258 550574
rect -5814 514658 -5578 514894
rect -5494 514658 -5258 514894
rect -5814 514338 -5578 514574
rect -5494 514338 -5258 514574
rect -5814 478658 -5578 478894
rect -5494 478658 -5258 478894
rect -5814 478338 -5578 478574
rect -5494 478338 -5258 478574
rect -5814 442658 -5578 442894
rect -5494 442658 -5258 442894
rect -5814 442338 -5578 442574
rect -5494 442338 -5258 442574
rect -5814 406658 -5578 406894
rect -5494 406658 -5258 406894
rect -5814 406338 -5578 406574
rect -5494 406338 -5258 406574
rect -5814 370658 -5578 370894
rect -5494 370658 -5258 370894
rect -5814 370338 -5578 370574
rect -5494 370338 -5258 370574
rect -5814 334658 -5578 334894
rect -5494 334658 -5258 334894
rect -5814 334338 -5578 334574
rect -5494 334338 -5258 334574
rect -5814 298658 -5578 298894
rect -5494 298658 -5258 298894
rect -5814 298338 -5578 298574
rect -5494 298338 -5258 298574
rect -5814 262658 -5578 262894
rect -5494 262658 -5258 262894
rect -5814 262338 -5578 262574
rect -5494 262338 -5258 262574
rect -5814 226658 -5578 226894
rect -5494 226658 -5258 226894
rect -5814 226338 -5578 226574
rect -5494 226338 -5258 226574
rect -5814 190658 -5578 190894
rect -5494 190658 -5258 190894
rect -5814 190338 -5578 190574
rect -5494 190338 -5258 190574
rect -5814 154658 -5578 154894
rect -5494 154658 -5258 154894
rect -5814 154338 -5578 154574
rect -5494 154338 -5258 154574
rect -5814 118658 -5578 118894
rect -5494 118658 -5258 118894
rect -5814 118338 -5578 118574
rect -5494 118338 -5258 118574
rect -5814 82658 -5578 82894
rect -5494 82658 -5258 82894
rect -5814 82338 -5578 82574
rect -5494 82338 -5258 82574
rect -5814 46658 -5578 46894
rect -5494 46658 -5258 46894
rect -5814 46338 -5578 46574
rect -5494 46338 -5258 46574
rect -5814 10658 -5578 10894
rect -5494 10658 -5258 10894
rect -5814 10338 -5578 10574
rect -5494 10338 -5258 10574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 672938 -4618 673174
rect -4534 672938 -4298 673174
rect -4854 672618 -4618 672854
rect -4534 672618 -4298 672854
rect -4854 636938 -4618 637174
rect -4534 636938 -4298 637174
rect -4854 636618 -4618 636854
rect -4534 636618 -4298 636854
rect -4854 600938 -4618 601174
rect -4534 600938 -4298 601174
rect -4854 600618 -4618 600854
rect -4534 600618 -4298 600854
rect -4854 564938 -4618 565174
rect -4534 564938 -4298 565174
rect -4854 564618 -4618 564854
rect -4534 564618 -4298 564854
rect -4854 528938 -4618 529174
rect -4534 528938 -4298 529174
rect -4854 528618 -4618 528854
rect -4534 528618 -4298 528854
rect -4854 492938 -4618 493174
rect -4534 492938 -4298 493174
rect -4854 492618 -4618 492854
rect -4534 492618 -4298 492854
rect -4854 456938 -4618 457174
rect -4534 456938 -4298 457174
rect -4854 456618 -4618 456854
rect -4534 456618 -4298 456854
rect -4854 420938 -4618 421174
rect -4534 420938 -4298 421174
rect -4854 420618 -4618 420854
rect -4534 420618 -4298 420854
rect -4854 384938 -4618 385174
rect -4534 384938 -4298 385174
rect -4854 384618 -4618 384854
rect -4534 384618 -4298 384854
rect -4854 348938 -4618 349174
rect -4534 348938 -4298 349174
rect -4854 348618 -4618 348854
rect -4534 348618 -4298 348854
rect -4854 312938 -4618 313174
rect -4534 312938 -4298 313174
rect -4854 312618 -4618 312854
rect -4534 312618 -4298 312854
rect -4854 276938 -4618 277174
rect -4534 276938 -4298 277174
rect -4854 276618 -4618 276854
rect -4534 276618 -4298 276854
rect -4854 240938 -4618 241174
rect -4534 240938 -4298 241174
rect -4854 240618 -4618 240854
rect -4534 240618 -4298 240854
rect -4854 204938 -4618 205174
rect -4534 204938 -4298 205174
rect -4854 204618 -4618 204854
rect -4534 204618 -4298 204854
rect -4854 168938 -4618 169174
rect -4534 168938 -4298 169174
rect -4854 168618 -4618 168854
rect -4534 168618 -4298 168854
rect -4854 132938 -4618 133174
rect -4534 132938 -4298 133174
rect -4854 132618 -4618 132854
rect -4534 132618 -4298 132854
rect -4854 96938 -4618 97174
rect -4534 96938 -4298 97174
rect -4854 96618 -4618 96854
rect -4534 96618 -4298 96854
rect -4854 60938 -4618 61174
rect -4534 60938 -4298 61174
rect -4854 60618 -4618 60854
rect -4534 60618 -4298 60854
rect -4854 24938 -4618 25174
rect -4534 24938 -4298 25174
rect -4854 24618 -4618 24854
rect -4534 24618 -4298 24854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 5546 706522 5782 706758
rect 5866 706522 6102 706758
rect 5546 706202 5782 706438
rect 5866 706202 6102 706438
rect -3894 690938 -3658 691174
rect -3574 690938 -3338 691174
rect -3894 690618 -3658 690854
rect -3574 690618 -3338 690854
rect -3894 654938 -3658 655174
rect -3574 654938 -3338 655174
rect -3894 654618 -3658 654854
rect -3574 654618 -3338 654854
rect -3894 618938 -3658 619174
rect -3574 618938 -3338 619174
rect -3894 618618 -3658 618854
rect -3574 618618 -3338 618854
rect -3894 582938 -3658 583174
rect -3574 582938 -3338 583174
rect -3894 582618 -3658 582854
rect -3574 582618 -3338 582854
rect -3894 546938 -3658 547174
rect -3574 546938 -3338 547174
rect -3894 546618 -3658 546854
rect -3574 546618 -3338 546854
rect -3894 510938 -3658 511174
rect -3574 510938 -3338 511174
rect -3894 510618 -3658 510854
rect -3574 510618 -3338 510854
rect -3894 474938 -3658 475174
rect -3574 474938 -3338 475174
rect -3894 474618 -3658 474854
rect -3574 474618 -3338 474854
rect -3894 438938 -3658 439174
rect -3574 438938 -3338 439174
rect -3894 438618 -3658 438854
rect -3574 438618 -3338 438854
rect -3894 402938 -3658 403174
rect -3574 402938 -3338 403174
rect -3894 402618 -3658 402854
rect -3574 402618 -3338 402854
rect -3894 366938 -3658 367174
rect -3574 366938 -3338 367174
rect -3894 366618 -3658 366854
rect -3574 366618 -3338 366854
rect -3894 330938 -3658 331174
rect -3574 330938 -3338 331174
rect -3894 330618 -3658 330854
rect -3574 330618 -3338 330854
rect -3894 294938 -3658 295174
rect -3574 294938 -3338 295174
rect -3894 294618 -3658 294854
rect -3574 294618 -3338 294854
rect -3894 258938 -3658 259174
rect -3574 258938 -3338 259174
rect -3894 258618 -3658 258854
rect -3574 258618 -3338 258854
rect -3894 222938 -3658 223174
rect -3574 222938 -3338 223174
rect -3894 222618 -3658 222854
rect -3574 222618 -3338 222854
rect -3894 186938 -3658 187174
rect -3574 186938 -3338 187174
rect -3894 186618 -3658 186854
rect -3574 186618 -3338 186854
rect -3894 150938 -3658 151174
rect -3574 150938 -3338 151174
rect -3894 150618 -3658 150854
rect -3574 150618 -3338 150854
rect -3894 114938 -3658 115174
rect -3574 114938 -3338 115174
rect -3894 114618 -3658 114854
rect -3574 114618 -3338 114854
rect -3894 78938 -3658 79174
rect -3574 78938 -3338 79174
rect -3894 78618 -3658 78854
rect -3574 78618 -3338 78854
rect -3894 42938 -3658 43174
rect -3574 42938 -3338 43174
rect -3894 42618 -3658 42854
rect -3574 42618 -3338 42854
rect -3894 6938 -3658 7174
rect -3574 6938 -3338 7174
rect -3894 6618 -3658 6854
rect -3574 6618 -3338 6854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 30986 711322 31222 711558
rect 31306 711322 31542 711558
rect 30986 711002 31222 711238
rect 31306 711002 31542 711238
rect 27266 709402 27502 709638
rect 27586 709402 27822 709638
rect 27266 709082 27502 709318
rect 27586 709082 27822 709318
rect 23546 707482 23782 707718
rect 23866 707482 24102 707718
rect 23546 707162 23782 707398
rect 23866 707162 24102 707398
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 48986 710362 49222 710598
rect 49306 710362 49542 710598
rect 48986 710042 49222 710278
rect 49306 710042 49542 710278
rect 45266 708442 45502 708678
rect 45586 708442 45822 708678
rect 45266 708122 45502 708358
rect 45586 708122 45822 708358
rect 41546 706522 41782 706758
rect 41866 706522 42102 706758
rect 41546 706202 41782 706438
rect 41866 706202 42102 706438
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 66986 711322 67222 711558
rect 67306 711322 67542 711558
rect 66986 711002 67222 711238
rect 67306 711002 67542 711238
rect 63266 709402 63502 709638
rect 63586 709402 63822 709638
rect 63266 709082 63502 709318
rect 63586 709082 63822 709318
rect 59546 707482 59782 707718
rect 59866 707482 60102 707718
rect 59546 707162 59782 707398
rect 59866 707162 60102 707398
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 84986 710362 85222 710598
rect 85306 710362 85542 710598
rect 84986 710042 85222 710278
rect 85306 710042 85542 710278
rect 81266 708442 81502 708678
rect 81586 708442 81822 708678
rect 81266 708122 81502 708358
rect 81586 708122 81822 708358
rect 77546 706522 77782 706758
rect 77866 706522 78102 706758
rect 77546 706202 77782 706438
rect 77866 706202 78102 706438
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 102986 711322 103222 711558
rect 103306 711322 103542 711558
rect 102986 711002 103222 711238
rect 103306 711002 103542 711238
rect 99266 709402 99502 709638
rect 99586 709402 99822 709638
rect 99266 709082 99502 709318
rect 99586 709082 99822 709318
rect 95546 707482 95782 707718
rect 95866 707482 96102 707718
rect 95546 707162 95782 707398
rect 95866 707162 96102 707398
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 120986 710362 121222 710598
rect 121306 710362 121542 710598
rect 120986 710042 121222 710278
rect 121306 710042 121542 710278
rect 117266 708442 117502 708678
rect 117586 708442 117822 708678
rect 117266 708122 117502 708358
rect 117586 708122 117822 708358
rect 113546 706522 113782 706758
rect 113866 706522 114102 706758
rect 113546 706202 113782 706438
rect 113866 706202 114102 706438
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 138986 711322 139222 711558
rect 139306 711322 139542 711558
rect 138986 711002 139222 711238
rect 139306 711002 139542 711238
rect 135266 709402 135502 709638
rect 135586 709402 135822 709638
rect 135266 709082 135502 709318
rect 135586 709082 135822 709318
rect 131546 707482 131782 707718
rect 131866 707482 132102 707718
rect 131546 707162 131782 707398
rect 131866 707162 132102 707398
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 156986 710362 157222 710598
rect 157306 710362 157542 710598
rect 156986 710042 157222 710278
rect 157306 710042 157542 710278
rect 153266 708442 153502 708678
rect 153586 708442 153822 708678
rect 153266 708122 153502 708358
rect 153586 708122 153822 708358
rect 149546 706522 149782 706758
rect 149866 706522 150102 706758
rect 149546 706202 149782 706438
rect 149866 706202 150102 706438
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 174986 711322 175222 711558
rect 175306 711322 175542 711558
rect 174986 711002 175222 711238
rect 175306 711002 175542 711238
rect 171266 709402 171502 709638
rect 171586 709402 171822 709638
rect 171266 709082 171502 709318
rect 171586 709082 171822 709318
rect 167546 707482 167782 707718
rect 167866 707482 168102 707718
rect 167546 707162 167782 707398
rect 167866 707162 168102 707398
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 192986 710362 193222 710598
rect 193306 710362 193542 710598
rect 192986 710042 193222 710278
rect 193306 710042 193542 710278
rect 189266 708442 189502 708678
rect 189586 708442 189822 708678
rect 189266 708122 189502 708358
rect 189586 708122 189822 708358
rect 185546 706522 185782 706758
rect 185866 706522 186102 706758
rect 185546 706202 185782 706438
rect 185866 706202 186102 706438
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 210986 711322 211222 711558
rect 211306 711322 211542 711558
rect 210986 711002 211222 711238
rect 211306 711002 211542 711238
rect 207266 709402 207502 709638
rect 207586 709402 207822 709638
rect 207266 709082 207502 709318
rect 207586 709082 207822 709318
rect 203546 707482 203782 707718
rect 203866 707482 204102 707718
rect 203546 707162 203782 707398
rect 203866 707162 204102 707398
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 228986 710362 229222 710598
rect 229306 710362 229542 710598
rect 228986 710042 229222 710278
rect 229306 710042 229542 710278
rect 225266 708442 225502 708678
rect 225586 708442 225822 708678
rect 225266 708122 225502 708358
rect 225586 708122 225822 708358
rect 221546 706522 221782 706758
rect 221866 706522 222102 706758
rect 221546 706202 221782 706438
rect 221866 706202 222102 706438
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 246986 711322 247222 711558
rect 247306 711322 247542 711558
rect 246986 711002 247222 711238
rect 247306 711002 247542 711238
rect 243266 709402 243502 709638
rect 243586 709402 243822 709638
rect 243266 709082 243502 709318
rect 243586 709082 243822 709318
rect 239546 707482 239782 707718
rect 239866 707482 240102 707718
rect 239546 707162 239782 707398
rect 239866 707162 240102 707398
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 264986 710362 265222 710598
rect 265306 710362 265542 710598
rect 264986 710042 265222 710278
rect 265306 710042 265542 710278
rect 261266 708442 261502 708678
rect 261586 708442 261822 708678
rect 261266 708122 261502 708358
rect 261586 708122 261822 708358
rect 257546 706522 257782 706758
rect 257866 706522 258102 706758
rect 257546 706202 257782 706438
rect 257866 706202 258102 706438
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 282986 711322 283222 711558
rect 283306 711322 283542 711558
rect 282986 711002 283222 711238
rect 283306 711002 283542 711238
rect 279266 709402 279502 709638
rect 279586 709402 279822 709638
rect 279266 709082 279502 709318
rect 279586 709082 279822 709318
rect 275546 707482 275782 707718
rect 275866 707482 276102 707718
rect 275546 707162 275782 707398
rect 275866 707162 276102 707398
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 300986 710362 301222 710598
rect 301306 710362 301542 710598
rect 300986 710042 301222 710278
rect 301306 710042 301542 710278
rect 297266 708442 297502 708678
rect 297586 708442 297822 708678
rect 297266 708122 297502 708358
rect 297586 708122 297822 708358
rect 293546 706522 293782 706758
rect 293866 706522 294102 706758
rect 293546 706202 293782 706438
rect 293866 706202 294102 706438
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 318986 711322 319222 711558
rect 319306 711322 319542 711558
rect 318986 711002 319222 711238
rect 319306 711002 319542 711238
rect 315266 709402 315502 709638
rect 315586 709402 315822 709638
rect 315266 709082 315502 709318
rect 315586 709082 315822 709318
rect 311546 707482 311782 707718
rect 311866 707482 312102 707718
rect 311546 707162 311782 707398
rect 311866 707162 312102 707398
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 336986 710362 337222 710598
rect 337306 710362 337542 710598
rect 336986 710042 337222 710278
rect 337306 710042 337542 710278
rect 333266 708442 333502 708678
rect 333586 708442 333822 708678
rect 333266 708122 333502 708358
rect 333586 708122 333822 708358
rect 329546 706522 329782 706758
rect 329866 706522 330102 706758
rect 329546 706202 329782 706438
rect 329866 706202 330102 706438
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 354986 711322 355222 711558
rect 355306 711322 355542 711558
rect 354986 711002 355222 711238
rect 355306 711002 355542 711238
rect 351266 709402 351502 709638
rect 351586 709402 351822 709638
rect 351266 709082 351502 709318
rect 351586 709082 351822 709318
rect 347546 707482 347782 707718
rect 347866 707482 348102 707718
rect 347546 707162 347782 707398
rect 347866 707162 348102 707398
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 372986 710362 373222 710598
rect 373306 710362 373542 710598
rect 372986 710042 373222 710278
rect 373306 710042 373542 710278
rect 369266 708442 369502 708678
rect 369586 708442 369822 708678
rect 369266 708122 369502 708358
rect 369586 708122 369822 708358
rect 365546 706522 365782 706758
rect 365866 706522 366102 706758
rect 365546 706202 365782 706438
rect 365866 706202 366102 706438
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 390986 711322 391222 711558
rect 391306 711322 391542 711558
rect 390986 711002 391222 711238
rect 391306 711002 391542 711238
rect 387266 709402 387502 709638
rect 387586 709402 387822 709638
rect 387266 709082 387502 709318
rect 387586 709082 387822 709318
rect 383546 707482 383782 707718
rect 383866 707482 384102 707718
rect 383546 707162 383782 707398
rect 383866 707162 384102 707398
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 408986 710362 409222 710598
rect 409306 710362 409542 710598
rect 408986 710042 409222 710278
rect 409306 710042 409542 710278
rect 405266 708442 405502 708678
rect 405586 708442 405822 708678
rect 405266 708122 405502 708358
rect 405586 708122 405822 708358
rect 401546 706522 401782 706758
rect 401866 706522 402102 706758
rect 401546 706202 401782 706438
rect 401866 706202 402102 706438
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 426986 711322 427222 711558
rect 427306 711322 427542 711558
rect 426986 711002 427222 711238
rect 427306 711002 427542 711238
rect 423266 709402 423502 709638
rect 423586 709402 423822 709638
rect 423266 709082 423502 709318
rect 423586 709082 423822 709318
rect 419546 707482 419782 707718
rect 419866 707482 420102 707718
rect 419546 707162 419782 707398
rect 419866 707162 420102 707398
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 444986 710362 445222 710598
rect 445306 710362 445542 710598
rect 444986 710042 445222 710278
rect 445306 710042 445542 710278
rect 441266 708442 441502 708678
rect 441586 708442 441822 708678
rect 441266 708122 441502 708358
rect 441586 708122 441822 708358
rect 437546 706522 437782 706758
rect 437866 706522 438102 706758
rect 437546 706202 437782 706438
rect 437866 706202 438102 706438
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 462986 711322 463222 711558
rect 463306 711322 463542 711558
rect 462986 711002 463222 711238
rect 463306 711002 463542 711238
rect 459266 709402 459502 709638
rect 459586 709402 459822 709638
rect 459266 709082 459502 709318
rect 459586 709082 459822 709318
rect 455546 707482 455782 707718
rect 455866 707482 456102 707718
rect 455546 707162 455782 707398
rect 455866 707162 456102 707398
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 480986 710362 481222 710598
rect 481306 710362 481542 710598
rect 480986 710042 481222 710278
rect 481306 710042 481542 710278
rect 477266 708442 477502 708678
rect 477586 708442 477822 708678
rect 477266 708122 477502 708358
rect 477586 708122 477822 708358
rect 473546 706522 473782 706758
rect 473866 706522 474102 706758
rect 473546 706202 473782 706438
rect 473866 706202 474102 706438
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 498986 711322 499222 711558
rect 499306 711322 499542 711558
rect 498986 711002 499222 711238
rect 499306 711002 499542 711238
rect 495266 709402 495502 709638
rect 495586 709402 495822 709638
rect 495266 709082 495502 709318
rect 495586 709082 495822 709318
rect 491546 707482 491782 707718
rect 491866 707482 492102 707718
rect 491546 707162 491782 707398
rect 491866 707162 492102 707398
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 516986 710362 517222 710598
rect 517306 710362 517542 710598
rect 516986 710042 517222 710278
rect 517306 710042 517542 710278
rect 513266 708442 513502 708678
rect 513586 708442 513822 708678
rect 513266 708122 513502 708358
rect 513586 708122 513822 708358
rect 509546 706522 509782 706758
rect 509866 706522 510102 706758
rect 509546 706202 509782 706438
rect 509866 706202 510102 706438
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 534986 711322 535222 711558
rect 535306 711322 535542 711558
rect 534986 711002 535222 711238
rect 535306 711002 535542 711238
rect 531266 709402 531502 709638
rect 531586 709402 531822 709638
rect 531266 709082 531502 709318
rect 531586 709082 531822 709318
rect 527546 707482 527782 707718
rect 527866 707482 528102 707718
rect 527546 707162 527782 707398
rect 527866 707162 528102 707398
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 552986 710362 553222 710598
rect 553306 710362 553542 710598
rect 552986 710042 553222 710278
rect 553306 710042 553542 710278
rect 549266 708442 549502 708678
rect 549586 708442 549822 708678
rect 549266 708122 549502 708358
rect 549586 708122 549822 708358
rect 545546 706522 545782 706758
rect 545866 706522 546102 706758
rect 545546 706202 545782 706438
rect 545866 706202 546102 706438
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 570986 711322 571222 711558
rect 571306 711322 571542 711558
rect 570986 711002 571222 711238
rect 571306 711002 571542 711238
rect 567266 709402 567502 709638
rect 567586 709402 567822 709638
rect 567266 709082 567502 709318
rect 567586 709082 567822 709318
rect 563546 707482 563782 707718
rect 563866 707482 564102 707718
rect 563546 707162 563782 707398
rect 563866 707162 564102 707398
rect 559826 705562 560062 705798
rect 560146 705562 560382 705798
rect 559826 705242 560062 705478
rect 560146 705242 560382 705478
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect 8250 687218 8486 687454
rect 8250 686898 8486 687134
rect 38970 687218 39206 687454
rect 38970 686898 39206 687134
rect 69690 687218 69926 687454
rect 69690 686898 69926 687134
rect 100410 687218 100646 687454
rect 100410 686898 100646 687134
rect 131130 687218 131366 687454
rect 131130 686898 131366 687134
rect 161850 687218 162086 687454
rect 161850 686898 162086 687134
rect 192570 687218 192806 687454
rect 192570 686898 192806 687134
rect 223290 687218 223526 687454
rect 223290 686898 223526 687134
rect 254010 687218 254246 687454
rect 254010 686898 254246 687134
rect 284730 687218 284966 687454
rect 284730 686898 284966 687134
rect 315450 687218 315686 687454
rect 315450 686898 315686 687134
rect 346170 687218 346406 687454
rect 346170 686898 346406 687134
rect 376890 687218 377126 687454
rect 376890 686898 377126 687134
rect 407610 687218 407846 687454
rect 407610 686898 407846 687134
rect 438330 687218 438566 687454
rect 438330 686898 438566 687134
rect 469050 687218 469286 687454
rect 469050 686898 469286 687134
rect 499770 687218 500006 687454
rect 499770 686898 500006 687134
rect 530490 687218 530726 687454
rect 530490 686898 530726 687134
rect 561210 687218 561446 687454
rect 561210 686898 561446 687134
rect 567266 676658 567502 676894
rect 567586 676658 567822 676894
rect 567266 676338 567502 676574
rect 567586 676338 567822 676574
rect 23610 669218 23846 669454
rect 23610 668898 23846 669134
rect 54330 669218 54566 669454
rect 54330 668898 54566 669134
rect 85050 669218 85286 669454
rect 85050 668898 85286 669134
rect 115770 669218 116006 669454
rect 115770 668898 116006 669134
rect 146490 669218 146726 669454
rect 146490 668898 146726 669134
rect 177210 669218 177446 669454
rect 177210 668898 177446 669134
rect 207930 669218 208166 669454
rect 207930 668898 208166 669134
rect 238650 669218 238886 669454
rect 238650 668898 238886 669134
rect 269370 669218 269606 669454
rect 269370 668898 269606 669134
rect 300090 669218 300326 669454
rect 300090 668898 300326 669134
rect 330810 669218 331046 669454
rect 330810 668898 331046 669134
rect 361530 669218 361766 669454
rect 361530 668898 361766 669134
rect 392250 669218 392486 669454
rect 392250 668898 392486 669134
rect 422970 669218 423206 669454
rect 422970 668898 423206 669134
rect 453690 669218 453926 669454
rect 453690 668898 453926 669134
rect 484410 669218 484646 669454
rect 484410 668898 484646 669134
rect 515130 669218 515366 669454
rect 515130 668898 515366 669134
rect 545850 669218 546086 669454
rect 545850 668898 546086 669134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect 8250 651218 8486 651454
rect 8250 650898 8486 651134
rect 38970 651218 39206 651454
rect 38970 650898 39206 651134
rect 69690 651218 69926 651454
rect 69690 650898 69926 651134
rect 100410 651218 100646 651454
rect 100410 650898 100646 651134
rect 131130 651218 131366 651454
rect 131130 650898 131366 651134
rect 161850 651218 162086 651454
rect 161850 650898 162086 651134
rect 192570 651218 192806 651454
rect 192570 650898 192806 651134
rect 223290 651218 223526 651454
rect 223290 650898 223526 651134
rect 254010 651218 254246 651454
rect 254010 650898 254246 651134
rect 284730 651218 284966 651454
rect 284730 650898 284966 651134
rect 315450 651218 315686 651454
rect 315450 650898 315686 651134
rect 346170 651218 346406 651454
rect 346170 650898 346406 651134
rect 376890 651218 377126 651454
rect 376890 650898 377126 651134
rect 407610 651218 407846 651454
rect 407610 650898 407846 651134
rect 438330 651218 438566 651454
rect 438330 650898 438566 651134
rect 469050 651218 469286 651454
rect 469050 650898 469286 651134
rect 499770 651218 500006 651454
rect 499770 650898 500006 651134
rect 530490 651218 530726 651454
rect 530490 650898 530726 651134
rect 561210 651218 561446 651454
rect 561210 650898 561446 651134
rect 567266 640658 567502 640894
rect 567586 640658 567822 640894
rect 567266 640338 567502 640574
rect 567586 640338 567822 640574
rect 23610 633218 23846 633454
rect 23610 632898 23846 633134
rect 54330 633218 54566 633454
rect 54330 632898 54566 633134
rect 85050 633218 85286 633454
rect 85050 632898 85286 633134
rect 115770 633218 116006 633454
rect 115770 632898 116006 633134
rect 146490 633218 146726 633454
rect 146490 632898 146726 633134
rect 177210 633218 177446 633454
rect 177210 632898 177446 633134
rect 207930 633218 208166 633454
rect 207930 632898 208166 633134
rect 238650 633218 238886 633454
rect 238650 632898 238886 633134
rect 269370 633218 269606 633454
rect 269370 632898 269606 633134
rect 300090 633218 300326 633454
rect 300090 632898 300326 633134
rect 330810 633218 331046 633454
rect 330810 632898 331046 633134
rect 361530 633218 361766 633454
rect 361530 632898 361766 633134
rect 392250 633218 392486 633454
rect 392250 632898 392486 633134
rect 422970 633218 423206 633454
rect 422970 632898 423206 633134
rect 453690 633218 453926 633454
rect 453690 632898 453926 633134
rect 484410 633218 484646 633454
rect 484410 632898 484646 633134
rect 515130 633218 515366 633454
rect 515130 632898 515366 633134
rect 545850 633218 546086 633454
rect 545850 632898 546086 633134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect 8250 615218 8486 615454
rect 8250 614898 8486 615134
rect 38970 615218 39206 615454
rect 38970 614898 39206 615134
rect 69690 615218 69926 615454
rect 69690 614898 69926 615134
rect 100410 615218 100646 615454
rect 100410 614898 100646 615134
rect 131130 615218 131366 615454
rect 131130 614898 131366 615134
rect 161850 615218 162086 615454
rect 161850 614898 162086 615134
rect 192570 615218 192806 615454
rect 192570 614898 192806 615134
rect 223290 615218 223526 615454
rect 223290 614898 223526 615134
rect 254010 615218 254246 615454
rect 254010 614898 254246 615134
rect 284730 615218 284966 615454
rect 284730 614898 284966 615134
rect 315450 615218 315686 615454
rect 315450 614898 315686 615134
rect 346170 615218 346406 615454
rect 346170 614898 346406 615134
rect 376890 615218 377126 615454
rect 376890 614898 377126 615134
rect 407610 615218 407846 615454
rect 407610 614898 407846 615134
rect 438330 615218 438566 615454
rect 438330 614898 438566 615134
rect 469050 615218 469286 615454
rect 469050 614898 469286 615134
rect 499770 615218 500006 615454
rect 499770 614898 500006 615134
rect 530490 615218 530726 615454
rect 530490 614898 530726 615134
rect 561210 615218 561446 615454
rect 561210 614898 561446 615134
rect 567266 604658 567502 604894
rect 567586 604658 567822 604894
rect 567266 604338 567502 604574
rect 567586 604338 567822 604574
rect 23610 597218 23846 597454
rect 23610 596898 23846 597134
rect 54330 597218 54566 597454
rect 54330 596898 54566 597134
rect 85050 597218 85286 597454
rect 85050 596898 85286 597134
rect 115770 597218 116006 597454
rect 115770 596898 116006 597134
rect 146490 597218 146726 597454
rect 146490 596898 146726 597134
rect 177210 597218 177446 597454
rect 177210 596898 177446 597134
rect 207930 597218 208166 597454
rect 207930 596898 208166 597134
rect 238650 597218 238886 597454
rect 238650 596898 238886 597134
rect 269370 597218 269606 597454
rect 269370 596898 269606 597134
rect 300090 597218 300326 597454
rect 300090 596898 300326 597134
rect 330810 597218 331046 597454
rect 330810 596898 331046 597134
rect 361530 597218 361766 597454
rect 361530 596898 361766 597134
rect 392250 597218 392486 597454
rect 392250 596898 392486 597134
rect 422970 597218 423206 597454
rect 422970 596898 423206 597134
rect 453690 597218 453926 597454
rect 453690 596898 453926 597134
rect 484410 597218 484646 597454
rect 484410 596898 484646 597134
rect 515130 597218 515366 597454
rect 515130 596898 515366 597134
rect 545850 597218 546086 597454
rect 545850 596898 546086 597134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect 8250 579218 8486 579454
rect 8250 578898 8486 579134
rect 38970 579218 39206 579454
rect 38970 578898 39206 579134
rect 69690 579218 69926 579454
rect 69690 578898 69926 579134
rect 100410 579218 100646 579454
rect 100410 578898 100646 579134
rect 131130 579218 131366 579454
rect 131130 578898 131366 579134
rect 161850 579218 162086 579454
rect 161850 578898 162086 579134
rect 192570 579218 192806 579454
rect 192570 578898 192806 579134
rect 223290 579218 223526 579454
rect 223290 578898 223526 579134
rect 254010 579218 254246 579454
rect 254010 578898 254246 579134
rect 284730 579218 284966 579454
rect 284730 578898 284966 579134
rect 315450 579218 315686 579454
rect 315450 578898 315686 579134
rect 346170 579218 346406 579454
rect 346170 578898 346406 579134
rect 376890 579218 377126 579454
rect 376890 578898 377126 579134
rect 407610 579218 407846 579454
rect 407610 578898 407846 579134
rect 438330 579218 438566 579454
rect 438330 578898 438566 579134
rect 469050 579218 469286 579454
rect 469050 578898 469286 579134
rect 499770 579218 500006 579454
rect 499770 578898 500006 579134
rect 530490 579218 530726 579454
rect 530490 578898 530726 579134
rect 561210 579218 561446 579454
rect 561210 578898 561446 579134
rect 567266 568658 567502 568894
rect 567586 568658 567822 568894
rect 567266 568338 567502 568574
rect 567586 568338 567822 568574
rect 23610 561218 23846 561454
rect 23610 560898 23846 561134
rect 54330 561218 54566 561454
rect 54330 560898 54566 561134
rect 85050 561218 85286 561454
rect 85050 560898 85286 561134
rect 115770 561218 116006 561454
rect 115770 560898 116006 561134
rect 146490 561218 146726 561454
rect 146490 560898 146726 561134
rect 177210 561218 177446 561454
rect 177210 560898 177446 561134
rect 207930 561218 208166 561454
rect 207930 560898 208166 561134
rect 238650 561218 238886 561454
rect 238650 560898 238886 561134
rect 269370 561218 269606 561454
rect 269370 560898 269606 561134
rect 300090 561218 300326 561454
rect 300090 560898 300326 561134
rect 330810 561218 331046 561454
rect 330810 560898 331046 561134
rect 361530 561218 361766 561454
rect 361530 560898 361766 561134
rect 392250 561218 392486 561454
rect 392250 560898 392486 561134
rect 422970 561218 423206 561454
rect 422970 560898 423206 561134
rect 453690 561218 453926 561454
rect 453690 560898 453926 561134
rect 484410 561218 484646 561454
rect 484410 560898 484646 561134
rect 515130 561218 515366 561454
rect 515130 560898 515366 561134
rect 545850 561218 546086 561454
rect 545850 560898 546086 561134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect 8250 543218 8486 543454
rect 8250 542898 8486 543134
rect 38970 543218 39206 543454
rect 38970 542898 39206 543134
rect 69690 543218 69926 543454
rect 69690 542898 69926 543134
rect 100410 543218 100646 543454
rect 100410 542898 100646 543134
rect 131130 543218 131366 543454
rect 131130 542898 131366 543134
rect 161850 543218 162086 543454
rect 161850 542898 162086 543134
rect 192570 543218 192806 543454
rect 192570 542898 192806 543134
rect 223290 543218 223526 543454
rect 223290 542898 223526 543134
rect 254010 543218 254246 543454
rect 254010 542898 254246 543134
rect 284730 543218 284966 543454
rect 284730 542898 284966 543134
rect 315450 543218 315686 543454
rect 315450 542898 315686 543134
rect 346170 543218 346406 543454
rect 346170 542898 346406 543134
rect 376890 543218 377126 543454
rect 376890 542898 377126 543134
rect 407610 543218 407846 543454
rect 407610 542898 407846 543134
rect 438330 543218 438566 543454
rect 438330 542898 438566 543134
rect 469050 543218 469286 543454
rect 469050 542898 469286 543134
rect 499770 543218 500006 543454
rect 499770 542898 500006 543134
rect 530490 543218 530726 543454
rect 530490 542898 530726 543134
rect 561210 543218 561446 543454
rect 561210 542898 561446 543134
rect 567266 532658 567502 532894
rect 567586 532658 567822 532894
rect 567266 532338 567502 532574
rect 567586 532338 567822 532574
rect 23610 525218 23846 525454
rect 23610 524898 23846 525134
rect 54330 525218 54566 525454
rect 54330 524898 54566 525134
rect 85050 525218 85286 525454
rect 85050 524898 85286 525134
rect 115770 525218 116006 525454
rect 115770 524898 116006 525134
rect 146490 525218 146726 525454
rect 146490 524898 146726 525134
rect 177210 525218 177446 525454
rect 177210 524898 177446 525134
rect 207930 525218 208166 525454
rect 207930 524898 208166 525134
rect 238650 525218 238886 525454
rect 238650 524898 238886 525134
rect 269370 525218 269606 525454
rect 269370 524898 269606 525134
rect 300090 525218 300326 525454
rect 300090 524898 300326 525134
rect 330810 525218 331046 525454
rect 330810 524898 331046 525134
rect 361530 525218 361766 525454
rect 361530 524898 361766 525134
rect 392250 525218 392486 525454
rect 392250 524898 392486 525134
rect 422970 525218 423206 525454
rect 422970 524898 423206 525134
rect 453690 525218 453926 525454
rect 453690 524898 453926 525134
rect 484410 525218 484646 525454
rect 484410 524898 484646 525134
rect 515130 525218 515366 525454
rect 515130 524898 515366 525134
rect 545850 525218 546086 525454
rect 545850 524898 546086 525134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect 8250 507218 8486 507454
rect 8250 506898 8486 507134
rect 38970 507218 39206 507454
rect 38970 506898 39206 507134
rect 69690 507218 69926 507454
rect 69690 506898 69926 507134
rect 100410 507218 100646 507454
rect 100410 506898 100646 507134
rect 131130 507218 131366 507454
rect 131130 506898 131366 507134
rect 161850 507218 162086 507454
rect 161850 506898 162086 507134
rect 192570 507218 192806 507454
rect 192570 506898 192806 507134
rect 223290 507218 223526 507454
rect 223290 506898 223526 507134
rect 254010 507218 254246 507454
rect 254010 506898 254246 507134
rect 284730 507218 284966 507454
rect 284730 506898 284966 507134
rect 315450 507218 315686 507454
rect 315450 506898 315686 507134
rect 346170 507218 346406 507454
rect 346170 506898 346406 507134
rect 376890 507218 377126 507454
rect 376890 506898 377126 507134
rect 407610 507218 407846 507454
rect 407610 506898 407846 507134
rect 438330 507218 438566 507454
rect 438330 506898 438566 507134
rect 469050 507218 469286 507454
rect 469050 506898 469286 507134
rect 499770 507218 500006 507454
rect 499770 506898 500006 507134
rect 530490 507218 530726 507454
rect 530490 506898 530726 507134
rect 561210 507218 561446 507454
rect 561210 506898 561446 507134
rect 567266 496658 567502 496894
rect 567586 496658 567822 496894
rect 567266 496338 567502 496574
rect 567586 496338 567822 496574
rect 23610 489218 23846 489454
rect 23610 488898 23846 489134
rect 54330 489218 54566 489454
rect 54330 488898 54566 489134
rect 85050 489218 85286 489454
rect 85050 488898 85286 489134
rect 115770 489218 116006 489454
rect 115770 488898 116006 489134
rect 146490 489218 146726 489454
rect 146490 488898 146726 489134
rect 177210 489218 177446 489454
rect 177210 488898 177446 489134
rect 207930 489218 208166 489454
rect 207930 488898 208166 489134
rect 238650 489218 238886 489454
rect 238650 488898 238886 489134
rect 269370 489218 269606 489454
rect 269370 488898 269606 489134
rect 300090 489218 300326 489454
rect 300090 488898 300326 489134
rect 330810 489218 331046 489454
rect 330810 488898 331046 489134
rect 361530 489218 361766 489454
rect 361530 488898 361766 489134
rect 392250 489218 392486 489454
rect 392250 488898 392486 489134
rect 422970 489218 423206 489454
rect 422970 488898 423206 489134
rect 453690 489218 453926 489454
rect 453690 488898 453926 489134
rect 484410 489218 484646 489454
rect 484410 488898 484646 489134
rect 515130 489218 515366 489454
rect 515130 488898 515366 489134
rect 545850 489218 546086 489454
rect 545850 488898 546086 489134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect 8250 471218 8486 471454
rect 8250 470898 8486 471134
rect 38970 471218 39206 471454
rect 38970 470898 39206 471134
rect 69690 471218 69926 471454
rect 69690 470898 69926 471134
rect 100410 471218 100646 471454
rect 100410 470898 100646 471134
rect 131130 471218 131366 471454
rect 131130 470898 131366 471134
rect 161850 471218 162086 471454
rect 161850 470898 162086 471134
rect 192570 471218 192806 471454
rect 192570 470898 192806 471134
rect 223290 471218 223526 471454
rect 223290 470898 223526 471134
rect 254010 471218 254246 471454
rect 254010 470898 254246 471134
rect 284730 471218 284966 471454
rect 284730 470898 284966 471134
rect 315450 471218 315686 471454
rect 315450 470898 315686 471134
rect 346170 471218 346406 471454
rect 346170 470898 346406 471134
rect 376890 471218 377126 471454
rect 376890 470898 377126 471134
rect 407610 471218 407846 471454
rect 407610 470898 407846 471134
rect 438330 471218 438566 471454
rect 438330 470898 438566 471134
rect 469050 471218 469286 471454
rect 469050 470898 469286 471134
rect 499770 471218 500006 471454
rect 499770 470898 500006 471134
rect 530490 471218 530726 471454
rect 530490 470898 530726 471134
rect 561210 471218 561446 471454
rect 561210 470898 561446 471134
rect 567266 460658 567502 460894
rect 567586 460658 567822 460894
rect 567266 460338 567502 460574
rect 567586 460338 567822 460574
rect 23610 453218 23846 453454
rect 23610 452898 23846 453134
rect 54330 453218 54566 453454
rect 54330 452898 54566 453134
rect 85050 453218 85286 453454
rect 85050 452898 85286 453134
rect 115770 453218 116006 453454
rect 115770 452898 116006 453134
rect 146490 453218 146726 453454
rect 146490 452898 146726 453134
rect 177210 453218 177446 453454
rect 177210 452898 177446 453134
rect 207930 453218 208166 453454
rect 207930 452898 208166 453134
rect 238650 453218 238886 453454
rect 238650 452898 238886 453134
rect 269370 453218 269606 453454
rect 269370 452898 269606 453134
rect 300090 453218 300326 453454
rect 300090 452898 300326 453134
rect 330810 453218 331046 453454
rect 330810 452898 331046 453134
rect 361530 453218 361766 453454
rect 361530 452898 361766 453134
rect 392250 453218 392486 453454
rect 392250 452898 392486 453134
rect 422970 453218 423206 453454
rect 422970 452898 423206 453134
rect 453690 453218 453926 453454
rect 453690 452898 453926 453134
rect 484410 453218 484646 453454
rect 484410 452898 484646 453134
rect 515130 453218 515366 453454
rect 515130 452898 515366 453134
rect 545850 453218 546086 453454
rect 545850 452898 546086 453134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect 8250 435218 8486 435454
rect 8250 434898 8486 435134
rect 38970 435218 39206 435454
rect 38970 434898 39206 435134
rect 69690 435218 69926 435454
rect 69690 434898 69926 435134
rect 100410 435218 100646 435454
rect 100410 434898 100646 435134
rect 131130 435218 131366 435454
rect 131130 434898 131366 435134
rect 161850 435218 162086 435454
rect 161850 434898 162086 435134
rect 192570 435218 192806 435454
rect 192570 434898 192806 435134
rect 223290 435218 223526 435454
rect 223290 434898 223526 435134
rect 254010 435218 254246 435454
rect 254010 434898 254246 435134
rect 284730 435218 284966 435454
rect 284730 434898 284966 435134
rect 315450 435218 315686 435454
rect 315450 434898 315686 435134
rect 346170 435218 346406 435454
rect 346170 434898 346406 435134
rect 376890 435218 377126 435454
rect 376890 434898 377126 435134
rect 407610 435218 407846 435454
rect 407610 434898 407846 435134
rect 438330 435218 438566 435454
rect 438330 434898 438566 435134
rect 469050 435218 469286 435454
rect 469050 434898 469286 435134
rect 499770 435218 500006 435454
rect 499770 434898 500006 435134
rect 530490 435218 530726 435454
rect 530490 434898 530726 435134
rect 561210 435218 561446 435454
rect 561210 434898 561446 435134
rect 567266 424658 567502 424894
rect 567586 424658 567822 424894
rect 567266 424338 567502 424574
rect 567586 424338 567822 424574
rect 23610 417218 23846 417454
rect 23610 416898 23846 417134
rect 54330 417218 54566 417454
rect 54330 416898 54566 417134
rect 85050 417218 85286 417454
rect 85050 416898 85286 417134
rect 115770 417218 116006 417454
rect 115770 416898 116006 417134
rect 146490 417218 146726 417454
rect 146490 416898 146726 417134
rect 177210 417218 177446 417454
rect 177210 416898 177446 417134
rect 207930 417218 208166 417454
rect 207930 416898 208166 417134
rect 238650 417218 238886 417454
rect 238650 416898 238886 417134
rect 269370 417218 269606 417454
rect 269370 416898 269606 417134
rect 300090 417218 300326 417454
rect 300090 416898 300326 417134
rect 330810 417218 331046 417454
rect 330810 416898 331046 417134
rect 361530 417218 361766 417454
rect 361530 416898 361766 417134
rect 392250 417218 392486 417454
rect 392250 416898 392486 417134
rect 422970 417218 423206 417454
rect 422970 416898 423206 417134
rect 453690 417218 453926 417454
rect 453690 416898 453926 417134
rect 484410 417218 484646 417454
rect 484410 416898 484646 417134
rect 515130 417218 515366 417454
rect 515130 416898 515366 417134
rect 545850 417218 546086 417454
rect 545850 416898 546086 417134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect 8250 399218 8486 399454
rect 8250 398898 8486 399134
rect 38970 399218 39206 399454
rect 38970 398898 39206 399134
rect 69690 399218 69926 399454
rect 69690 398898 69926 399134
rect 100410 399218 100646 399454
rect 100410 398898 100646 399134
rect 131130 399218 131366 399454
rect 131130 398898 131366 399134
rect 161850 399218 162086 399454
rect 161850 398898 162086 399134
rect 192570 399218 192806 399454
rect 192570 398898 192806 399134
rect 223290 399218 223526 399454
rect 223290 398898 223526 399134
rect 254010 399218 254246 399454
rect 254010 398898 254246 399134
rect 284730 399218 284966 399454
rect 284730 398898 284966 399134
rect 315450 399218 315686 399454
rect 315450 398898 315686 399134
rect 346170 399218 346406 399454
rect 346170 398898 346406 399134
rect 376890 399218 377126 399454
rect 376890 398898 377126 399134
rect 407610 399218 407846 399454
rect 407610 398898 407846 399134
rect 438330 399218 438566 399454
rect 438330 398898 438566 399134
rect 469050 399218 469286 399454
rect 469050 398898 469286 399134
rect 499770 399218 500006 399454
rect 499770 398898 500006 399134
rect 530490 399218 530726 399454
rect 530490 398898 530726 399134
rect 561210 399218 561446 399454
rect 561210 398898 561446 399134
rect 567266 388658 567502 388894
rect 567586 388658 567822 388894
rect 567266 388338 567502 388574
rect 567586 388338 567822 388574
rect 23610 381218 23846 381454
rect 23610 380898 23846 381134
rect 54330 381218 54566 381454
rect 54330 380898 54566 381134
rect 85050 381218 85286 381454
rect 85050 380898 85286 381134
rect 115770 381218 116006 381454
rect 115770 380898 116006 381134
rect 146490 381218 146726 381454
rect 146490 380898 146726 381134
rect 177210 381218 177446 381454
rect 177210 380898 177446 381134
rect 207930 381218 208166 381454
rect 207930 380898 208166 381134
rect 238650 381218 238886 381454
rect 238650 380898 238886 381134
rect 269370 381218 269606 381454
rect 269370 380898 269606 381134
rect 300090 381218 300326 381454
rect 300090 380898 300326 381134
rect 330810 381218 331046 381454
rect 330810 380898 331046 381134
rect 361530 381218 361766 381454
rect 361530 380898 361766 381134
rect 392250 381218 392486 381454
rect 392250 380898 392486 381134
rect 422970 381218 423206 381454
rect 422970 380898 423206 381134
rect 453690 381218 453926 381454
rect 453690 380898 453926 381134
rect 484410 381218 484646 381454
rect 484410 380898 484646 381134
rect 515130 381218 515366 381454
rect 515130 380898 515366 381134
rect 545850 381218 546086 381454
rect 545850 380898 546086 381134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect 8250 363218 8486 363454
rect 8250 362898 8486 363134
rect 38970 363218 39206 363454
rect 38970 362898 39206 363134
rect 69690 363218 69926 363454
rect 69690 362898 69926 363134
rect 100410 363218 100646 363454
rect 100410 362898 100646 363134
rect 131130 363218 131366 363454
rect 131130 362898 131366 363134
rect 161850 363218 162086 363454
rect 161850 362898 162086 363134
rect 192570 363218 192806 363454
rect 192570 362898 192806 363134
rect 223290 363218 223526 363454
rect 223290 362898 223526 363134
rect 254010 363218 254246 363454
rect 254010 362898 254246 363134
rect 284730 363218 284966 363454
rect 284730 362898 284966 363134
rect 315450 363218 315686 363454
rect 315450 362898 315686 363134
rect 346170 363218 346406 363454
rect 346170 362898 346406 363134
rect 376890 363218 377126 363454
rect 376890 362898 377126 363134
rect 407610 363218 407846 363454
rect 407610 362898 407846 363134
rect 438330 363218 438566 363454
rect 438330 362898 438566 363134
rect 469050 363218 469286 363454
rect 469050 362898 469286 363134
rect 499770 363218 500006 363454
rect 499770 362898 500006 363134
rect 530490 363218 530726 363454
rect 530490 362898 530726 363134
rect 561210 363218 561446 363454
rect 561210 362898 561446 363134
rect 567266 352658 567502 352894
rect 567586 352658 567822 352894
rect 567266 352338 567502 352574
rect 567586 352338 567822 352574
rect 23610 345218 23846 345454
rect 23610 344898 23846 345134
rect 54330 345218 54566 345454
rect 54330 344898 54566 345134
rect 85050 345218 85286 345454
rect 85050 344898 85286 345134
rect 115770 345218 116006 345454
rect 115770 344898 116006 345134
rect 146490 345218 146726 345454
rect 146490 344898 146726 345134
rect 177210 345218 177446 345454
rect 177210 344898 177446 345134
rect 207930 345218 208166 345454
rect 207930 344898 208166 345134
rect 238650 345218 238886 345454
rect 238650 344898 238886 345134
rect 269370 345218 269606 345454
rect 269370 344898 269606 345134
rect 300090 345218 300326 345454
rect 300090 344898 300326 345134
rect 330810 345218 331046 345454
rect 330810 344898 331046 345134
rect 361530 345218 361766 345454
rect 361530 344898 361766 345134
rect 392250 345218 392486 345454
rect 392250 344898 392486 345134
rect 422970 345218 423206 345454
rect 422970 344898 423206 345134
rect 453690 345218 453926 345454
rect 453690 344898 453926 345134
rect 484410 345218 484646 345454
rect 484410 344898 484646 345134
rect 515130 345218 515366 345454
rect 515130 344898 515366 345134
rect 545850 345218 546086 345454
rect 545850 344898 546086 345134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect 8250 327218 8486 327454
rect 8250 326898 8486 327134
rect 38970 327218 39206 327454
rect 38970 326898 39206 327134
rect 69690 327218 69926 327454
rect 69690 326898 69926 327134
rect 100410 327218 100646 327454
rect 100410 326898 100646 327134
rect 131130 327218 131366 327454
rect 131130 326898 131366 327134
rect 161850 327218 162086 327454
rect 161850 326898 162086 327134
rect 192570 327218 192806 327454
rect 192570 326898 192806 327134
rect 223290 327218 223526 327454
rect 223290 326898 223526 327134
rect 254010 327218 254246 327454
rect 254010 326898 254246 327134
rect 284730 327218 284966 327454
rect 284730 326898 284966 327134
rect 315450 327218 315686 327454
rect 315450 326898 315686 327134
rect 346170 327218 346406 327454
rect 346170 326898 346406 327134
rect 376890 327218 377126 327454
rect 376890 326898 377126 327134
rect 407610 327218 407846 327454
rect 407610 326898 407846 327134
rect 438330 327218 438566 327454
rect 438330 326898 438566 327134
rect 469050 327218 469286 327454
rect 469050 326898 469286 327134
rect 499770 327218 500006 327454
rect 499770 326898 500006 327134
rect 530490 327218 530726 327454
rect 530490 326898 530726 327134
rect 561210 327218 561446 327454
rect 561210 326898 561446 327134
rect 567266 316658 567502 316894
rect 567586 316658 567822 316894
rect 567266 316338 567502 316574
rect 567586 316338 567822 316574
rect 23610 309218 23846 309454
rect 23610 308898 23846 309134
rect 54330 309218 54566 309454
rect 54330 308898 54566 309134
rect 85050 309218 85286 309454
rect 85050 308898 85286 309134
rect 115770 309218 116006 309454
rect 115770 308898 116006 309134
rect 146490 309218 146726 309454
rect 146490 308898 146726 309134
rect 177210 309218 177446 309454
rect 177210 308898 177446 309134
rect 207930 309218 208166 309454
rect 207930 308898 208166 309134
rect 238650 309218 238886 309454
rect 238650 308898 238886 309134
rect 269370 309218 269606 309454
rect 269370 308898 269606 309134
rect 300090 309218 300326 309454
rect 300090 308898 300326 309134
rect 330810 309218 331046 309454
rect 330810 308898 331046 309134
rect 361530 309218 361766 309454
rect 361530 308898 361766 309134
rect 392250 309218 392486 309454
rect 392250 308898 392486 309134
rect 422970 309218 423206 309454
rect 422970 308898 423206 309134
rect 453690 309218 453926 309454
rect 453690 308898 453926 309134
rect 484410 309218 484646 309454
rect 484410 308898 484646 309134
rect 515130 309218 515366 309454
rect 515130 308898 515366 309134
rect 545850 309218 546086 309454
rect 545850 308898 546086 309134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect 8250 291218 8486 291454
rect 8250 290898 8486 291134
rect 38970 291218 39206 291454
rect 38970 290898 39206 291134
rect 69690 291218 69926 291454
rect 69690 290898 69926 291134
rect 100410 291218 100646 291454
rect 100410 290898 100646 291134
rect 131130 291218 131366 291454
rect 131130 290898 131366 291134
rect 161850 291218 162086 291454
rect 161850 290898 162086 291134
rect 192570 291218 192806 291454
rect 192570 290898 192806 291134
rect 223290 291218 223526 291454
rect 223290 290898 223526 291134
rect 254010 291218 254246 291454
rect 254010 290898 254246 291134
rect 284730 291218 284966 291454
rect 284730 290898 284966 291134
rect 315450 291218 315686 291454
rect 315450 290898 315686 291134
rect 346170 291218 346406 291454
rect 346170 290898 346406 291134
rect 376890 291218 377126 291454
rect 376890 290898 377126 291134
rect 407610 291218 407846 291454
rect 407610 290898 407846 291134
rect 438330 291218 438566 291454
rect 438330 290898 438566 291134
rect 469050 291218 469286 291454
rect 469050 290898 469286 291134
rect 499770 291218 500006 291454
rect 499770 290898 500006 291134
rect 530490 291218 530726 291454
rect 530490 290898 530726 291134
rect 561210 291218 561446 291454
rect 561210 290898 561446 291134
rect 567266 280658 567502 280894
rect 567586 280658 567822 280894
rect 567266 280338 567502 280574
rect 567586 280338 567822 280574
rect 23610 273218 23846 273454
rect 23610 272898 23846 273134
rect 54330 273218 54566 273454
rect 54330 272898 54566 273134
rect 85050 273218 85286 273454
rect 85050 272898 85286 273134
rect 115770 273218 116006 273454
rect 115770 272898 116006 273134
rect 146490 273218 146726 273454
rect 146490 272898 146726 273134
rect 177210 273218 177446 273454
rect 177210 272898 177446 273134
rect 207930 273218 208166 273454
rect 207930 272898 208166 273134
rect 238650 273218 238886 273454
rect 238650 272898 238886 273134
rect 269370 273218 269606 273454
rect 269370 272898 269606 273134
rect 300090 273218 300326 273454
rect 300090 272898 300326 273134
rect 330810 273218 331046 273454
rect 330810 272898 331046 273134
rect 361530 273218 361766 273454
rect 361530 272898 361766 273134
rect 392250 273218 392486 273454
rect 392250 272898 392486 273134
rect 422970 273218 423206 273454
rect 422970 272898 423206 273134
rect 453690 273218 453926 273454
rect 453690 272898 453926 273134
rect 484410 273218 484646 273454
rect 484410 272898 484646 273134
rect 515130 273218 515366 273454
rect 515130 272898 515366 273134
rect 545850 273218 546086 273454
rect 545850 272898 546086 273134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect 8250 255218 8486 255454
rect 8250 254898 8486 255134
rect 38970 255218 39206 255454
rect 38970 254898 39206 255134
rect 69690 255218 69926 255454
rect 69690 254898 69926 255134
rect 100410 255218 100646 255454
rect 100410 254898 100646 255134
rect 131130 255218 131366 255454
rect 131130 254898 131366 255134
rect 161850 255218 162086 255454
rect 161850 254898 162086 255134
rect 192570 255218 192806 255454
rect 192570 254898 192806 255134
rect 223290 255218 223526 255454
rect 223290 254898 223526 255134
rect 254010 255218 254246 255454
rect 254010 254898 254246 255134
rect 284730 255218 284966 255454
rect 284730 254898 284966 255134
rect 315450 255218 315686 255454
rect 315450 254898 315686 255134
rect 346170 255218 346406 255454
rect 346170 254898 346406 255134
rect 376890 255218 377126 255454
rect 376890 254898 377126 255134
rect 407610 255218 407846 255454
rect 407610 254898 407846 255134
rect 438330 255218 438566 255454
rect 438330 254898 438566 255134
rect 469050 255218 469286 255454
rect 469050 254898 469286 255134
rect 499770 255218 500006 255454
rect 499770 254898 500006 255134
rect 530490 255218 530726 255454
rect 530490 254898 530726 255134
rect 561210 255218 561446 255454
rect 561210 254898 561446 255134
rect 567266 244658 567502 244894
rect 567586 244658 567822 244894
rect 567266 244338 567502 244574
rect 567586 244338 567822 244574
rect 23610 237218 23846 237454
rect 23610 236898 23846 237134
rect 54330 237218 54566 237454
rect 54330 236898 54566 237134
rect 85050 237218 85286 237454
rect 85050 236898 85286 237134
rect 115770 237218 116006 237454
rect 115770 236898 116006 237134
rect 146490 237218 146726 237454
rect 146490 236898 146726 237134
rect 177210 237218 177446 237454
rect 177210 236898 177446 237134
rect 207930 237218 208166 237454
rect 207930 236898 208166 237134
rect 238650 237218 238886 237454
rect 238650 236898 238886 237134
rect 269370 237218 269606 237454
rect 269370 236898 269606 237134
rect 300090 237218 300326 237454
rect 300090 236898 300326 237134
rect 330810 237218 331046 237454
rect 330810 236898 331046 237134
rect 361530 237218 361766 237454
rect 361530 236898 361766 237134
rect 392250 237218 392486 237454
rect 392250 236898 392486 237134
rect 422970 237218 423206 237454
rect 422970 236898 423206 237134
rect 453690 237218 453926 237454
rect 453690 236898 453926 237134
rect 484410 237218 484646 237454
rect 484410 236898 484646 237134
rect 515130 237218 515366 237454
rect 515130 236898 515366 237134
rect 545850 237218 546086 237454
rect 545850 236898 546086 237134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect 8250 219218 8486 219454
rect 8250 218898 8486 219134
rect 38970 219218 39206 219454
rect 38970 218898 39206 219134
rect 69690 219218 69926 219454
rect 69690 218898 69926 219134
rect 100410 219218 100646 219454
rect 100410 218898 100646 219134
rect 131130 219218 131366 219454
rect 131130 218898 131366 219134
rect 161850 219218 162086 219454
rect 161850 218898 162086 219134
rect 192570 219218 192806 219454
rect 192570 218898 192806 219134
rect 223290 219218 223526 219454
rect 223290 218898 223526 219134
rect 254010 219218 254246 219454
rect 254010 218898 254246 219134
rect 284730 219218 284966 219454
rect 284730 218898 284966 219134
rect 315450 219218 315686 219454
rect 315450 218898 315686 219134
rect 346170 219218 346406 219454
rect 346170 218898 346406 219134
rect 376890 219218 377126 219454
rect 376890 218898 377126 219134
rect 407610 219218 407846 219454
rect 407610 218898 407846 219134
rect 438330 219218 438566 219454
rect 438330 218898 438566 219134
rect 469050 219218 469286 219454
rect 469050 218898 469286 219134
rect 499770 219218 500006 219454
rect 499770 218898 500006 219134
rect 530490 219218 530726 219454
rect 530490 218898 530726 219134
rect 561210 219218 561446 219454
rect 561210 218898 561446 219134
rect 567266 208658 567502 208894
rect 567586 208658 567822 208894
rect 567266 208338 567502 208574
rect 567586 208338 567822 208574
rect 23610 201218 23846 201454
rect 23610 200898 23846 201134
rect 54330 201218 54566 201454
rect 54330 200898 54566 201134
rect 85050 201218 85286 201454
rect 85050 200898 85286 201134
rect 115770 201218 116006 201454
rect 115770 200898 116006 201134
rect 146490 201218 146726 201454
rect 146490 200898 146726 201134
rect 177210 201218 177446 201454
rect 177210 200898 177446 201134
rect 207930 201218 208166 201454
rect 207930 200898 208166 201134
rect 238650 201218 238886 201454
rect 238650 200898 238886 201134
rect 269370 201218 269606 201454
rect 269370 200898 269606 201134
rect 300090 201218 300326 201454
rect 300090 200898 300326 201134
rect 330810 201218 331046 201454
rect 330810 200898 331046 201134
rect 361530 201218 361766 201454
rect 361530 200898 361766 201134
rect 392250 201218 392486 201454
rect 392250 200898 392486 201134
rect 422970 201218 423206 201454
rect 422970 200898 423206 201134
rect 453690 201218 453926 201454
rect 453690 200898 453926 201134
rect 484410 201218 484646 201454
rect 484410 200898 484646 201134
rect 515130 201218 515366 201454
rect 515130 200898 515366 201134
rect 545850 201218 546086 201454
rect 545850 200898 546086 201134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect 8250 183218 8486 183454
rect 8250 182898 8486 183134
rect 38970 183218 39206 183454
rect 38970 182898 39206 183134
rect 69690 183218 69926 183454
rect 69690 182898 69926 183134
rect 100410 183218 100646 183454
rect 100410 182898 100646 183134
rect 131130 183218 131366 183454
rect 131130 182898 131366 183134
rect 161850 183218 162086 183454
rect 161850 182898 162086 183134
rect 192570 183218 192806 183454
rect 192570 182898 192806 183134
rect 223290 183218 223526 183454
rect 223290 182898 223526 183134
rect 254010 183218 254246 183454
rect 254010 182898 254246 183134
rect 284730 183218 284966 183454
rect 284730 182898 284966 183134
rect 315450 183218 315686 183454
rect 315450 182898 315686 183134
rect 346170 183218 346406 183454
rect 346170 182898 346406 183134
rect 376890 183218 377126 183454
rect 376890 182898 377126 183134
rect 407610 183218 407846 183454
rect 407610 182898 407846 183134
rect 438330 183218 438566 183454
rect 438330 182898 438566 183134
rect 469050 183218 469286 183454
rect 469050 182898 469286 183134
rect 499770 183218 500006 183454
rect 499770 182898 500006 183134
rect 530490 183218 530726 183454
rect 530490 182898 530726 183134
rect 561210 183218 561446 183454
rect 561210 182898 561446 183134
rect 567266 172658 567502 172894
rect 567586 172658 567822 172894
rect 567266 172338 567502 172574
rect 567586 172338 567822 172574
rect 23610 165218 23846 165454
rect 23610 164898 23846 165134
rect 54330 165218 54566 165454
rect 54330 164898 54566 165134
rect 85050 165218 85286 165454
rect 85050 164898 85286 165134
rect 115770 165218 116006 165454
rect 115770 164898 116006 165134
rect 146490 165218 146726 165454
rect 146490 164898 146726 165134
rect 177210 165218 177446 165454
rect 177210 164898 177446 165134
rect 207930 165218 208166 165454
rect 207930 164898 208166 165134
rect 238650 165218 238886 165454
rect 238650 164898 238886 165134
rect 269370 165218 269606 165454
rect 269370 164898 269606 165134
rect 300090 165218 300326 165454
rect 300090 164898 300326 165134
rect 330810 165218 331046 165454
rect 330810 164898 331046 165134
rect 361530 165218 361766 165454
rect 361530 164898 361766 165134
rect 392250 165218 392486 165454
rect 392250 164898 392486 165134
rect 422970 165218 423206 165454
rect 422970 164898 423206 165134
rect 453690 165218 453926 165454
rect 453690 164898 453926 165134
rect 484410 165218 484646 165454
rect 484410 164898 484646 165134
rect 515130 165218 515366 165454
rect 515130 164898 515366 165134
rect 545850 165218 546086 165454
rect 545850 164898 546086 165134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect 8250 147218 8486 147454
rect 8250 146898 8486 147134
rect 38970 147218 39206 147454
rect 38970 146898 39206 147134
rect 69690 147218 69926 147454
rect 69690 146898 69926 147134
rect 100410 147218 100646 147454
rect 100410 146898 100646 147134
rect 131130 147218 131366 147454
rect 131130 146898 131366 147134
rect 161850 147218 162086 147454
rect 161850 146898 162086 147134
rect 192570 147218 192806 147454
rect 192570 146898 192806 147134
rect 223290 147218 223526 147454
rect 223290 146898 223526 147134
rect 254010 147218 254246 147454
rect 254010 146898 254246 147134
rect 284730 147218 284966 147454
rect 284730 146898 284966 147134
rect 315450 147218 315686 147454
rect 315450 146898 315686 147134
rect 346170 147218 346406 147454
rect 346170 146898 346406 147134
rect 376890 147218 377126 147454
rect 376890 146898 377126 147134
rect 407610 147218 407846 147454
rect 407610 146898 407846 147134
rect 438330 147218 438566 147454
rect 438330 146898 438566 147134
rect 469050 147218 469286 147454
rect 469050 146898 469286 147134
rect 499770 147218 500006 147454
rect 499770 146898 500006 147134
rect 530490 147218 530726 147454
rect 530490 146898 530726 147134
rect 561210 147218 561446 147454
rect 561210 146898 561446 147134
rect 567266 136658 567502 136894
rect 567586 136658 567822 136894
rect 567266 136338 567502 136574
rect 567586 136338 567822 136574
rect 23610 129218 23846 129454
rect 23610 128898 23846 129134
rect 54330 129218 54566 129454
rect 54330 128898 54566 129134
rect 85050 129218 85286 129454
rect 85050 128898 85286 129134
rect 115770 129218 116006 129454
rect 115770 128898 116006 129134
rect 146490 129218 146726 129454
rect 146490 128898 146726 129134
rect 177210 129218 177446 129454
rect 177210 128898 177446 129134
rect 207930 129218 208166 129454
rect 207930 128898 208166 129134
rect 238650 129218 238886 129454
rect 238650 128898 238886 129134
rect 269370 129218 269606 129454
rect 269370 128898 269606 129134
rect 300090 129218 300326 129454
rect 300090 128898 300326 129134
rect 330810 129218 331046 129454
rect 330810 128898 331046 129134
rect 361530 129218 361766 129454
rect 361530 128898 361766 129134
rect 392250 129218 392486 129454
rect 392250 128898 392486 129134
rect 422970 129218 423206 129454
rect 422970 128898 423206 129134
rect 453690 129218 453926 129454
rect 453690 128898 453926 129134
rect 484410 129218 484646 129454
rect 484410 128898 484646 129134
rect 515130 129218 515366 129454
rect 515130 128898 515366 129134
rect 545850 129218 546086 129454
rect 545850 128898 546086 129134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect 8250 111218 8486 111454
rect 8250 110898 8486 111134
rect 38970 111218 39206 111454
rect 38970 110898 39206 111134
rect 69690 111218 69926 111454
rect 69690 110898 69926 111134
rect 100410 111218 100646 111454
rect 100410 110898 100646 111134
rect 131130 111218 131366 111454
rect 131130 110898 131366 111134
rect 161850 111218 162086 111454
rect 161850 110898 162086 111134
rect 192570 111218 192806 111454
rect 192570 110898 192806 111134
rect 223290 111218 223526 111454
rect 223290 110898 223526 111134
rect 254010 111218 254246 111454
rect 254010 110898 254246 111134
rect 284730 111218 284966 111454
rect 284730 110898 284966 111134
rect 315450 111218 315686 111454
rect 315450 110898 315686 111134
rect 346170 111218 346406 111454
rect 346170 110898 346406 111134
rect 376890 111218 377126 111454
rect 376890 110898 377126 111134
rect 407610 111218 407846 111454
rect 407610 110898 407846 111134
rect 438330 111218 438566 111454
rect 438330 110898 438566 111134
rect 469050 111218 469286 111454
rect 469050 110898 469286 111134
rect 499770 111218 500006 111454
rect 499770 110898 500006 111134
rect 530490 111218 530726 111454
rect 530490 110898 530726 111134
rect 561210 111218 561446 111454
rect 561210 110898 561446 111134
rect 567266 100658 567502 100894
rect 567586 100658 567822 100894
rect 567266 100338 567502 100574
rect 567586 100338 567822 100574
rect 23610 93218 23846 93454
rect 23610 92898 23846 93134
rect 54330 93218 54566 93454
rect 54330 92898 54566 93134
rect 85050 93218 85286 93454
rect 85050 92898 85286 93134
rect 115770 93218 116006 93454
rect 115770 92898 116006 93134
rect 146490 93218 146726 93454
rect 146490 92898 146726 93134
rect 177210 93218 177446 93454
rect 177210 92898 177446 93134
rect 207930 93218 208166 93454
rect 207930 92898 208166 93134
rect 238650 93218 238886 93454
rect 238650 92898 238886 93134
rect 269370 93218 269606 93454
rect 269370 92898 269606 93134
rect 300090 93218 300326 93454
rect 300090 92898 300326 93134
rect 330810 93218 331046 93454
rect 330810 92898 331046 93134
rect 361530 93218 361766 93454
rect 361530 92898 361766 93134
rect 392250 93218 392486 93454
rect 392250 92898 392486 93134
rect 422970 93218 423206 93454
rect 422970 92898 423206 93134
rect 453690 93218 453926 93454
rect 453690 92898 453926 93134
rect 484410 93218 484646 93454
rect 484410 92898 484646 93134
rect 515130 93218 515366 93454
rect 515130 92898 515366 93134
rect 545850 93218 546086 93454
rect 545850 92898 546086 93134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect 8250 75218 8486 75454
rect 8250 74898 8486 75134
rect 38970 75218 39206 75454
rect 38970 74898 39206 75134
rect 69690 75218 69926 75454
rect 69690 74898 69926 75134
rect 100410 75218 100646 75454
rect 100410 74898 100646 75134
rect 131130 75218 131366 75454
rect 131130 74898 131366 75134
rect 161850 75218 162086 75454
rect 161850 74898 162086 75134
rect 192570 75218 192806 75454
rect 192570 74898 192806 75134
rect 223290 75218 223526 75454
rect 223290 74898 223526 75134
rect 254010 75218 254246 75454
rect 254010 74898 254246 75134
rect 284730 75218 284966 75454
rect 284730 74898 284966 75134
rect 315450 75218 315686 75454
rect 315450 74898 315686 75134
rect 346170 75218 346406 75454
rect 346170 74898 346406 75134
rect 376890 75218 377126 75454
rect 376890 74898 377126 75134
rect 407610 75218 407846 75454
rect 407610 74898 407846 75134
rect 438330 75218 438566 75454
rect 438330 74898 438566 75134
rect 469050 75218 469286 75454
rect 469050 74898 469286 75134
rect 499770 75218 500006 75454
rect 499770 74898 500006 75134
rect 530490 75218 530726 75454
rect 530490 74898 530726 75134
rect 561210 75218 561446 75454
rect 561210 74898 561446 75134
rect 567266 64658 567502 64894
rect 567586 64658 567822 64894
rect 567266 64338 567502 64574
rect 567586 64338 567822 64574
rect 23610 57218 23846 57454
rect 23610 56898 23846 57134
rect 54330 57218 54566 57454
rect 54330 56898 54566 57134
rect 85050 57218 85286 57454
rect 85050 56898 85286 57134
rect 115770 57218 116006 57454
rect 115770 56898 116006 57134
rect 146490 57218 146726 57454
rect 146490 56898 146726 57134
rect 177210 57218 177446 57454
rect 177210 56898 177446 57134
rect 207930 57218 208166 57454
rect 207930 56898 208166 57134
rect 238650 57218 238886 57454
rect 238650 56898 238886 57134
rect 269370 57218 269606 57454
rect 269370 56898 269606 57134
rect 300090 57218 300326 57454
rect 300090 56898 300326 57134
rect 330810 57218 331046 57454
rect 330810 56898 331046 57134
rect 361530 57218 361766 57454
rect 361530 56898 361766 57134
rect 392250 57218 392486 57454
rect 392250 56898 392486 57134
rect 422970 57218 423206 57454
rect 422970 56898 423206 57134
rect 453690 57218 453926 57454
rect 453690 56898 453926 57134
rect 484410 57218 484646 57454
rect 484410 56898 484646 57134
rect 515130 57218 515366 57454
rect 515130 56898 515366 57134
rect 545850 57218 546086 57454
rect 545850 56898 546086 57134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect 8250 39218 8486 39454
rect 8250 38898 8486 39134
rect 38970 39218 39206 39454
rect 38970 38898 39206 39134
rect 69690 39218 69926 39454
rect 69690 38898 69926 39134
rect 100410 39218 100646 39454
rect 100410 38898 100646 39134
rect 131130 39218 131366 39454
rect 131130 38898 131366 39134
rect 161850 39218 162086 39454
rect 161850 38898 162086 39134
rect 192570 39218 192806 39454
rect 192570 38898 192806 39134
rect 223290 39218 223526 39454
rect 223290 38898 223526 39134
rect 254010 39218 254246 39454
rect 254010 38898 254246 39134
rect 284730 39218 284966 39454
rect 284730 38898 284966 39134
rect 315450 39218 315686 39454
rect 315450 38898 315686 39134
rect 346170 39218 346406 39454
rect 346170 38898 346406 39134
rect 376890 39218 377126 39454
rect 376890 38898 377126 39134
rect 407610 39218 407846 39454
rect 407610 38898 407846 39134
rect 438330 39218 438566 39454
rect 438330 38898 438566 39134
rect 469050 39218 469286 39454
rect 469050 38898 469286 39134
rect 499770 39218 500006 39454
rect 499770 38898 500006 39134
rect 530490 39218 530726 39454
rect 530490 38898 530726 39134
rect 561210 39218 561446 39454
rect 561210 38898 561446 39134
rect 567266 28658 567502 28894
rect 567586 28658 567822 28894
rect 567266 28338 567502 28574
rect 567586 28338 567822 28574
rect 23610 21218 23846 21454
rect 23610 20898 23846 21134
rect 54330 21218 54566 21454
rect 54330 20898 54566 21134
rect 85050 21218 85286 21454
rect 85050 20898 85286 21134
rect 115770 21218 116006 21454
rect 115770 20898 116006 21134
rect 146490 21218 146726 21454
rect 146490 20898 146726 21134
rect 177210 21218 177446 21454
rect 177210 20898 177446 21134
rect 207930 21218 208166 21454
rect 207930 20898 208166 21134
rect 238650 21218 238886 21454
rect 238650 20898 238886 21134
rect 269370 21218 269606 21454
rect 269370 20898 269606 21134
rect 300090 21218 300326 21454
rect 300090 20898 300326 21134
rect 330810 21218 331046 21454
rect 330810 20898 331046 21134
rect 361530 21218 361766 21454
rect 361530 20898 361766 21134
rect 392250 21218 392486 21454
rect 392250 20898 392486 21134
rect 422970 21218 423206 21454
rect 422970 20898 423206 21134
rect 453690 21218 453926 21454
rect 453690 20898 453926 21134
rect 484410 21218 484646 21454
rect 484410 20898 484646 21134
rect 515130 21218 515366 21454
rect 515130 20898 515366 21134
rect 545850 21218 546086 21454
rect 545850 20898 546086 21134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect 8250 3218 8486 3454
rect 8250 2898 8486 3134
rect 38970 3218 39206 3454
rect 38970 2898 39206 3134
rect 69690 3218 69926 3454
rect 69690 2898 69926 3134
rect 100410 3218 100646 3454
rect 100410 2898 100646 3134
rect 131130 3218 131366 3454
rect 131130 2898 131366 3134
rect 161850 3218 162086 3454
rect 161850 2898 162086 3134
rect 192570 3218 192806 3454
rect 192570 2898 192806 3134
rect 223290 3218 223526 3454
rect 223290 2898 223526 3134
rect 254010 3218 254246 3454
rect 254010 2898 254246 3134
rect 284730 3218 284966 3454
rect 284730 2898 284966 3134
rect 315450 3218 315686 3454
rect 315450 2898 315686 3134
rect 346170 3218 346406 3454
rect 346170 2898 346406 3134
rect 376890 3218 377126 3454
rect 376890 2898 377126 3134
rect 407610 3218 407846 3454
rect 407610 2898 407846 3134
rect 438330 3218 438566 3454
rect 438330 2898 438566 3134
rect 469050 3218 469286 3454
rect 469050 2898 469286 3134
rect 499770 3218 500006 3454
rect 499770 2898 500006 3134
rect 530490 3218 530726 3454
rect 530490 2898 530726 3134
rect 561210 3218 561446 3454
rect 561210 2898 561446 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 5546 -2502 5782 -2266
rect 5866 -2502 6102 -2266
rect 5546 -2822 5782 -2586
rect 5866 -2822 6102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 9266 -4422 9502 -4186
rect 9586 -4422 9822 -4186
rect 9266 -4742 9502 -4506
rect 9586 -4742 9822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 23546 -3462 23782 -3226
rect 23866 -3462 24102 -3226
rect 23546 -3782 23782 -3546
rect 23866 -3782 24102 -3546
rect 27266 -5382 27502 -5146
rect 27586 -5382 27822 -5146
rect 27266 -5702 27502 -5466
rect 27586 -5702 27822 -5466
rect 12986 -6342 13222 -6106
rect 13306 -6342 13542 -6106
rect 12986 -6662 13222 -6426
rect 13306 -6662 13542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 41546 -2502 41782 -2266
rect 41866 -2502 42102 -2266
rect 41546 -2822 41782 -2586
rect 41866 -2822 42102 -2586
rect 45266 -4422 45502 -4186
rect 45586 -4422 45822 -4186
rect 45266 -4742 45502 -4506
rect 45586 -4742 45822 -4506
rect 30986 -7302 31222 -7066
rect 31306 -7302 31542 -7066
rect 30986 -7622 31222 -7386
rect 31306 -7622 31542 -7386
rect 59546 -3462 59782 -3226
rect 59866 -3462 60102 -3226
rect 59546 -3782 59782 -3546
rect 59866 -3782 60102 -3546
rect 63266 -5382 63502 -5146
rect 63586 -5382 63822 -5146
rect 63266 -5702 63502 -5466
rect 63586 -5702 63822 -5466
rect 48986 -6342 49222 -6106
rect 49306 -6342 49542 -6106
rect 48986 -6662 49222 -6426
rect 49306 -6662 49542 -6426
rect 77546 -2502 77782 -2266
rect 77866 -2502 78102 -2266
rect 77546 -2822 77782 -2586
rect 77866 -2822 78102 -2586
rect 81266 -4422 81502 -4186
rect 81586 -4422 81822 -4186
rect 81266 -4742 81502 -4506
rect 81586 -4742 81822 -4506
rect 66986 -7302 67222 -7066
rect 67306 -7302 67542 -7066
rect 66986 -7622 67222 -7386
rect 67306 -7622 67542 -7386
rect 95546 -3462 95782 -3226
rect 95866 -3462 96102 -3226
rect 95546 -3782 95782 -3546
rect 95866 -3782 96102 -3546
rect 99266 -5382 99502 -5146
rect 99586 -5382 99822 -5146
rect 99266 -5702 99502 -5466
rect 99586 -5702 99822 -5466
rect 84986 -6342 85222 -6106
rect 85306 -6342 85542 -6106
rect 84986 -6662 85222 -6426
rect 85306 -6662 85542 -6426
rect 113546 -2502 113782 -2266
rect 113866 -2502 114102 -2266
rect 113546 -2822 113782 -2586
rect 113866 -2822 114102 -2586
rect 117266 -4422 117502 -4186
rect 117586 -4422 117822 -4186
rect 117266 -4742 117502 -4506
rect 117586 -4742 117822 -4506
rect 102986 -7302 103222 -7066
rect 103306 -7302 103542 -7066
rect 102986 -7622 103222 -7386
rect 103306 -7622 103542 -7386
rect 131546 -3462 131782 -3226
rect 131866 -3462 132102 -3226
rect 131546 -3782 131782 -3546
rect 131866 -3782 132102 -3546
rect 135266 -5382 135502 -5146
rect 135586 -5382 135822 -5146
rect 135266 -5702 135502 -5466
rect 135586 -5702 135822 -5466
rect 120986 -6342 121222 -6106
rect 121306 -6342 121542 -6106
rect 120986 -6662 121222 -6426
rect 121306 -6662 121542 -6426
rect 149546 -2502 149782 -2266
rect 149866 -2502 150102 -2266
rect 149546 -2822 149782 -2586
rect 149866 -2822 150102 -2586
rect 153266 -4422 153502 -4186
rect 153586 -4422 153822 -4186
rect 153266 -4742 153502 -4506
rect 153586 -4742 153822 -4506
rect 138986 -7302 139222 -7066
rect 139306 -7302 139542 -7066
rect 138986 -7622 139222 -7386
rect 139306 -7622 139542 -7386
rect 167546 -3462 167782 -3226
rect 167866 -3462 168102 -3226
rect 167546 -3782 167782 -3546
rect 167866 -3782 168102 -3546
rect 171266 -5382 171502 -5146
rect 171586 -5382 171822 -5146
rect 171266 -5702 171502 -5466
rect 171586 -5702 171822 -5466
rect 156986 -6342 157222 -6106
rect 157306 -6342 157542 -6106
rect 156986 -6662 157222 -6426
rect 157306 -6662 157542 -6426
rect 185546 -2502 185782 -2266
rect 185866 -2502 186102 -2266
rect 185546 -2822 185782 -2586
rect 185866 -2822 186102 -2586
rect 189266 -4422 189502 -4186
rect 189586 -4422 189822 -4186
rect 189266 -4742 189502 -4506
rect 189586 -4742 189822 -4506
rect 174986 -7302 175222 -7066
rect 175306 -7302 175542 -7066
rect 174986 -7622 175222 -7386
rect 175306 -7622 175542 -7386
rect 203546 -3462 203782 -3226
rect 203866 -3462 204102 -3226
rect 203546 -3782 203782 -3546
rect 203866 -3782 204102 -3546
rect 207266 -5382 207502 -5146
rect 207586 -5382 207822 -5146
rect 207266 -5702 207502 -5466
rect 207586 -5702 207822 -5466
rect 192986 -6342 193222 -6106
rect 193306 -6342 193542 -6106
rect 192986 -6662 193222 -6426
rect 193306 -6662 193542 -6426
rect 221546 -2502 221782 -2266
rect 221866 -2502 222102 -2266
rect 221546 -2822 221782 -2586
rect 221866 -2822 222102 -2586
rect 225266 -4422 225502 -4186
rect 225586 -4422 225822 -4186
rect 225266 -4742 225502 -4506
rect 225586 -4742 225822 -4506
rect 210986 -7302 211222 -7066
rect 211306 -7302 211542 -7066
rect 210986 -7622 211222 -7386
rect 211306 -7622 211542 -7386
rect 239546 -3462 239782 -3226
rect 239866 -3462 240102 -3226
rect 239546 -3782 239782 -3546
rect 239866 -3782 240102 -3546
rect 243266 -5382 243502 -5146
rect 243586 -5382 243822 -5146
rect 243266 -5702 243502 -5466
rect 243586 -5702 243822 -5466
rect 228986 -6342 229222 -6106
rect 229306 -6342 229542 -6106
rect 228986 -6662 229222 -6426
rect 229306 -6662 229542 -6426
rect 257546 -2502 257782 -2266
rect 257866 -2502 258102 -2266
rect 257546 -2822 257782 -2586
rect 257866 -2822 258102 -2586
rect 261266 -4422 261502 -4186
rect 261586 -4422 261822 -4186
rect 261266 -4742 261502 -4506
rect 261586 -4742 261822 -4506
rect 246986 -7302 247222 -7066
rect 247306 -7302 247542 -7066
rect 246986 -7622 247222 -7386
rect 247306 -7622 247542 -7386
rect 275546 -3462 275782 -3226
rect 275866 -3462 276102 -3226
rect 275546 -3782 275782 -3546
rect 275866 -3782 276102 -3546
rect 279266 -5382 279502 -5146
rect 279586 -5382 279822 -5146
rect 279266 -5702 279502 -5466
rect 279586 -5702 279822 -5466
rect 264986 -6342 265222 -6106
rect 265306 -6342 265542 -6106
rect 264986 -6662 265222 -6426
rect 265306 -6662 265542 -6426
rect 293546 -2502 293782 -2266
rect 293866 -2502 294102 -2266
rect 293546 -2822 293782 -2586
rect 293866 -2822 294102 -2586
rect 297266 -4422 297502 -4186
rect 297586 -4422 297822 -4186
rect 297266 -4742 297502 -4506
rect 297586 -4742 297822 -4506
rect 282986 -7302 283222 -7066
rect 283306 -7302 283542 -7066
rect 282986 -7622 283222 -7386
rect 283306 -7622 283542 -7386
rect 311546 -3462 311782 -3226
rect 311866 -3462 312102 -3226
rect 311546 -3782 311782 -3546
rect 311866 -3782 312102 -3546
rect 315266 -5382 315502 -5146
rect 315586 -5382 315822 -5146
rect 315266 -5702 315502 -5466
rect 315586 -5702 315822 -5466
rect 300986 -6342 301222 -6106
rect 301306 -6342 301542 -6106
rect 300986 -6662 301222 -6426
rect 301306 -6662 301542 -6426
rect 329546 -2502 329782 -2266
rect 329866 -2502 330102 -2266
rect 329546 -2822 329782 -2586
rect 329866 -2822 330102 -2586
rect 333266 -4422 333502 -4186
rect 333586 -4422 333822 -4186
rect 333266 -4742 333502 -4506
rect 333586 -4742 333822 -4506
rect 318986 -7302 319222 -7066
rect 319306 -7302 319542 -7066
rect 318986 -7622 319222 -7386
rect 319306 -7622 319542 -7386
rect 347546 -3462 347782 -3226
rect 347866 -3462 348102 -3226
rect 347546 -3782 347782 -3546
rect 347866 -3782 348102 -3546
rect 351266 -5382 351502 -5146
rect 351586 -5382 351822 -5146
rect 351266 -5702 351502 -5466
rect 351586 -5702 351822 -5466
rect 336986 -6342 337222 -6106
rect 337306 -6342 337542 -6106
rect 336986 -6662 337222 -6426
rect 337306 -6662 337542 -6426
rect 365546 -2502 365782 -2266
rect 365866 -2502 366102 -2266
rect 365546 -2822 365782 -2586
rect 365866 -2822 366102 -2586
rect 369266 -4422 369502 -4186
rect 369586 -4422 369822 -4186
rect 369266 -4742 369502 -4506
rect 369586 -4742 369822 -4506
rect 354986 -7302 355222 -7066
rect 355306 -7302 355542 -7066
rect 354986 -7622 355222 -7386
rect 355306 -7622 355542 -7386
rect 383546 -3462 383782 -3226
rect 383866 -3462 384102 -3226
rect 383546 -3782 383782 -3546
rect 383866 -3782 384102 -3546
rect 387266 -5382 387502 -5146
rect 387586 -5382 387822 -5146
rect 387266 -5702 387502 -5466
rect 387586 -5702 387822 -5466
rect 372986 -6342 373222 -6106
rect 373306 -6342 373542 -6106
rect 372986 -6662 373222 -6426
rect 373306 -6662 373542 -6426
rect 401546 -2502 401782 -2266
rect 401866 -2502 402102 -2266
rect 401546 -2822 401782 -2586
rect 401866 -2822 402102 -2586
rect 405266 -4422 405502 -4186
rect 405586 -4422 405822 -4186
rect 405266 -4742 405502 -4506
rect 405586 -4742 405822 -4506
rect 390986 -7302 391222 -7066
rect 391306 -7302 391542 -7066
rect 390986 -7622 391222 -7386
rect 391306 -7622 391542 -7386
rect 419546 -3462 419782 -3226
rect 419866 -3462 420102 -3226
rect 419546 -3782 419782 -3546
rect 419866 -3782 420102 -3546
rect 423266 -5382 423502 -5146
rect 423586 -5382 423822 -5146
rect 423266 -5702 423502 -5466
rect 423586 -5702 423822 -5466
rect 408986 -6342 409222 -6106
rect 409306 -6342 409542 -6106
rect 408986 -6662 409222 -6426
rect 409306 -6662 409542 -6426
rect 437546 -2502 437782 -2266
rect 437866 -2502 438102 -2266
rect 437546 -2822 437782 -2586
rect 437866 -2822 438102 -2586
rect 441266 -4422 441502 -4186
rect 441586 -4422 441822 -4186
rect 441266 -4742 441502 -4506
rect 441586 -4742 441822 -4506
rect 426986 -7302 427222 -7066
rect 427306 -7302 427542 -7066
rect 426986 -7622 427222 -7386
rect 427306 -7622 427542 -7386
rect 455546 -3462 455782 -3226
rect 455866 -3462 456102 -3226
rect 455546 -3782 455782 -3546
rect 455866 -3782 456102 -3546
rect 459266 -5382 459502 -5146
rect 459586 -5382 459822 -5146
rect 459266 -5702 459502 -5466
rect 459586 -5702 459822 -5466
rect 444986 -6342 445222 -6106
rect 445306 -6342 445542 -6106
rect 444986 -6662 445222 -6426
rect 445306 -6662 445542 -6426
rect 473546 -2502 473782 -2266
rect 473866 -2502 474102 -2266
rect 473546 -2822 473782 -2586
rect 473866 -2822 474102 -2586
rect 477266 -4422 477502 -4186
rect 477586 -4422 477822 -4186
rect 477266 -4742 477502 -4506
rect 477586 -4742 477822 -4506
rect 462986 -7302 463222 -7066
rect 463306 -7302 463542 -7066
rect 462986 -7622 463222 -7386
rect 463306 -7622 463542 -7386
rect 491546 -3462 491782 -3226
rect 491866 -3462 492102 -3226
rect 491546 -3782 491782 -3546
rect 491866 -3782 492102 -3546
rect 495266 -5382 495502 -5146
rect 495586 -5382 495822 -5146
rect 495266 -5702 495502 -5466
rect 495586 -5702 495822 -5466
rect 480986 -6342 481222 -6106
rect 481306 -6342 481542 -6106
rect 480986 -6662 481222 -6426
rect 481306 -6662 481542 -6426
rect 509546 -2502 509782 -2266
rect 509866 -2502 510102 -2266
rect 509546 -2822 509782 -2586
rect 509866 -2822 510102 -2586
rect 513266 -4422 513502 -4186
rect 513586 -4422 513822 -4186
rect 513266 -4742 513502 -4506
rect 513586 -4742 513822 -4506
rect 498986 -7302 499222 -7066
rect 499306 -7302 499542 -7066
rect 498986 -7622 499222 -7386
rect 499306 -7622 499542 -7386
rect 527546 -3462 527782 -3226
rect 527866 -3462 528102 -3226
rect 527546 -3782 527782 -3546
rect 527866 -3782 528102 -3546
rect 531266 -5382 531502 -5146
rect 531586 -5382 531822 -5146
rect 531266 -5702 531502 -5466
rect 531586 -5702 531822 -5466
rect 516986 -6342 517222 -6106
rect 517306 -6342 517542 -6106
rect 516986 -6662 517222 -6426
rect 517306 -6662 517542 -6426
rect 545546 -2502 545782 -2266
rect 545866 -2502 546102 -2266
rect 545546 -2822 545782 -2586
rect 545866 -2822 546102 -2586
rect 549266 -4422 549502 -4186
rect 549586 -4422 549822 -4186
rect 549266 -4742 549502 -4506
rect 549586 -4742 549822 -4506
rect 534986 -7302 535222 -7066
rect 535306 -7302 535542 -7066
rect 534986 -7622 535222 -7386
rect 535306 -7622 535542 -7386
rect 563546 -3462 563782 -3226
rect 563866 -3462 564102 -3226
rect 563546 -3782 563782 -3546
rect 563866 -3782 564102 -3546
rect 567266 -5382 567502 -5146
rect 567586 -5382 567822 -5146
rect 567266 -5702 567502 -5466
rect 567586 -5702 567822 -5466
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 581546 706522 581782 706758
rect 581866 706522 582102 706758
rect 581546 706202 581782 706438
rect 581866 706202 582102 706438
rect 570986 680378 571222 680614
rect 571306 680378 571542 680614
rect 570986 680058 571222 680294
rect 571306 680058 571542 680294
rect 570986 644378 571222 644614
rect 571306 644378 571542 644614
rect 570986 644058 571222 644294
rect 571306 644058 571542 644294
rect 570986 608378 571222 608614
rect 571306 608378 571542 608614
rect 570986 608058 571222 608294
rect 571306 608058 571542 608294
rect 570986 572378 571222 572614
rect 571306 572378 571542 572614
rect 570986 572058 571222 572294
rect 571306 572058 571542 572294
rect 570986 536378 571222 536614
rect 571306 536378 571542 536614
rect 570986 536058 571222 536294
rect 571306 536058 571542 536294
rect 570986 500378 571222 500614
rect 571306 500378 571542 500614
rect 570986 500058 571222 500294
rect 571306 500058 571542 500294
rect 570986 464378 571222 464614
rect 571306 464378 571542 464614
rect 570986 464058 571222 464294
rect 571306 464058 571542 464294
rect 570986 428378 571222 428614
rect 571306 428378 571542 428614
rect 570986 428058 571222 428294
rect 571306 428058 571542 428294
rect 570986 392378 571222 392614
rect 571306 392378 571542 392614
rect 570986 392058 571222 392294
rect 571306 392058 571542 392294
rect 570986 356378 571222 356614
rect 571306 356378 571542 356614
rect 570986 356058 571222 356294
rect 571306 356058 571542 356294
rect 570986 320378 571222 320614
rect 571306 320378 571542 320614
rect 570986 320058 571222 320294
rect 571306 320058 571542 320294
rect 570986 284378 571222 284614
rect 571306 284378 571542 284614
rect 570986 284058 571222 284294
rect 571306 284058 571542 284294
rect 570986 248378 571222 248614
rect 571306 248378 571542 248614
rect 570986 248058 571222 248294
rect 571306 248058 571542 248294
rect 570986 212378 571222 212614
rect 571306 212378 571542 212614
rect 570986 212058 571222 212294
rect 571306 212058 571542 212294
rect 570986 176378 571222 176614
rect 571306 176378 571542 176614
rect 570986 176058 571222 176294
rect 571306 176058 571542 176294
rect 570986 140378 571222 140614
rect 571306 140378 571542 140614
rect 570986 140058 571222 140294
rect 571306 140058 571542 140294
rect 570986 104378 571222 104614
rect 571306 104378 571542 104614
rect 570986 104058 571222 104294
rect 571306 104058 571542 104294
rect 570986 68378 571222 68614
rect 571306 68378 571542 68614
rect 570986 68058 571222 68294
rect 571306 68058 571542 68294
rect 570986 32378 571222 32614
rect 571306 32378 571542 32614
rect 570986 32058 571222 32294
rect 571306 32058 571542 32294
rect 552986 -6342 553222 -6106
rect 553306 -6342 553542 -6106
rect 552986 -6662 553222 -6426
rect 553306 -6662 553542 -6426
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 690938 587498 691174
rect 587582 690938 587818 691174
rect 587262 690618 587498 690854
rect 587582 690618 587818 690854
rect 587262 654938 587498 655174
rect 587582 654938 587818 655174
rect 587262 654618 587498 654854
rect 587582 654618 587818 654854
rect 587262 618938 587498 619174
rect 587582 618938 587818 619174
rect 587262 618618 587498 618854
rect 587582 618618 587818 618854
rect 587262 582938 587498 583174
rect 587582 582938 587818 583174
rect 587262 582618 587498 582854
rect 587582 582618 587818 582854
rect 587262 546938 587498 547174
rect 587582 546938 587818 547174
rect 587262 546618 587498 546854
rect 587582 546618 587818 546854
rect 587262 510938 587498 511174
rect 587582 510938 587818 511174
rect 587262 510618 587498 510854
rect 587582 510618 587818 510854
rect 587262 474938 587498 475174
rect 587582 474938 587818 475174
rect 587262 474618 587498 474854
rect 587582 474618 587818 474854
rect 587262 438938 587498 439174
rect 587582 438938 587818 439174
rect 587262 438618 587498 438854
rect 587582 438618 587818 438854
rect 587262 402938 587498 403174
rect 587582 402938 587818 403174
rect 587262 402618 587498 402854
rect 587582 402618 587818 402854
rect 587262 366938 587498 367174
rect 587582 366938 587818 367174
rect 587262 366618 587498 366854
rect 587582 366618 587818 366854
rect 587262 330938 587498 331174
rect 587582 330938 587818 331174
rect 587262 330618 587498 330854
rect 587582 330618 587818 330854
rect 587262 294938 587498 295174
rect 587582 294938 587818 295174
rect 587262 294618 587498 294854
rect 587582 294618 587818 294854
rect 587262 258938 587498 259174
rect 587582 258938 587818 259174
rect 587262 258618 587498 258854
rect 587582 258618 587818 258854
rect 587262 222938 587498 223174
rect 587582 222938 587818 223174
rect 587262 222618 587498 222854
rect 587582 222618 587818 222854
rect 587262 186938 587498 187174
rect 587582 186938 587818 187174
rect 587262 186618 587498 186854
rect 587582 186618 587818 186854
rect 587262 150938 587498 151174
rect 587582 150938 587818 151174
rect 587262 150618 587498 150854
rect 587582 150618 587818 150854
rect 587262 114938 587498 115174
rect 587582 114938 587818 115174
rect 587262 114618 587498 114854
rect 587582 114618 587818 114854
rect 587262 78938 587498 79174
rect 587582 78938 587818 79174
rect 587262 78618 587498 78854
rect 587582 78618 587818 78854
rect 587262 42938 587498 43174
rect 587582 42938 587818 43174
rect 587262 42618 587498 42854
rect 587582 42618 587818 42854
rect 587262 6938 587498 7174
rect 587582 6938 587818 7174
rect 587262 6618 587498 6854
rect 587582 6618 587818 6854
rect 581546 -2502 581782 -2266
rect 581866 -2502 582102 -2266
rect 581546 -2822 581782 -2586
rect 581866 -2822 582102 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 672938 588458 673174
rect 588542 672938 588778 673174
rect 588222 672618 588458 672854
rect 588542 672618 588778 672854
rect 588222 636938 588458 637174
rect 588542 636938 588778 637174
rect 588222 636618 588458 636854
rect 588542 636618 588778 636854
rect 588222 600938 588458 601174
rect 588542 600938 588778 601174
rect 588222 600618 588458 600854
rect 588542 600618 588778 600854
rect 588222 564938 588458 565174
rect 588542 564938 588778 565174
rect 588222 564618 588458 564854
rect 588542 564618 588778 564854
rect 588222 528938 588458 529174
rect 588542 528938 588778 529174
rect 588222 528618 588458 528854
rect 588542 528618 588778 528854
rect 588222 492938 588458 493174
rect 588542 492938 588778 493174
rect 588222 492618 588458 492854
rect 588542 492618 588778 492854
rect 588222 456938 588458 457174
rect 588542 456938 588778 457174
rect 588222 456618 588458 456854
rect 588542 456618 588778 456854
rect 588222 420938 588458 421174
rect 588542 420938 588778 421174
rect 588222 420618 588458 420854
rect 588542 420618 588778 420854
rect 588222 384938 588458 385174
rect 588542 384938 588778 385174
rect 588222 384618 588458 384854
rect 588542 384618 588778 384854
rect 588222 348938 588458 349174
rect 588542 348938 588778 349174
rect 588222 348618 588458 348854
rect 588542 348618 588778 348854
rect 588222 312938 588458 313174
rect 588542 312938 588778 313174
rect 588222 312618 588458 312854
rect 588542 312618 588778 312854
rect 588222 276938 588458 277174
rect 588542 276938 588778 277174
rect 588222 276618 588458 276854
rect 588542 276618 588778 276854
rect 588222 240938 588458 241174
rect 588542 240938 588778 241174
rect 588222 240618 588458 240854
rect 588542 240618 588778 240854
rect 588222 204938 588458 205174
rect 588542 204938 588778 205174
rect 588222 204618 588458 204854
rect 588542 204618 588778 204854
rect 588222 168938 588458 169174
rect 588542 168938 588778 169174
rect 588222 168618 588458 168854
rect 588542 168618 588778 168854
rect 588222 132938 588458 133174
rect 588542 132938 588778 133174
rect 588222 132618 588458 132854
rect 588542 132618 588778 132854
rect 588222 96938 588458 97174
rect 588542 96938 588778 97174
rect 588222 96618 588458 96854
rect 588542 96618 588778 96854
rect 588222 60938 588458 61174
rect 588542 60938 588778 61174
rect 588222 60618 588458 60854
rect 588542 60618 588778 60854
rect 588222 24938 588458 25174
rect 588542 24938 588778 25174
rect 588222 24618 588458 24854
rect 588542 24618 588778 24854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 694658 589418 694894
rect 589502 694658 589738 694894
rect 589182 694338 589418 694574
rect 589502 694338 589738 694574
rect 589182 658658 589418 658894
rect 589502 658658 589738 658894
rect 589182 658338 589418 658574
rect 589502 658338 589738 658574
rect 589182 622658 589418 622894
rect 589502 622658 589738 622894
rect 589182 622338 589418 622574
rect 589502 622338 589738 622574
rect 589182 586658 589418 586894
rect 589502 586658 589738 586894
rect 589182 586338 589418 586574
rect 589502 586338 589738 586574
rect 589182 550658 589418 550894
rect 589502 550658 589738 550894
rect 589182 550338 589418 550574
rect 589502 550338 589738 550574
rect 589182 514658 589418 514894
rect 589502 514658 589738 514894
rect 589182 514338 589418 514574
rect 589502 514338 589738 514574
rect 589182 478658 589418 478894
rect 589502 478658 589738 478894
rect 589182 478338 589418 478574
rect 589502 478338 589738 478574
rect 589182 442658 589418 442894
rect 589502 442658 589738 442894
rect 589182 442338 589418 442574
rect 589502 442338 589738 442574
rect 589182 406658 589418 406894
rect 589502 406658 589738 406894
rect 589182 406338 589418 406574
rect 589502 406338 589738 406574
rect 589182 370658 589418 370894
rect 589502 370658 589738 370894
rect 589182 370338 589418 370574
rect 589502 370338 589738 370574
rect 589182 334658 589418 334894
rect 589502 334658 589738 334894
rect 589182 334338 589418 334574
rect 589502 334338 589738 334574
rect 589182 298658 589418 298894
rect 589502 298658 589738 298894
rect 589182 298338 589418 298574
rect 589502 298338 589738 298574
rect 589182 262658 589418 262894
rect 589502 262658 589738 262894
rect 589182 262338 589418 262574
rect 589502 262338 589738 262574
rect 589182 226658 589418 226894
rect 589502 226658 589738 226894
rect 589182 226338 589418 226574
rect 589502 226338 589738 226574
rect 589182 190658 589418 190894
rect 589502 190658 589738 190894
rect 589182 190338 589418 190574
rect 589502 190338 589738 190574
rect 589182 154658 589418 154894
rect 589502 154658 589738 154894
rect 589182 154338 589418 154574
rect 589502 154338 589738 154574
rect 589182 118658 589418 118894
rect 589502 118658 589738 118894
rect 589182 118338 589418 118574
rect 589502 118338 589738 118574
rect 589182 82658 589418 82894
rect 589502 82658 589738 82894
rect 589182 82338 589418 82574
rect 589502 82338 589738 82574
rect 589182 46658 589418 46894
rect 589502 46658 589738 46894
rect 589182 46338 589418 46574
rect 589502 46338 589738 46574
rect 589182 10658 589418 10894
rect 589502 10658 589738 10894
rect 589182 10338 589418 10574
rect 589502 10338 589738 10574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 676658 590378 676894
rect 590462 676658 590698 676894
rect 590142 676338 590378 676574
rect 590462 676338 590698 676574
rect 590142 640658 590378 640894
rect 590462 640658 590698 640894
rect 590142 640338 590378 640574
rect 590462 640338 590698 640574
rect 590142 604658 590378 604894
rect 590462 604658 590698 604894
rect 590142 604338 590378 604574
rect 590462 604338 590698 604574
rect 590142 568658 590378 568894
rect 590462 568658 590698 568894
rect 590142 568338 590378 568574
rect 590462 568338 590698 568574
rect 590142 532658 590378 532894
rect 590462 532658 590698 532894
rect 590142 532338 590378 532574
rect 590462 532338 590698 532574
rect 590142 496658 590378 496894
rect 590462 496658 590698 496894
rect 590142 496338 590378 496574
rect 590462 496338 590698 496574
rect 590142 460658 590378 460894
rect 590462 460658 590698 460894
rect 590142 460338 590378 460574
rect 590462 460338 590698 460574
rect 590142 424658 590378 424894
rect 590462 424658 590698 424894
rect 590142 424338 590378 424574
rect 590462 424338 590698 424574
rect 590142 388658 590378 388894
rect 590462 388658 590698 388894
rect 590142 388338 590378 388574
rect 590462 388338 590698 388574
rect 590142 352658 590378 352894
rect 590462 352658 590698 352894
rect 590142 352338 590378 352574
rect 590462 352338 590698 352574
rect 590142 316658 590378 316894
rect 590462 316658 590698 316894
rect 590142 316338 590378 316574
rect 590462 316338 590698 316574
rect 590142 280658 590378 280894
rect 590462 280658 590698 280894
rect 590142 280338 590378 280574
rect 590462 280338 590698 280574
rect 590142 244658 590378 244894
rect 590462 244658 590698 244894
rect 590142 244338 590378 244574
rect 590462 244338 590698 244574
rect 590142 208658 590378 208894
rect 590462 208658 590698 208894
rect 590142 208338 590378 208574
rect 590462 208338 590698 208574
rect 590142 172658 590378 172894
rect 590462 172658 590698 172894
rect 590142 172338 590378 172574
rect 590462 172338 590698 172574
rect 590142 136658 590378 136894
rect 590462 136658 590698 136894
rect 590142 136338 590378 136574
rect 590462 136338 590698 136574
rect 590142 100658 590378 100894
rect 590462 100658 590698 100894
rect 590142 100338 590378 100574
rect 590462 100338 590698 100574
rect 590142 64658 590378 64894
rect 590462 64658 590698 64894
rect 590142 64338 590378 64574
rect 590462 64338 590698 64574
rect 590142 28658 590378 28894
rect 590462 28658 590698 28894
rect 590142 28338 590378 28574
rect 590462 28338 590698 28574
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 698378 591338 698614
rect 591422 698378 591658 698614
rect 591102 698058 591338 698294
rect 591422 698058 591658 698294
rect 591102 662378 591338 662614
rect 591422 662378 591658 662614
rect 591102 662058 591338 662294
rect 591422 662058 591658 662294
rect 591102 626378 591338 626614
rect 591422 626378 591658 626614
rect 591102 626058 591338 626294
rect 591422 626058 591658 626294
rect 591102 590378 591338 590614
rect 591422 590378 591658 590614
rect 591102 590058 591338 590294
rect 591422 590058 591658 590294
rect 591102 554378 591338 554614
rect 591422 554378 591658 554614
rect 591102 554058 591338 554294
rect 591422 554058 591658 554294
rect 591102 518378 591338 518614
rect 591422 518378 591658 518614
rect 591102 518058 591338 518294
rect 591422 518058 591658 518294
rect 591102 482378 591338 482614
rect 591422 482378 591658 482614
rect 591102 482058 591338 482294
rect 591422 482058 591658 482294
rect 591102 446378 591338 446614
rect 591422 446378 591658 446614
rect 591102 446058 591338 446294
rect 591422 446058 591658 446294
rect 591102 410378 591338 410614
rect 591422 410378 591658 410614
rect 591102 410058 591338 410294
rect 591422 410058 591658 410294
rect 591102 374378 591338 374614
rect 591422 374378 591658 374614
rect 591102 374058 591338 374294
rect 591422 374058 591658 374294
rect 591102 338378 591338 338614
rect 591422 338378 591658 338614
rect 591102 338058 591338 338294
rect 591422 338058 591658 338294
rect 591102 302378 591338 302614
rect 591422 302378 591658 302614
rect 591102 302058 591338 302294
rect 591422 302058 591658 302294
rect 591102 266378 591338 266614
rect 591422 266378 591658 266614
rect 591102 266058 591338 266294
rect 591422 266058 591658 266294
rect 591102 230378 591338 230614
rect 591422 230378 591658 230614
rect 591102 230058 591338 230294
rect 591422 230058 591658 230294
rect 591102 194378 591338 194614
rect 591422 194378 591658 194614
rect 591102 194058 591338 194294
rect 591422 194058 591658 194294
rect 591102 158378 591338 158614
rect 591422 158378 591658 158614
rect 591102 158058 591338 158294
rect 591422 158058 591658 158294
rect 591102 122378 591338 122614
rect 591422 122378 591658 122614
rect 591102 122058 591338 122294
rect 591422 122058 591658 122294
rect 591102 86378 591338 86614
rect 591422 86378 591658 86614
rect 591102 86058 591338 86294
rect 591422 86058 591658 86294
rect 591102 50378 591338 50614
rect 591422 50378 591658 50614
rect 591102 50058 591338 50294
rect 591422 50058 591658 50294
rect 591102 14378 591338 14614
rect 591422 14378 591658 14614
rect 591102 14058 591338 14294
rect 591422 14058 591658 14294
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 680378 592298 680614
rect 592382 680378 592618 680614
rect 592062 680058 592298 680294
rect 592382 680058 592618 680294
rect 592062 644378 592298 644614
rect 592382 644378 592618 644614
rect 592062 644058 592298 644294
rect 592382 644058 592618 644294
rect 592062 608378 592298 608614
rect 592382 608378 592618 608614
rect 592062 608058 592298 608294
rect 592382 608058 592618 608294
rect 592062 572378 592298 572614
rect 592382 572378 592618 572614
rect 592062 572058 592298 572294
rect 592382 572058 592618 572294
rect 592062 536378 592298 536614
rect 592382 536378 592618 536614
rect 592062 536058 592298 536294
rect 592382 536058 592618 536294
rect 592062 500378 592298 500614
rect 592382 500378 592618 500614
rect 592062 500058 592298 500294
rect 592382 500058 592618 500294
rect 592062 464378 592298 464614
rect 592382 464378 592618 464614
rect 592062 464058 592298 464294
rect 592382 464058 592618 464294
rect 592062 428378 592298 428614
rect 592382 428378 592618 428614
rect 592062 428058 592298 428294
rect 592382 428058 592618 428294
rect 592062 392378 592298 392614
rect 592382 392378 592618 392614
rect 592062 392058 592298 392294
rect 592382 392058 592618 392294
rect 592062 356378 592298 356614
rect 592382 356378 592618 356614
rect 592062 356058 592298 356294
rect 592382 356058 592618 356294
rect 592062 320378 592298 320614
rect 592382 320378 592618 320614
rect 592062 320058 592298 320294
rect 592382 320058 592618 320294
rect 592062 284378 592298 284614
rect 592382 284378 592618 284614
rect 592062 284058 592298 284294
rect 592382 284058 592618 284294
rect 592062 248378 592298 248614
rect 592382 248378 592618 248614
rect 592062 248058 592298 248294
rect 592382 248058 592618 248294
rect 592062 212378 592298 212614
rect 592382 212378 592618 212614
rect 592062 212058 592298 212294
rect 592382 212058 592618 212294
rect 592062 176378 592298 176614
rect 592382 176378 592618 176614
rect 592062 176058 592298 176294
rect 592382 176058 592618 176294
rect 592062 140378 592298 140614
rect 592382 140378 592618 140614
rect 592062 140058 592298 140294
rect 592382 140058 592618 140294
rect 592062 104378 592298 104614
rect 592382 104378 592618 104614
rect 592062 104058 592298 104294
rect 592382 104058 592618 104294
rect 592062 68378 592298 68614
rect 592382 68378 592618 68614
rect 592062 68058 592298 68294
rect 592382 68058 592618 68294
rect 592062 32378 592298 32614
rect 592382 32378 592618 32614
rect 592062 32058 592298 32294
rect 592382 32058 592618 32294
rect 570986 -7302 571222 -7066
rect 571306 -7302 571542 -7066
rect 570986 -7622 571222 -7386
rect 571306 -7622 571542 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 592650 698294
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 590730 694894
rect -6806 694574 590730 694658
rect -6806 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 590730 694574
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 588810 691174
rect -4886 690854 588810 690938
rect -4886 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 588810 690854
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 8250 687454
rect 8486 687218 38970 687454
rect 39206 687218 69690 687454
rect 69926 687218 100410 687454
rect 100646 687218 131130 687454
rect 131366 687218 161850 687454
rect 162086 687218 192570 687454
rect 192806 687218 223290 687454
rect 223526 687218 254010 687454
rect 254246 687218 284730 687454
rect 284966 687218 315450 687454
rect 315686 687218 346170 687454
rect 346406 687218 376890 687454
rect 377126 687218 407610 687454
rect 407846 687218 438330 687454
rect 438566 687218 469050 687454
rect 469286 687218 499770 687454
rect 500006 687218 530490 687454
rect 530726 687218 561210 687454
rect 561446 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 8250 687134
rect 8486 686898 38970 687134
rect 39206 686898 69690 687134
rect 69926 686898 100410 687134
rect 100646 686898 131130 687134
rect 131366 686898 161850 687134
rect 162086 686898 192570 687134
rect 192806 686898 223290 687134
rect 223526 686898 254010 687134
rect 254246 686898 284730 687134
rect 284966 686898 315450 687134
rect 315686 686898 346170 687134
rect 346406 686898 376890 687134
rect 377126 686898 407610 687134
rect 407846 686898 438330 687134
rect 438566 686898 469050 687134
rect 469286 686898 499770 687134
rect 500006 686898 530490 687134
rect 530726 686898 561210 687134
rect 561446 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect -8726 680294 592650 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect -6806 676574 590730 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect -4886 672854 588810 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 23610 669454
rect 23846 669218 54330 669454
rect 54566 669218 85050 669454
rect 85286 669218 115770 669454
rect 116006 669218 146490 669454
rect 146726 669218 177210 669454
rect 177446 669218 207930 669454
rect 208166 669218 238650 669454
rect 238886 669218 269370 669454
rect 269606 669218 300090 669454
rect 300326 669218 330810 669454
rect 331046 669218 361530 669454
rect 361766 669218 392250 669454
rect 392486 669218 422970 669454
rect 423206 669218 453690 669454
rect 453926 669218 484410 669454
rect 484646 669218 515130 669454
rect 515366 669218 545850 669454
rect 546086 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 23610 669134
rect 23846 668898 54330 669134
rect 54566 668898 85050 669134
rect 85286 668898 115770 669134
rect 116006 668898 146490 669134
rect 146726 668898 177210 669134
rect 177446 668898 207930 669134
rect 208166 668898 238650 669134
rect 238886 668898 269370 669134
rect 269606 668898 300090 669134
rect 300326 668898 330810 669134
rect 331046 668898 361530 669134
rect 361766 668898 392250 669134
rect 392486 668898 422970 669134
rect 423206 668898 453690 669134
rect 453926 668898 484410 669134
rect 484646 668898 515130 669134
rect 515366 668898 545850 669134
rect 546086 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 592650 662294
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 590730 658894
rect -6806 658574 590730 658658
rect -6806 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 590730 658574
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 588810 655174
rect -4886 654854 588810 654938
rect -4886 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 588810 654854
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 8250 651454
rect 8486 651218 38970 651454
rect 39206 651218 69690 651454
rect 69926 651218 100410 651454
rect 100646 651218 131130 651454
rect 131366 651218 161850 651454
rect 162086 651218 192570 651454
rect 192806 651218 223290 651454
rect 223526 651218 254010 651454
rect 254246 651218 284730 651454
rect 284966 651218 315450 651454
rect 315686 651218 346170 651454
rect 346406 651218 376890 651454
rect 377126 651218 407610 651454
rect 407846 651218 438330 651454
rect 438566 651218 469050 651454
rect 469286 651218 499770 651454
rect 500006 651218 530490 651454
rect 530726 651218 561210 651454
rect 561446 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 8250 651134
rect 8486 650898 38970 651134
rect 39206 650898 69690 651134
rect 69926 650898 100410 651134
rect 100646 650898 131130 651134
rect 131366 650898 161850 651134
rect 162086 650898 192570 651134
rect 192806 650898 223290 651134
rect 223526 650898 254010 651134
rect 254246 650898 284730 651134
rect 284966 650898 315450 651134
rect 315686 650898 346170 651134
rect 346406 650898 376890 651134
rect 377126 650898 407610 651134
rect 407846 650898 438330 651134
rect 438566 650898 469050 651134
rect 469286 650898 499770 651134
rect 500006 650898 530490 651134
rect 530726 650898 561210 651134
rect 561446 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect -8726 644294 592650 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect -6806 640574 590730 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect -4886 636854 588810 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 23610 633454
rect 23846 633218 54330 633454
rect 54566 633218 85050 633454
rect 85286 633218 115770 633454
rect 116006 633218 146490 633454
rect 146726 633218 177210 633454
rect 177446 633218 207930 633454
rect 208166 633218 238650 633454
rect 238886 633218 269370 633454
rect 269606 633218 300090 633454
rect 300326 633218 330810 633454
rect 331046 633218 361530 633454
rect 361766 633218 392250 633454
rect 392486 633218 422970 633454
rect 423206 633218 453690 633454
rect 453926 633218 484410 633454
rect 484646 633218 515130 633454
rect 515366 633218 545850 633454
rect 546086 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 23610 633134
rect 23846 632898 54330 633134
rect 54566 632898 85050 633134
rect 85286 632898 115770 633134
rect 116006 632898 146490 633134
rect 146726 632898 177210 633134
rect 177446 632898 207930 633134
rect 208166 632898 238650 633134
rect 238886 632898 269370 633134
rect 269606 632898 300090 633134
rect 300326 632898 330810 633134
rect 331046 632898 361530 633134
rect 361766 632898 392250 633134
rect 392486 632898 422970 633134
rect 423206 632898 453690 633134
rect 453926 632898 484410 633134
rect 484646 632898 515130 633134
rect 515366 632898 545850 633134
rect 546086 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 592650 626294
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 590730 622894
rect -6806 622574 590730 622658
rect -6806 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 590730 622574
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 588810 619174
rect -4886 618854 588810 618938
rect -4886 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 588810 618854
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 8250 615454
rect 8486 615218 38970 615454
rect 39206 615218 69690 615454
rect 69926 615218 100410 615454
rect 100646 615218 131130 615454
rect 131366 615218 161850 615454
rect 162086 615218 192570 615454
rect 192806 615218 223290 615454
rect 223526 615218 254010 615454
rect 254246 615218 284730 615454
rect 284966 615218 315450 615454
rect 315686 615218 346170 615454
rect 346406 615218 376890 615454
rect 377126 615218 407610 615454
rect 407846 615218 438330 615454
rect 438566 615218 469050 615454
rect 469286 615218 499770 615454
rect 500006 615218 530490 615454
rect 530726 615218 561210 615454
rect 561446 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 8250 615134
rect 8486 614898 38970 615134
rect 39206 614898 69690 615134
rect 69926 614898 100410 615134
rect 100646 614898 131130 615134
rect 131366 614898 161850 615134
rect 162086 614898 192570 615134
rect 192806 614898 223290 615134
rect 223526 614898 254010 615134
rect 254246 614898 284730 615134
rect 284966 614898 315450 615134
rect 315686 614898 346170 615134
rect 346406 614898 376890 615134
rect 377126 614898 407610 615134
rect 407846 614898 438330 615134
rect 438566 614898 469050 615134
rect 469286 614898 499770 615134
rect 500006 614898 530490 615134
rect 530726 614898 561210 615134
rect 561446 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect -8726 608294 592650 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect -6806 604574 590730 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect -4886 600854 588810 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 23610 597454
rect 23846 597218 54330 597454
rect 54566 597218 85050 597454
rect 85286 597218 115770 597454
rect 116006 597218 146490 597454
rect 146726 597218 177210 597454
rect 177446 597218 207930 597454
rect 208166 597218 238650 597454
rect 238886 597218 269370 597454
rect 269606 597218 300090 597454
rect 300326 597218 330810 597454
rect 331046 597218 361530 597454
rect 361766 597218 392250 597454
rect 392486 597218 422970 597454
rect 423206 597218 453690 597454
rect 453926 597218 484410 597454
rect 484646 597218 515130 597454
rect 515366 597218 545850 597454
rect 546086 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 23610 597134
rect 23846 596898 54330 597134
rect 54566 596898 85050 597134
rect 85286 596898 115770 597134
rect 116006 596898 146490 597134
rect 146726 596898 177210 597134
rect 177446 596898 207930 597134
rect 208166 596898 238650 597134
rect 238886 596898 269370 597134
rect 269606 596898 300090 597134
rect 300326 596898 330810 597134
rect 331046 596898 361530 597134
rect 361766 596898 392250 597134
rect 392486 596898 422970 597134
rect 423206 596898 453690 597134
rect 453926 596898 484410 597134
rect 484646 596898 515130 597134
rect 515366 596898 545850 597134
rect 546086 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 592650 590294
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 590730 586894
rect -6806 586574 590730 586658
rect -6806 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 590730 586574
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 588810 583174
rect -4886 582854 588810 582938
rect -4886 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 588810 582854
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 8250 579454
rect 8486 579218 38970 579454
rect 39206 579218 69690 579454
rect 69926 579218 100410 579454
rect 100646 579218 131130 579454
rect 131366 579218 161850 579454
rect 162086 579218 192570 579454
rect 192806 579218 223290 579454
rect 223526 579218 254010 579454
rect 254246 579218 284730 579454
rect 284966 579218 315450 579454
rect 315686 579218 346170 579454
rect 346406 579218 376890 579454
rect 377126 579218 407610 579454
rect 407846 579218 438330 579454
rect 438566 579218 469050 579454
rect 469286 579218 499770 579454
rect 500006 579218 530490 579454
rect 530726 579218 561210 579454
rect 561446 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 8250 579134
rect 8486 578898 38970 579134
rect 39206 578898 69690 579134
rect 69926 578898 100410 579134
rect 100646 578898 131130 579134
rect 131366 578898 161850 579134
rect 162086 578898 192570 579134
rect 192806 578898 223290 579134
rect 223526 578898 254010 579134
rect 254246 578898 284730 579134
rect 284966 578898 315450 579134
rect 315686 578898 346170 579134
rect 346406 578898 376890 579134
rect 377126 578898 407610 579134
rect 407846 578898 438330 579134
rect 438566 578898 469050 579134
rect 469286 578898 499770 579134
rect 500006 578898 530490 579134
rect 530726 578898 561210 579134
rect 561446 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect -8726 572294 592650 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect -6806 568574 590730 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect -4886 564854 588810 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect -4886 564586 588810 564618
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 23610 561454
rect 23846 561218 54330 561454
rect 54566 561218 85050 561454
rect 85286 561218 115770 561454
rect 116006 561218 146490 561454
rect 146726 561218 177210 561454
rect 177446 561218 207930 561454
rect 208166 561218 238650 561454
rect 238886 561218 269370 561454
rect 269606 561218 300090 561454
rect 300326 561218 330810 561454
rect 331046 561218 361530 561454
rect 361766 561218 392250 561454
rect 392486 561218 422970 561454
rect 423206 561218 453690 561454
rect 453926 561218 484410 561454
rect 484646 561218 515130 561454
rect 515366 561218 545850 561454
rect 546086 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 23610 561134
rect 23846 560898 54330 561134
rect 54566 560898 85050 561134
rect 85286 560898 115770 561134
rect 116006 560898 146490 561134
rect 146726 560898 177210 561134
rect 177446 560898 207930 561134
rect 208166 560898 238650 561134
rect 238886 560898 269370 561134
rect 269606 560898 300090 561134
rect 300326 560898 330810 561134
rect 331046 560898 361530 561134
rect 361766 560898 392250 561134
rect 392486 560898 422970 561134
rect 423206 560898 453690 561134
rect 453926 560898 484410 561134
rect 484646 560898 515130 561134
rect 515366 560898 545850 561134
rect 546086 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 592650 554294
rect -8726 554026 592650 554058
rect -6806 550894 590730 550926
rect -6806 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 590730 550894
rect -6806 550574 590730 550658
rect -6806 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 590730 550574
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 588810 547174
rect -4886 546854 588810 546938
rect -4886 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 588810 546854
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 8250 543454
rect 8486 543218 38970 543454
rect 39206 543218 69690 543454
rect 69926 543218 100410 543454
rect 100646 543218 131130 543454
rect 131366 543218 161850 543454
rect 162086 543218 192570 543454
rect 192806 543218 223290 543454
rect 223526 543218 254010 543454
rect 254246 543218 284730 543454
rect 284966 543218 315450 543454
rect 315686 543218 346170 543454
rect 346406 543218 376890 543454
rect 377126 543218 407610 543454
rect 407846 543218 438330 543454
rect 438566 543218 469050 543454
rect 469286 543218 499770 543454
rect 500006 543218 530490 543454
rect 530726 543218 561210 543454
rect 561446 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 8250 543134
rect 8486 542898 38970 543134
rect 39206 542898 69690 543134
rect 69926 542898 100410 543134
rect 100646 542898 131130 543134
rect 131366 542898 161850 543134
rect 162086 542898 192570 543134
rect 192806 542898 223290 543134
rect 223526 542898 254010 543134
rect 254246 542898 284730 543134
rect 284966 542898 315450 543134
rect 315686 542898 346170 543134
rect 346406 542898 376890 543134
rect 377126 542898 407610 543134
rect 407846 542898 438330 543134
rect 438566 542898 469050 543134
rect 469286 542898 499770 543134
rect 500006 542898 530490 543134
rect 530726 542898 561210 543134
rect 561446 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect -8726 536294 592650 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect -6806 532574 590730 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect -4886 528854 588810 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 23610 525454
rect 23846 525218 54330 525454
rect 54566 525218 85050 525454
rect 85286 525218 115770 525454
rect 116006 525218 146490 525454
rect 146726 525218 177210 525454
rect 177446 525218 207930 525454
rect 208166 525218 238650 525454
rect 238886 525218 269370 525454
rect 269606 525218 300090 525454
rect 300326 525218 330810 525454
rect 331046 525218 361530 525454
rect 361766 525218 392250 525454
rect 392486 525218 422970 525454
rect 423206 525218 453690 525454
rect 453926 525218 484410 525454
rect 484646 525218 515130 525454
rect 515366 525218 545850 525454
rect 546086 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 23610 525134
rect 23846 524898 54330 525134
rect 54566 524898 85050 525134
rect 85286 524898 115770 525134
rect 116006 524898 146490 525134
rect 146726 524898 177210 525134
rect 177446 524898 207930 525134
rect 208166 524898 238650 525134
rect 238886 524898 269370 525134
rect 269606 524898 300090 525134
rect 300326 524898 330810 525134
rect 331046 524898 361530 525134
rect 361766 524898 392250 525134
rect 392486 524898 422970 525134
rect 423206 524898 453690 525134
rect 453926 524898 484410 525134
rect 484646 524898 515130 525134
rect 515366 524898 545850 525134
rect 546086 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 592650 518294
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 590730 514894
rect -6806 514574 590730 514658
rect -6806 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 590730 514574
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 588810 511174
rect -4886 510854 588810 510938
rect -4886 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 588810 510854
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 8250 507454
rect 8486 507218 38970 507454
rect 39206 507218 69690 507454
rect 69926 507218 100410 507454
rect 100646 507218 131130 507454
rect 131366 507218 161850 507454
rect 162086 507218 192570 507454
rect 192806 507218 223290 507454
rect 223526 507218 254010 507454
rect 254246 507218 284730 507454
rect 284966 507218 315450 507454
rect 315686 507218 346170 507454
rect 346406 507218 376890 507454
rect 377126 507218 407610 507454
rect 407846 507218 438330 507454
rect 438566 507218 469050 507454
rect 469286 507218 499770 507454
rect 500006 507218 530490 507454
rect 530726 507218 561210 507454
rect 561446 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 8250 507134
rect 8486 506898 38970 507134
rect 39206 506898 69690 507134
rect 69926 506898 100410 507134
rect 100646 506898 131130 507134
rect 131366 506898 161850 507134
rect 162086 506898 192570 507134
rect 192806 506898 223290 507134
rect 223526 506898 254010 507134
rect 254246 506898 284730 507134
rect 284966 506898 315450 507134
rect 315686 506898 346170 507134
rect 346406 506898 376890 507134
rect 377126 506898 407610 507134
rect 407846 506898 438330 507134
rect 438566 506898 469050 507134
rect 469286 506898 499770 507134
rect 500006 506898 530490 507134
rect 530726 506898 561210 507134
rect 561446 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect -8726 500294 592650 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect -6806 496574 590730 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect -4886 492854 588810 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 23610 489454
rect 23846 489218 54330 489454
rect 54566 489218 85050 489454
rect 85286 489218 115770 489454
rect 116006 489218 146490 489454
rect 146726 489218 177210 489454
rect 177446 489218 207930 489454
rect 208166 489218 238650 489454
rect 238886 489218 269370 489454
rect 269606 489218 300090 489454
rect 300326 489218 330810 489454
rect 331046 489218 361530 489454
rect 361766 489218 392250 489454
rect 392486 489218 422970 489454
rect 423206 489218 453690 489454
rect 453926 489218 484410 489454
rect 484646 489218 515130 489454
rect 515366 489218 545850 489454
rect 546086 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 23610 489134
rect 23846 488898 54330 489134
rect 54566 488898 85050 489134
rect 85286 488898 115770 489134
rect 116006 488898 146490 489134
rect 146726 488898 177210 489134
rect 177446 488898 207930 489134
rect 208166 488898 238650 489134
rect 238886 488898 269370 489134
rect 269606 488898 300090 489134
rect 300326 488898 330810 489134
rect 331046 488898 361530 489134
rect 361766 488898 392250 489134
rect 392486 488898 422970 489134
rect 423206 488898 453690 489134
rect 453926 488898 484410 489134
rect 484646 488898 515130 489134
rect 515366 488898 545850 489134
rect 546086 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 592650 482294
rect -8726 482026 592650 482058
rect -6806 478894 590730 478926
rect -6806 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 590730 478894
rect -6806 478574 590730 478658
rect -6806 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 590730 478574
rect -6806 478306 590730 478338
rect -4886 475174 588810 475206
rect -4886 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 588810 475174
rect -4886 474854 588810 474938
rect -4886 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 588810 474854
rect -4886 474586 588810 474618
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 8250 471454
rect 8486 471218 38970 471454
rect 39206 471218 69690 471454
rect 69926 471218 100410 471454
rect 100646 471218 131130 471454
rect 131366 471218 161850 471454
rect 162086 471218 192570 471454
rect 192806 471218 223290 471454
rect 223526 471218 254010 471454
rect 254246 471218 284730 471454
rect 284966 471218 315450 471454
rect 315686 471218 346170 471454
rect 346406 471218 376890 471454
rect 377126 471218 407610 471454
rect 407846 471218 438330 471454
rect 438566 471218 469050 471454
rect 469286 471218 499770 471454
rect 500006 471218 530490 471454
rect 530726 471218 561210 471454
rect 561446 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 8250 471134
rect 8486 470898 38970 471134
rect 39206 470898 69690 471134
rect 69926 470898 100410 471134
rect 100646 470898 131130 471134
rect 131366 470898 161850 471134
rect 162086 470898 192570 471134
rect 192806 470898 223290 471134
rect 223526 470898 254010 471134
rect 254246 470898 284730 471134
rect 284966 470898 315450 471134
rect 315686 470898 346170 471134
rect 346406 470898 376890 471134
rect 377126 470898 407610 471134
rect 407846 470898 438330 471134
rect 438566 470898 469050 471134
rect 469286 470898 499770 471134
rect 500006 470898 530490 471134
rect 530726 470898 561210 471134
rect 561446 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect -8726 464294 592650 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect -6806 460574 590730 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect -4886 456854 588810 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 23610 453454
rect 23846 453218 54330 453454
rect 54566 453218 85050 453454
rect 85286 453218 115770 453454
rect 116006 453218 146490 453454
rect 146726 453218 177210 453454
rect 177446 453218 207930 453454
rect 208166 453218 238650 453454
rect 238886 453218 269370 453454
rect 269606 453218 300090 453454
rect 300326 453218 330810 453454
rect 331046 453218 361530 453454
rect 361766 453218 392250 453454
rect 392486 453218 422970 453454
rect 423206 453218 453690 453454
rect 453926 453218 484410 453454
rect 484646 453218 515130 453454
rect 515366 453218 545850 453454
rect 546086 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 23610 453134
rect 23846 452898 54330 453134
rect 54566 452898 85050 453134
rect 85286 452898 115770 453134
rect 116006 452898 146490 453134
rect 146726 452898 177210 453134
rect 177446 452898 207930 453134
rect 208166 452898 238650 453134
rect 238886 452898 269370 453134
rect 269606 452898 300090 453134
rect 300326 452898 330810 453134
rect 331046 452898 361530 453134
rect 361766 452898 392250 453134
rect 392486 452898 422970 453134
rect 423206 452898 453690 453134
rect 453926 452898 484410 453134
rect 484646 452898 515130 453134
rect 515366 452898 545850 453134
rect 546086 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 592650 446294
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 590730 442894
rect -6806 442574 590730 442658
rect -6806 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 590730 442574
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 588810 439174
rect -4886 438854 588810 438938
rect -4886 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 588810 438854
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 8250 435454
rect 8486 435218 38970 435454
rect 39206 435218 69690 435454
rect 69926 435218 100410 435454
rect 100646 435218 131130 435454
rect 131366 435218 161850 435454
rect 162086 435218 192570 435454
rect 192806 435218 223290 435454
rect 223526 435218 254010 435454
rect 254246 435218 284730 435454
rect 284966 435218 315450 435454
rect 315686 435218 346170 435454
rect 346406 435218 376890 435454
rect 377126 435218 407610 435454
rect 407846 435218 438330 435454
rect 438566 435218 469050 435454
rect 469286 435218 499770 435454
rect 500006 435218 530490 435454
rect 530726 435218 561210 435454
rect 561446 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 8250 435134
rect 8486 434898 38970 435134
rect 39206 434898 69690 435134
rect 69926 434898 100410 435134
rect 100646 434898 131130 435134
rect 131366 434898 161850 435134
rect 162086 434898 192570 435134
rect 192806 434898 223290 435134
rect 223526 434898 254010 435134
rect 254246 434898 284730 435134
rect 284966 434898 315450 435134
rect 315686 434898 346170 435134
rect 346406 434898 376890 435134
rect 377126 434898 407610 435134
rect 407846 434898 438330 435134
rect 438566 434898 469050 435134
rect 469286 434898 499770 435134
rect 500006 434898 530490 435134
rect 530726 434898 561210 435134
rect 561446 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect -8726 428294 592650 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect -6806 424574 590730 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect -4886 420854 588810 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 23610 417454
rect 23846 417218 54330 417454
rect 54566 417218 85050 417454
rect 85286 417218 115770 417454
rect 116006 417218 146490 417454
rect 146726 417218 177210 417454
rect 177446 417218 207930 417454
rect 208166 417218 238650 417454
rect 238886 417218 269370 417454
rect 269606 417218 300090 417454
rect 300326 417218 330810 417454
rect 331046 417218 361530 417454
rect 361766 417218 392250 417454
rect 392486 417218 422970 417454
rect 423206 417218 453690 417454
rect 453926 417218 484410 417454
rect 484646 417218 515130 417454
rect 515366 417218 545850 417454
rect 546086 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 23610 417134
rect 23846 416898 54330 417134
rect 54566 416898 85050 417134
rect 85286 416898 115770 417134
rect 116006 416898 146490 417134
rect 146726 416898 177210 417134
rect 177446 416898 207930 417134
rect 208166 416898 238650 417134
rect 238886 416898 269370 417134
rect 269606 416898 300090 417134
rect 300326 416898 330810 417134
rect 331046 416898 361530 417134
rect 361766 416898 392250 417134
rect 392486 416898 422970 417134
rect 423206 416898 453690 417134
rect 453926 416898 484410 417134
rect 484646 416898 515130 417134
rect 515366 416898 545850 417134
rect 546086 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 592650 410294
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 590730 406894
rect -6806 406574 590730 406658
rect -6806 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 590730 406574
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 588810 403174
rect -4886 402854 588810 402938
rect -4886 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 588810 402854
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 8250 399454
rect 8486 399218 38970 399454
rect 39206 399218 69690 399454
rect 69926 399218 100410 399454
rect 100646 399218 131130 399454
rect 131366 399218 161850 399454
rect 162086 399218 192570 399454
rect 192806 399218 223290 399454
rect 223526 399218 254010 399454
rect 254246 399218 284730 399454
rect 284966 399218 315450 399454
rect 315686 399218 346170 399454
rect 346406 399218 376890 399454
rect 377126 399218 407610 399454
rect 407846 399218 438330 399454
rect 438566 399218 469050 399454
rect 469286 399218 499770 399454
rect 500006 399218 530490 399454
rect 530726 399218 561210 399454
rect 561446 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 8250 399134
rect 8486 398898 38970 399134
rect 39206 398898 69690 399134
rect 69926 398898 100410 399134
rect 100646 398898 131130 399134
rect 131366 398898 161850 399134
rect 162086 398898 192570 399134
rect 192806 398898 223290 399134
rect 223526 398898 254010 399134
rect 254246 398898 284730 399134
rect 284966 398898 315450 399134
rect 315686 398898 346170 399134
rect 346406 398898 376890 399134
rect 377126 398898 407610 399134
rect 407846 398898 438330 399134
rect 438566 398898 469050 399134
rect 469286 398898 499770 399134
rect 500006 398898 530490 399134
rect 530726 398898 561210 399134
rect 561446 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect -8726 392294 592650 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect -8726 392026 592650 392058
rect -6806 388894 590730 388926
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect -6806 388574 590730 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect -4886 384854 588810 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 23610 381454
rect 23846 381218 54330 381454
rect 54566 381218 85050 381454
rect 85286 381218 115770 381454
rect 116006 381218 146490 381454
rect 146726 381218 177210 381454
rect 177446 381218 207930 381454
rect 208166 381218 238650 381454
rect 238886 381218 269370 381454
rect 269606 381218 300090 381454
rect 300326 381218 330810 381454
rect 331046 381218 361530 381454
rect 361766 381218 392250 381454
rect 392486 381218 422970 381454
rect 423206 381218 453690 381454
rect 453926 381218 484410 381454
rect 484646 381218 515130 381454
rect 515366 381218 545850 381454
rect 546086 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect -2966 381134 586890 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 23610 381134
rect 23846 380898 54330 381134
rect 54566 380898 85050 381134
rect 85286 380898 115770 381134
rect 116006 380898 146490 381134
rect 146726 380898 177210 381134
rect 177446 380898 207930 381134
rect 208166 380898 238650 381134
rect 238886 380898 269370 381134
rect 269606 380898 300090 381134
rect 300326 380898 330810 381134
rect 331046 380898 361530 381134
rect 361766 380898 392250 381134
rect 392486 380898 422970 381134
rect 423206 380898 453690 381134
rect 453926 380898 484410 381134
rect 484646 380898 515130 381134
rect 515366 380898 545850 381134
rect 546086 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 592650 374294
rect -8726 374026 592650 374058
rect -6806 370894 590730 370926
rect -6806 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 590730 370894
rect -6806 370574 590730 370658
rect -6806 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 590730 370574
rect -6806 370306 590730 370338
rect -4886 367174 588810 367206
rect -4886 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 588810 367174
rect -4886 366854 588810 366938
rect -4886 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 588810 366854
rect -4886 366586 588810 366618
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 8250 363454
rect 8486 363218 38970 363454
rect 39206 363218 69690 363454
rect 69926 363218 100410 363454
rect 100646 363218 131130 363454
rect 131366 363218 161850 363454
rect 162086 363218 192570 363454
rect 192806 363218 223290 363454
rect 223526 363218 254010 363454
rect 254246 363218 284730 363454
rect 284966 363218 315450 363454
rect 315686 363218 346170 363454
rect 346406 363218 376890 363454
rect 377126 363218 407610 363454
rect 407846 363218 438330 363454
rect 438566 363218 469050 363454
rect 469286 363218 499770 363454
rect 500006 363218 530490 363454
rect 530726 363218 561210 363454
rect 561446 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 8250 363134
rect 8486 362898 38970 363134
rect 39206 362898 69690 363134
rect 69926 362898 100410 363134
rect 100646 362898 131130 363134
rect 131366 362898 161850 363134
rect 162086 362898 192570 363134
rect 192806 362898 223290 363134
rect 223526 362898 254010 363134
rect 254246 362898 284730 363134
rect 284966 362898 315450 363134
rect 315686 362898 346170 363134
rect 346406 362898 376890 363134
rect 377126 362898 407610 363134
rect 407846 362898 438330 363134
rect 438566 362898 469050 363134
rect 469286 362898 499770 363134
rect 500006 362898 530490 363134
rect 530726 362898 561210 363134
rect 561446 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect -8726 356614 592650 356646
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect -8726 356294 592650 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect -6806 352574 590730 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect -4886 348854 588810 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect -4886 348586 588810 348618
rect -2966 345454 586890 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 23610 345454
rect 23846 345218 54330 345454
rect 54566 345218 85050 345454
rect 85286 345218 115770 345454
rect 116006 345218 146490 345454
rect 146726 345218 177210 345454
rect 177446 345218 207930 345454
rect 208166 345218 238650 345454
rect 238886 345218 269370 345454
rect 269606 345218 300090 345454
rect 300326 345218 330810 345454
rect 331046 345218 361530 345454
rect 361766 345218 392250 345454
rect 392486 345218 422970 345454
rect 423206 345218 453690 345454
rect 453926 345218 484410 345454
rect 484646 345218 515130 345454
rect 515366 345218 545850 345454
rect 546086 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect -2966 345134 586890 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 23610 345134
rect 23846 344898 54330 345134
rect 54566 344898 85050 345134
rect 85286 344898 115770 345134
rect 116006 344898 146490 345134
rect 146726 344898 177210 345134
rect 177446 344898 207930 345134
rect 208166 344898 238650 345134
rect 238886 344898 269370 345134
rect 269606 344898 300090 345134
rect 300326 344898 330810 345134
rect 331046 344898 361530 345134
rect 361766 344898 392250 345134
rect 392486 344898 422970 345134
rect 423206 344898 453690 345134
rect 453926 344898 484410 345134
rect 484646 344898 515130 345134
rect 515366 344898 545850 345134
rect 546086 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect -2966 344866 586890 344898
rect -8726 338614 592650 338646
rect -8726 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 592650 338294
rect -8726 338026 592650 338058
rect -6806 334894 590730 334926
rect -6806 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 590730 334894
rect -6806 334574 590730 334658
rect -6806 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 590730 334574
rect -6806 334306 590730 334338
rect -4886 331174 588810 331206
rect -4886 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 588810 331174
rect -4886 330854 588810 330938
rect -4886 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 588810 330854
rect -4886 330586 588810 330618
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 8250 327454
rect 8486 327218 38970 327454
rect 39206 327218 69690 327454
rect 69926 327218 100410 327454
rect 100646 327218 131130 327454
rect 131366 327218 161850 327454
rect 162086 327218 192570 327454
rect 192806 327218 223290 327454
rect 223526 327218 254010 327454
rect 254246 327218 284730 327454
rect 284966 327218 315450 327454
rect 315686 327218 346170 327454
rect 346406 327218 376890 327454
rect 377126 327218 407610 327454
rect 407846 327218 438330 327454
rect 438566 327218 469050 327454
rect 469286 327218 499770 327454
rect 500006 327218 530490 327454
rect 530726 327218 561210 327454
rect 561446 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 8250 327134
rect 8486 326898 38970 327134
rect 39206 326898 69690 327134
rect 69926 326898 100410 327134
rect 100646 326898 131130 327134
rect 131366 326898 161850 327134
rect 162086 326898 192570 327134
rect 192806 326898 223290 327134
rect 223526 326898 254010 327134
rect 254246 326898 284730 327134
rect 284966 326898 315450 327134
rect 315686 326898 346170 327134
rect 346406 326898 376890 327134
rect 377126 326898 407610 327134
rect 407846 326898 438330 327134
rect 438566 326898 469050 327134
rect 469286 326898 499770 327134
rect 500006 326898 530490 327134
rect 530726 326898 561210 327134
rect 561446 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect -8726 320294 592650 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect -6806 316574 590730 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect -4886 312854 588810 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 23610 309454
rect 23846 309218 54330 309454
rect 54566 309218 85050 309454
rect 85286 309218 115770 309454
rect 116006 309218 146490 309454
rect 146726 309218 177210 309454
rect 177446 309218 207930 309454
rect 208166 309218 238650 309454
rect 238886 309218 269370 309454
rect 269606 309218 300090 309454
rect 300326 309218 330810 309454
rect 331046 309218 361530 309454
rect 361766 309218 392250 309454
rect 392486 309218 422970 309454
rect 423206 309218 453690 309454
rect 453926 309218 484410 309454
rect 484646 309218 515130 309454
rect 515366 309218 545850 309454
rect 546086 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect -2966 309134 586890 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 23610 309134
rect 23846 308898 54330 309134
rect 54566 308898 85050 309134
rect 85286 308898 115770 309134
rect 116006 308898 146490 309134
rect 146726 308898 177210 309134
rect 177446 308898 207930 309134
rect 208166 308898 238650 309134
rect 238886 308898 269370 309134
rect 269606 308898 300090 309134
rect 300326 308898 330810 309134
rect 331046 308898 361530 309134
rect 361766 308898 392250 309134
rect 392486 308898 422970 309134
rect 423206 308898 453690 309134
rect 453926 308898 484410 309134
rect 484646 308898 515130 309134
rect 515366 308898 545850 309134
rect 546086 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect -2966 308866 586890 308898
rect -8726 302614 592650 302646
rect -8726 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 592650 302294
rect -8726 302026 592650 302058
rect -6806 298894 590730 298926
rect -6806 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 590730 298894
rect -6806 298574 590730 298658
rect -6806 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 590730 298574
rect -6806 298306 590730 298338
rect -4886 295174 588810 295206
rect -4886 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 588810 295174
rect -4886 294854 588810 294938
rect -4886 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 588810 294854
rect -4886 294586 588810 294618
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 8250 291454
rect 8486 291218 38970 291454
rect 39206 291218 69690 291454
rect 69926 291218 100410 291454
rect 100646 291218 131130 291454
rect 131366 291218 161850 291454
rect 162086 291218 192570 291454
rect 192806 291218 223290 291454
rect 223526 291218 254010 291454
rect 254246 291218 284730 291454
rect 284966 291218 315450 291454
rect 315686 291218 346170 291454
rect 346406 291218 376890 291454
rect 377126 291218 407610 291454
rect 407846 291218 438330 291454
rect 438566 291218 469050 291454
rect 469286 291218 499770 291454
rect 500006 291218 530490 291454
rect 530726 291218 561210 291454
rect 561446 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 8250 291134
rect 8486 290898 38970 291134
rect 39206 290898 69690 291134
rect 69926 290898 100410 291134
rect 100646 290898 131130 291134
rect 131366 290898 161850 291134
rect 162086 290898 192570 291134
rect 192806 290898 223290 291134
rect 223526 290898 254010 291134
rect 254246 290898 284730 291134
rect 284966 290898 315450 291134
rect 315686 290898 346170 291134
rect 346406 290898 376890 291134
rect 377126 290898 407610 291134
rect 407846 290898 438330 291134
rect 438566 290898 469050 291134
rect 469286 290898 499770 291134
rect 500006 290898 530490 291134
rect 530726 290898 561210 291134
rect 561446 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect -8726 284294 592650 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect -6806 280574 590730 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect -4886 276854 588810 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect -4886 276586 588810 276618
rect -2966 273454 586890 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 23610 273454
rect 23846 273218 54330 273454
rect 54566 273218 85050 273454
rect 85286 273218 115770 273454
rect 116006 273218 146490 273454
rect 146726 273218 177210 273454
rect 177446 273218 207930 273454
rect 208166 273218 238650 273454
rect 238886 273218 269370 273454
rect 269606 273218 300090 273454
rect 300326 273218 330810 273454
rect 331046 273218 361530 273454
rect 361766 273218 392250 273454
rect 392486 273218 422970 273454
rect 423206 273218 453690 273454
rect 453926 273218 484410 273454
rect 484646 273218 515130 273454
rect 515366 273218 545850 273454
rect 546086 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect -2966 273134 586890 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 23610 273134
rect 23846 272898 54330 273134
rect 54566 272898 85050 273134
rect 85286 272898 115770 273134
rect 116006 272898 146490 273134
rect 146726 272898 177210 273134
rect 177446 272898 207930 273134
rect 208166 272898 238650 273134
rect 238886 272898 269370 273134
rect 269606 272898 300090 273134
rect 300326 272898 330810 273134
rect 331046 272898 361530 273134
rect 361766 272898 392250 273134
rect 392486 272898 422970 273134
rect 423206 272898 453690 273134
rect 453926 272898 484410 273134
rect 484646 272898 515130 273134
rect 515366 272898 545850 273134
rect 546086 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 592650 266294
rect -8726 266026 592650 266058
rect -6806 262894 590730 262926
rect -6806 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 590730 262894
rect -6806 262574 590730 262658
rect -6806 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 590730 262574
rect -6806 262306 590730 262338
rect -4886 259174 588810 259206
rect -4886 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 588810 259174
rect -4886 258854 588810 258938
rect -4886 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 588810 258854
rect -4886 258586 588810 258618
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 8250 255454
rect 8486 255218 38970 255454
rect 39206 255218 69690 255454
rect 69926 255218 100410 255454
rect 100646 255218 131130 255454
rect 131366 255218 161850 255454
rect 162086 255218 192570 255454
rect 192806 255218 223290 255454
rect 223526 255218 254010 255454
rect 254246 255218 284730 255454
rect 284966 255218 315450 255454
rect 315686 255218 346170 255454
rect 346406 255218 376890 255454
rect 377126 255218 407610 255454
rect 407846 255218 438330 255454
rect 438566 255218 469050 255454
rect 469286 255218 499770 255454
rect 500006 255218 530490 255454
rect 530726 255218 561210 255454
rect 561446 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 8250 255134
rect 8486 254898 38970 255134
rect 39206 254898 69690 255134
rect 69926 254898 100410 255134
rect 100646 254898 131130 255134
rect 131366 254898 161850 255134
rect 162086 254898 192570 255134
rect 192806 254898 223290 255134
rect 223526 254898 254010 255134
rect 254246 254898 284730 255134
rect 284966 254898 315450 255134
rect 315686 254898 346170 255134
rect 346406 254898 376890 255134
rect 377126 254898 407610 255134
rect 407846 254898 438330 255134
rect 438566 254898 469050 255134
rect 469286 254898 499770 255134
rect 500006 254898 530490 255134
rect 530726 254898 561210 255134
rect 561446 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -8726 248614 592650 248646
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect -8726 248294 592650 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect -6806 244574 590730 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect -4886 240854 588810 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 23610 237454
rect 23846 237218 54330 237454
rect 54566 237218 85050 237454
rect 85286 237218 115770 237454
rect 116006 237218 146490 237454
rect 146726 237218 177210 237454
rect 177446 237218 207930 237454
rect 208166 237218 238650 237454
rect 238886 237218 269370 237454
rect 269606 237218 300090 237454
rect 300326 237218 330810 237454
rect 331046 237218 361530 237454
rect 361766 237218 392250 237454
rect 392486 237218 422970 237454
rect 423206 237218 453690 237454
rect 453926 237218 484410 237454
rect 484646 237218 515130 237454
rect 515366 237218 545850 237454
rect 546086 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect -2966 237134 586890 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 23610 237134
rect 23846 236898 54330 237134
rect 54566 236898 85050 237134
rect 85286 236898 115770 237134
rect 116006 236898 146490 237134
rect 146726 236898 177210 237134
rect 177446 236898 207930 237134
rect 208166 236898 238650 237134
rect 238886 236898 269370 237134
rect 269606 236898 300090 237134
rect 300326 236898 330810 237134
rect 331046 236898 361530 237134
rect 361766 236898 392250 237134
rect 392486 236898 422970 237134
rect 423206 236898 453690 237134
rect 453926 236898 484410 237134
rect 484646 236898 515130 237134
rect 515366 236898 545850 237134
rect 546086 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 592650 230294
rect -8726 230026 592650 230058
rect -6806 226894 590730 226926
rect -6806 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 590730 226894
rect -6806 226574 590730 226658
rect -6806 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 590730 226574
rect -6806 226306 590730 226338
rect -4886 223174 588810 223206
rect -4886 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 588810 223174
rect -4886 222854 588810 222938
rect -4886 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 588810 222854
rect -4886 222586 588810 222618
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 8250 219454
rect 8486 219218 38970 219454
rect 39206 219218 69690 219454
rect 69926 219218 100410 219454
rect 100646 219218 131130 219454
rect 131366 219218 161850 219454
rect 162086 219218 192570 219454
rect 192806 219218 223290 219454
rect 223526 219218 254010 219454
rect 254246 219218 284730 219454
rect 284966 219218 315450 219454
rect 315686 219218 346170 219454
rect 346406 219218 376890 219454
rect 377126 219218 407610 219454
rect 407846 219218 438330 219454
rect 438566 219218 469050 219454
rect 469286 219218 499770 219454
rect 500006 219218 530490 219454
rect 530726 219218 561210 219454
rect 561446 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 8250 219134
rect 8486 218898 38970 219134
rect 39206 218898 69690 219134
rect 69926 218898 100410 219134
rect 100646 218898 131130 219134
rect 131366 218898 161850 219134
rect 162086 218898 192570 219134
rect 192806 218898 223290 219134
rect 223526 218898 254010 219134
rect 254246 218898 284730 219134
rect 284966 218898 315450 219134
rect 315686 218898 346170 219134
rect 346406 218898 376890 219134
rect 377126 218898 407610 219134
rect 407846 218898 438330 219134
rect 438566 218898 469050 219134
rect 469286 218898 499770 219134
rect 500006 218898 530490 219134
rect 530726 218898 561210 219134
rect 561446 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -8726 212614 592650 212646
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect -8726 212294 592650 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect -6806 208574 590730 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect -4886 204854 588810 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 23610 201454
rect 23846 201218 54330 201454
rect 54566 201218 85050 201454
rect 85286 201218 115770 201454
rect 116006 201218 146490 201454
rect 146726 201218 177210 201454
rect 177446 201218 207930 201454
rect 208166 201218 238650 201454
rect 238886 201218 269370 201454
rect 269606 201218 300090 201454
rect 300326 201218 330810 201454
rect 331046 201218 361530 201454
rect 361766 201218 392250 201454
rect 392486 201218 422970 201454
rect 423206 201218 453690 201454
rect 453926 201218 484410 201454
rect 484646 201218 515130 201454
rect 515366 201218 545850 201454
rect 546086 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect -2966 201134 586890 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 23610 201134
rect 23846 200898 54330 201134
rect 54566 200898 85050 201134
rect 85286 200898 115770 201134
rect 116006 200898 146490 201134
rect 146726 200898 177210 201134
rect 177446 200898 207930 201134
rect 208166 200898 238650 201134
rect 238886 200898 269370 201134
rect 269606 200898 300090 201134
rect 300326 200898 330810 201134
rect 331046 200898 361530 201134
rect 361766 200898 392250 201134
rect 392486 200898 422970 201134
rect 423206 200898 453690 201134
rect 453926 200898 484410 201134
rect 484646 200898 515130 201134
rect 515366 200898 545850 201134
rect 546086 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 592650 194294
rect -8726 194026 592650 194058
rect -6806 190894 590730 190926
rect -6806 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 590730 190894
rect -6806 190574 590730 190658
rect -6806 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 590730 190574
rect -6806 190306 590730 190338
rect -4886 187174 588810 187206
rect -4886 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 588810 187174
rect -4886 186854 588810 186938
rect -4886 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 588810 186854
rect -4886 186586 588810 186618
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 8250 183454
rect 8486 183218 38970 183454
rect 39206 183218 69690 183454
rect 69926 183218 100410 183454
rect 100646 183218 131130 183454
rect 131366 183218 161850 183454
rect 162086 183218 192570 183454
rect 192806 183218 223290 183454
rect 223526 183218 254010 183454
rect 254246 183218 284730 183454
rect 284966 183218 315450 183454
rect 315686 183218 346170 183454
rect 346406 183218 376890 183454
rect 377126 183218 407610 183454
rect 407846 183218 438330 183454
rect 438566 183218 469050 183454
rect 469286 183218 499770 183454
rect 500006 183218 530490 183454
rect 530726 183218 561210 183454
rect 561446 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 8250 183134
rect 8486 182898 38970 183134
rect 39206 182898 69690 183134
rect 69926 182898 100410 183134
rect 100646 182898 131130 183134
rect 131366 182898 161850 183134
rect 162086 182898 192570 183134
rect 192806 182898 223290 183134
rect 223526 182898 254010 183134
rect 254246 182898 284730 183134
rect 284966 182898 315450 183134
rect 315686 182898 346170 183134
rect 346406 182898 376890 183134
rect 377126 182898 407610 183134
rect 407846 182898 438330 183134
rect 438566 182898 469050 183134
rect 469286 182898 499770 183134
rect 500006 182898 530490 183134
rect 530726 182898 561210 183134
rect 561446 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect -8726 176614 592650 176646
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect -8726 176294 592650 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect -8726 176026 592650 176058
rect -6806 172894 590730 172926
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect -6806 172574 590730 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect -6806 172306 590730 172338
rect -4886 169174 588810 169206
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect -4886 168854 588810 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect -4886 168586 588810 168618
rect -2966 165454 586890 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 23610 165454
rect 23846 165218 54330 165454
rect 54566 165218 85050 165454
rect 85286 165218 115770 165454
rect 116006 165218 146490 165454
rect 146726 165218 177210 165454
rect 177446 165218 207930 165454
rect 208166 165218 238650 165454
rect 238886 165218 269370 165454
rect 269606 165218 300090 165454
rect 300326 165218 330810 165454
rect 331046 165218 361530 165454
rect 361766 165218 392250 165454
rect 392486 165218 422970 165454
rect 423206 165218 453690 165454
rect 453926 165218 484410 165454
rect 484646 165218 515130 165454
rect 515366 165218 545850 165454
rect 546086 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect -2966 165134 586890 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 23610 165134
rect 23846 164898 54330 165134
rect 54566 164898 85050 165134
rect 85286 164898 115770 165134
rect 116006 164898 146490 165134
rect 146726 164898 177210 165134
rect 177446 164898 207930 165134
rect 208166 164898 238650 165134
rect 238886 164898 269370 165134
rect 269606 164898 300090 165134
rect 300326 164898 330810 165134
rect 331046 164898 361530 165134
rect 361766 164898 392250 165134
rect 392486 164898 422970 165134
rect 423206 164898 453690 165134
rect 453926 164898 484410 165134
rect 484646 164898 515130 165134
rect 515366 164898 545850 165134
rect 546086 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect -2966 164866 586890 164898
rect -8726 158614 592650 158646
rect -8726 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 592650 158294
rect -8726 158026 592650 158058
rect -6806 154894 590730 154926
rect -6806 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 590730 154894
rect -6806 154574 590730 154658
rect -6806 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 590730 154574
rect -6806 154306 590730 154338
rect -4886 151174 588810 151206
rect -4886 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 588810 151174
rect -4886 150854 588810 150938
rect -4886 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 588810 150854
rect -4886 150586 588810 150618
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 8250 147454
rect 8486 147218 38970 147454
rect 39206 147218 69690 147454
rect 69926 147218 100410 147454
rect 100646 147218 131130 147454
rect 131366 147218 161850 147454
rect 162086 147218 192570 147454
rect 192806 147218 223290 147454
rect 223526 147218 254010 147454
rect 254246 147218 284730 147454
rect 284966 147218 315450 147454
rect 315686 147218 346170 147454
rect 346406 147218 376890 147454
rect 377126 147218 407610 147454
rect 407846 147218 438330 147454
rect 438566 147218 469050 147454
rect 469286 147218 499770 147454
rect 500006 147218 530490 147454
rect 530726 147218 561210 147454
rect 561446 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 8250 147134
rect 8486 146898 38970 147134
rect 39206 146898 69690 147134
rect 69926 146898 100410 147134
rect 100646 146898 131130 147134
rect 131366 146898 161850 147134
rect 162086 146898 192570 147134
rect 192806 146898 223290 147134
rect 223526 146898 254010 147134
rect 254246 146898 284730 147134
rect 284966 146898 315450 147134
rect 315686 146898 346170 147134
rect 346406 146898 376890 147134
rect 377126 146898 407610 147134
rect 407846 146898 438330 147134
rect 438566 146898 469050 147134
rect 469286 146898 499770 147134
rect 500006 146898 530490 147134
rect 530726 146898 561210 147134
rect 561446 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -8726 140614 592650 140646
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect -8726 140294 592650 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect -8726 140026 592650 140058
rect -6806 136894 590730 136926
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect -6806 136574 590730 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect -6806 136306 590730 136338
rect -4886 133174 588810 133206
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect -4886 132854 588810 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect -4886 132586 588810 132618
rect -2966 129454 586890 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 23610 129454
rect 23846 129218 54330 129454
rect 54566 129218 85050 129454
rect 85286 129218 115770 129454
rect 116006 129218 146490 129454
rect 146726 129218 177210 129454
rect 177446 129218 207930 129454
rect 208166 129218 238650 129454
rect 238886 129218 269370 129454
rect 269606 129218 300090 129454
rect 300326 129218 330810 129454
rect 331046 129218 361530 129454
rect 361766 129218 392250 129454
rect 392486 129218 422970 129454
rect 423206 129218 453690 129454
rect 453926 129218 484410 129454
rect 484646 129218 515130 129454
rect 515366 129218 545850 129454
rect 546086 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect -2966 129134 586890 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 23610 129134
rect 23846 128898 54330 129134
rect 54566 128898 85050 129134
rect 85286 128898 115770 129134
rect 116006 128898 146490 129134
rect 146726 128898 177210 129134
rect 177446 128898 207930 129134
rect 208166 128898 238650 129134
rect 238886 128898 269370 129134
rect 269606 128898 300090 129134
rect 300326 128898 330810 129134
rect 331046 128898 361530 129134
rect 361766 128898 392250 129134
rect 392486 128898 422970 129134
rect 423206 128898 453690 129134
rect 453926 128898 484410 129134
rect 484646 128898 515130 129134
rect 515366 128898 545850 129134
rect 546086 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect -2966 128866 586890 128898
rect -8726 122614 592650 122646
rect -8726 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 592650 122294
rect -8726 122026 592650 122058
rect -6806 118894 590730 118926
rect -6806 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 590730 118894
rect -6806 118574 590730 118658
rect -6806 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 590730 118574
rect -6806 118306 590730 118338
rect -4886 115174 588810 115206
rect -4886 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 588810 115174
rect -4886 114854 588810 114938
rect -4886 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 588810 114854
rect -4886 114586 588810 114618
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 8250 111454
rect 8486 111218 38970 111454
rect 39206 111218 69690 111454
rect 69926 111218 100410 111454
rect 100646 111218 131130 111454
rect 131366 111218 161850 111454
rect 162086 111218 192570 111454
rect 192806 111218 223290 111454
rect 223526 111218 254010 111454
rect 254246 111218 284730 111454
rect 284966 111218 315450 111454
rect 315686 111218 346170 111454
rect 346406 111218 376890 111454
rect 377126 111218 407610 111454
rect 407846 111218 438330 111454
rect 438566 111218 469050 111454
rect 469286 111218 499770 111454
rect 500006 111218 530490 111454
rect 530726 111218 561210 111454
rect 561446 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 8250 111134
rect 8486 110898 38970 111134
rect 39206 110898 69690 111134
rect 69926 110898 100410 111134
rect 100646 110898 131130 111134
rect 131366 110898 161850 111134
rect 162086 110898 192570 111134
rect 192806 110898 223290 111134
rect 223526 110898 254010 111134
rect 254246 110898 284730 111134
rect 284966 110898 315450 111134
rect 315686 110898 346170 111134
rect 346406 110898 376890 111134
rect 377126 110898 407610 111134
rect 407846 110898 438330 111134
rect 438566 110898 469050 111134
rect 469286 110898 499770 111134
rect 500006 110898 530490 111134
rect 530726 110898 561210 111134
rect 561446 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -8726 104614 592650 104646
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect -8726 104294 592650 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect -8726 104026 592650 104058
rect -6806 100894 590730 100926
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect -6806 100574 590730 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect -6806 100306 590730 100338
rect -4886 97174 588810 97206
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect -4886 96854 588810 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect -4886 96586 588810 96618
rect -2966 93454 586890 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 23610 93454
rect 23846 93218 54330 93454
rect 54566 93218 85050 93454
rect 85286 93218 115770 93454
rect 116006 93218 146490 93454
rect 146726 93218 177210 93454
rect 177446 93218 207930 93454
rect 208166 93218 238650 93454
rect 238886 93218 269370 93454
rect 269606 93218 300090 93454
rect 300326 93218 330810 93454
rect 331046 93218 361530 93454
rect 361766 93218 392250 93454
rect 392486 93218 422970 93454
rect 423206 93218 453690 93454
rect 453926 93218 484410 93454
rect 484646 93218 515130 93454
rect 515366 93218 545850 93454
rect 546086 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect -2966 93134 586890 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 23610 93134
rect 23846 92898 54330 93134
rect 54566 92898 85050 93134
rect 85286 92898 115770 93134
rect 116006 92898 146490 93134
rect 146726 92898 177210 93134
rect 177446 92898 207930 93134
rect 208166 92898 238650 93134
rect 238886 92898 269370 93134
rect 269606 92898 300090 93134
rect 300326 92898 330810 93134
rect 331046 92898 361530 93134
rect 361766 92898 392250 93134
rect 392486 92898 422970 93134
rect 423206 92898 453690 93134
rect 453926 92898 484410 93134
rect 484646 92898 515130 93134
rect 515366 92898 545850 93134
rect 546086 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect -2966 92866 586890 92898
rect -8726 86614 592650 86646
rect -8726 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 592650 86294
rect -8726 86026 592650 86058
rect -6806 82894 590730 82926
rect -6806 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 590730 82894
rect -6806 82574 590730 82658
rect -6806 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 590730 82574
rect -6806 82306 590730 82338
rect -4886 79174 588810 79206
rect -4886 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 588810 79174
rect -4886 78854 588810 78938
rect -4886 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 588810 78854
rect -4886 78586 588810 78618
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 8250 75454
rect 8486 75218 38970 75454
rect 39206 75218 69690 75454
rect 69926 75218 100410 75454
rect 100646 75218 131130 75454
rect 131366 75218 161850 75454
rect 162086 75218 192570 75454
rect 192806 75218 223290 75454
rect 223526 75218 254010 75454
rect 254246 75218 284730 75454
rect 284966 75218 315450 75454
rect 315686 75218 346170 75454
rect 346406 75218 376890 75454
rect 377126 75218 407610 75454
rect 407846 75218 438330 75454
rect 438566 75218 469050 75454
rect 469286 75218 499770 75454
rect 500006 75218 530490 75454
rect 530726 75218 561210 75454
rect 561446 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 8250 75134
rect 8486 74898 38970 75134
rect 39206 74898 69690 75134
rect 69926 74898 100410 75134
rect 100646 74898 131130 75134
rect 131366 74898 161850 75134
rect 162086 74898 192570 75134
rect 192806 74898 223290 75134
rect 223526 74898 254010 75134
rect 254246 74898 284730 75134
rect 284966 74898 315450 75134
rect 315686 74898 346170 75134
rect 346406 74898 376890 75134
rect 377126 74898 407610 75134
rect 407846 74898 438330 75134
rect 438566 74898 469050 75134
rect 469286 74898 499770 75134
rect 500006 74898 530490 75134
rect 530726 74898 561210 75134
rect 561446 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -8726 68614 592650 68646
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect -8726 68294 592650 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect -8726 68026 592650 68058
rect -6806 64894 590730 64926
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect -6806 64574 590730 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect -6806 64306 590730 64338
rect -4886 61174 588810 61206
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect -4886 60854 588810 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect -4886 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 23610 57454
rect 23846 57218 54330 57454
rect 54566 57218 85050 57454
rect 85286 57218 115770 57454
rect 116006 57218 146490 57454
rect 146726 57218 177210 57454
rect 177446 57218 207930 57454
rect 208166 57218 238650 57454
rect 238886 57218 269370 57454
rect 269606 57218 300090 57454
rect 300326 57218 330810 57454
rect 331046 57218 361530 57454
rect 361766 57218 392250 57454
rect 392486 57218 422970 57454
rect 423206 57218 453690 57454
rect 453926 57218 484410 57454
rect 484646 57218 515130 57454
rect 515366 57218 545850 57454
rect 546086 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 23610 57134
rect 23846 56898 54330 57134
rect 54566 56898 85050 57134
rect 85286 56898 115770 57134
rect 116006 56898 146490 57134
rect 146726 56898 177210 57134
rect 177446 56898 207930 57134
rect 208166 56898 238650 57134
rect 238886 56898 269370 57134
rect 269606 56898 300090 57134
rect 300326 56898 330810 57134
rect 331046 56898 361530 57134
rect 361766 56898 392250 57134
rect 392486 56898 422970 57134
rect 423206 56898 453690 57134
rect 453926 56898 484410 57134
rect 484646 56898 515130 57134
rect 515366 56898 545850 57134
rect 546086 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 592650 50294
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 590730 46894
rect -6806 46574 590730 46658
rect -6806 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 590730 46574
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 588810 43174
rect -4886 42854 588810 42938
rect -4886 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 588810 42854
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 8250 39454
rect 8486 39218 38970 39454
rect 39206 39218 69690 39454
rect 69926 39218 100410 39454
rect 100646 39218 131130 39454
rect 131366 39218 161850 39454
rect 162086 39218 192570 39454
rect 192806 39218 223290 39454
rect 223526 39218 254010 39454
rect 254246 39218 284730 39454
rect 284966 39218 315450 39454
rect 315686 39218 346170 39454
rect 346406 39218 376890 39454
rect 377126 39218 407610 39454
rect 407846 39218 438330 39454
rect 438566 39218 469050 39454
rect 469286 39218 499770 39454
rect 500006 39218 530490 39454
rect 530726 39218 561210 39454
rect 561446 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 8250 39134
rect 8486 38898 38970 39134
rect 39206 38898 69690 39134
rect 69926 38898 100410 39134
rect 100646 38898 131130 39134
rect 131366 38898 161850 39134
rect 162086 38898 192570 39134
rect 192806 38898 223290 39134
rect 223526 38898 254010 39134
rect 254246 38898 284730 39134
rect 284966 38898 315450 39134
rect 315686 38898 346170 39134
rect 346406 38898 376890 39134
rect 377126 38898 407610 39134
rect 407846 38898 438330 39134
rect 438566 38898 469050 39134
rect 469286 38898 499770 39134
rect 500006 38898 530490 39134
rect 530726 38898 561210 39134
rect 561446 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect -8726 32294 592650 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect -6806 28574 590730 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect -4886 24854 588810 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 23610 21454
rect 23846 21218 54330 21454
rect 54566 21218 85050 21454
rect 85286 21218 115770 21454
rect 116006 21218 146490 21454
rect 146726 21218 177210 21454
rect 177446 21218 207930 21454
rect 208166 21218 238650 21454
rect 238886 21218 269370 21454
rect 269606 21218 300090 21454
rect 300326 21218 330810 21454
rect 331046 21218 361530 21454
rect 361766 21218 392250 21454
rect 392486 21218 422970 21454
rect 423206 21218 453690 21454
rect 453926 21218 484410 21454
rect 484646 21218 515130 21454
rect 515366 21218 545850 21454
rect 546086 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 23610 21134
rect 23846 20898 54330 21134
rect 54566 20898 85050 21134
rect 85286 20898 115770 21134
rect 116006 20898 146490 21134
rect 146726 20898 177210 21134
rect 177446 20898 207930 21134
rect 208166 20898 238650 21134
rect 238886 20898 269370 21134
rect 269606 20898 300090 21134
rect 300326 20898 330810 21134
rect 331046 20898 361530 21134
rect 361766 20898 392250 21134
rect 392486 20898 422970 21134
rect 423206 20898 453690 21134
rect 453926 20898 484410 21134
rect 484646 20898 515130 21134
rect 515366 20898 545850 21134
rect 546086 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 592650 14294
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 590730 10894
rect -6806 10574 590730 10658
rect -6806 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 590730 10574
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 588810 7174
rect -4886 6854 588810 6938
rect -4886 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 588810 6854
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 8250 3454
rect 8486 3218 38970 3454
rect 39206 3218 69690 3454
rect 69926 3218 100410 3454
rect 100646 3218 131130 3454
rect 131366 3218 161850 3454
rect 162086 3218 192570 3454
rect 192806 3218 223290 3454
rect 223526 3218 254010 3454
rect 254246 3218 284730 3454
rect 284966 3218 315450 3454
rect 315686 3218 346170 3454
rect 346406 3218 376890 3454
rect 377126 3218 407610 3454
rect 407846 3218 438330 3454
rect 438566 3218 469050 3454
rect 469286 3218 499770 3454
rect 500006 3218 530490 3454
rect 530726 3218 561210 3454
rect 561446 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 8250 3134
rect 8486 2898 38970 3134
rect 39206 2898 69690 3134
rect 69926 2898 100410 3134
rect 100646 2898 131130 3134
rect 131366 2898 161850 3134
rect 162086 2898 192570 3134
rect 192806 2898 223290 3134
rect 223526 2898 254010 3134
rect 254246 2898 284730 3134
rect 284966 2898 315450 3134
rect 315686 2898 346170 3134
rect 346406 2898 376890 3134
rect 377126 2898 407610 3134
rect 407846 2898 438330 3134
rect 438566 2898 469050 3134
rect 469286 2898 499770 3134
rect 500006 2898 530490 3134
rect 530726 2898 561210 3134
rect 561446 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use user_proj  mprj
timestamp 1639754316
transform 1 0 4000 0 1 0
box 566 0 559438 700000
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 702000 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 702000 38414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 702000 74414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 702000 110414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 702000 146414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 702000 182414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 702000 218414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 702000 254414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 702000 290414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 702000 326414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 702000 362414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 702000 398414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 702000 434414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 702000 470414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 702000 506414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 702000 542414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 -3814 6134 -2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 41514 -3814 42134 -2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 77514 -3814 78134 -2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 113514 -3814 114134 -2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 149514 -3814 150134 -2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 185514 -3814 186134 -2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 221514 -3814 222134 -2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 257514 -3814 258134 -2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 293514 -3814 294134 -2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 329514 -3814 330134 -2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 365514 -3814 366134 -2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 401514 -3814 402134 -2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 437514 -3814 438134 -2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 473514 -3814 474134 -2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 509514 -3814 510134 -2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 545514 -3814 546134 -2000 8 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 702000 6134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 702000 42134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 702000 78134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 702000 114134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 702000 150134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 702000 186134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 702000 222134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 702000 258134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 702000 294134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 702000 330134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 702000 366134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 702000 402134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 702000 438134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 702000 474134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 702000 510134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 702000 546134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 581514 -3814 582134 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 -5734 9854 -2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 45234 -5734 45854 -2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 81234 -5734 81854 -2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 117234 -5734 117854 -2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 153234 -5734 153854 -2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 189234 -5734 189854 -2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 225234 -5734 225854 -2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 261234 -5734 261854 -2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 297234 -5734 297854 -2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 333234 -5734 333854 -2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 369234 -5734 369854 -2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 405234 -5734 405854 -2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 441234 -5734 441854 -2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 477234 -5734 477854 -2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 513234 -5734 513854 -2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 549234 -5734 549854 -2000 8 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 702000 9854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 702000 45854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 702000 81854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 702000 117854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 702000 153854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 702000 189854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 702000 225854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 702000 261854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 702000 297854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 702000 333854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 702000 369854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 702000 405854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 702000 441854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 702000 477854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 702000 513854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 702000 549854 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 -7654 13574 -2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 48954 -7654 49574 -2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 84954 -7654 85574 -2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 120954 -7654 121574 -2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 156954 -7654 157574 -2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 192954 -7654 193574 -2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 228954 -7654 229574 -2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 264954 -7654 265574 -2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 300954 -7654 301574 -2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 336954 -7654 337574 -2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 372954 -7654 373574 -2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 408954 -7654 409574 -2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 444954 -7654 445574 -2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 480954 -7654 481574 -2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 516954 -7654 517574 -2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 552954 -7654 553574 -2000 8 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 702000 13574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 702000 49574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 702000 85574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 702000 121574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 702000 157574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 702000 193574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 702000 229574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 702000 265574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 702000 301574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 702000 337574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 702000 373574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 702000 409574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 702000 445574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 702000 481574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 702000 517574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 702000 553574 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 -5734 27854 -2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 -5734 63854 -2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 -5734 99854 -2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 -5734 135854 -2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 -5734 171854 -2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 -5734 207854 -2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 -5734 243854 -2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 -5734 279854 -2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 -5734 315854 -2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 -5734 351854 -2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 -5734 387854 -2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 -5734 423854 -2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 -5734 459854 -2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 -5734 495854 -2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 -5734 531854 -2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 702000 27854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 702000 63854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 702000 99854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 702000 135854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 702000 171854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 702000 207854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 702000 243854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 702000 279854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 702000 315854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 702000 351854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 702000 387854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 702000 423854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 702000 459854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 702000 495854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 702000 531854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 -5734 567854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 -7654 31574 -2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 -7654 67574 -2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 -7654 103574 -2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 -7654 139574 -2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 -7654 175574 -2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 -7654 211574 -2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 -7654 247574 -2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 -7654 283574 -2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 -7654 319574 -2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 -7654 355574 -2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 -7654 391574 -2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 -7654 427574 -2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 -7654 463574 -2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 -7654 499574 -2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 -7654 535574 -2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 702000 31574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 702000 67574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 702000 103574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 702000 139574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 702000 175574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 702000 211574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 702000 247574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 702000 283574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 702000 319574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 702000 355574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 702000 391574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 702000 427574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 702000 463574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 702000 499574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 702000 535574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 -7654 571574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 702000 20414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 702000 56414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 702000 92414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 702000 128414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 702000 164414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 702000 200414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 702000 236414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 702000 272414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 702000 308414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 702000 344414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 702000 380414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 702000 416414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 702000 452414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 702000 488414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 702000 524414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 702000 560414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 -3814 24134 -2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 -3814 60134 -2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 -3814 96134 -2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 -3814 132134 -2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 -3814 168134 -2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 -3814 204134 -2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 -3814 240134 -2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 -3814 276134 -2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 -3814 312134 -2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 -3814 348134 -2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 -3814 384134 -2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 -3814 420134 -2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 -3814 456134 -2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 -3814 492134 -2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 -3814 528134 -2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 -3814 564134 -2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 702000 24134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 702000 60134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 702000 96134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 702000 132134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 702000 168134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 702000 204134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 702000 240134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 702000 276134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 702000 312134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 702000 348134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 702000 384134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 702000 420134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 702000 456134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 702000 492134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 702000 528134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 702000 564134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
