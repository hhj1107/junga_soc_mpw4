magic
tech sky130A
magscale 1 2
timestamp 1640370137
<< obsli1 >>
rect 1104 1649 164467 164305
<< obsm1 >>
rect 106 484 164482 164336
<< metal2 >>
rect 478 165875 534 166675
rect 1398 165875 1454 166675
rect 2318 165875 2374 166675
rect 3330 165875 3386 166675
rect 4250 165875 4306 166675
rect 5170 165875 5226 166675
rect 6182 165875 6238 166675
rect 7102 165875 7158 166675
rect 8022 165875 8078 166675
rect 9034 165875 9090 166675
rect 9954 165875 10010 166675
rect 10874 165875 10930 166675
rect 11886 165875 11942 166675
rect 12806 165875 12862 166675
rect 13726 165875 13782 166675
rect 14738 165875 14794 166675
rect 15658 165875 15714 166675
rect 16578 165875 16634 166675
rect 17590 165875 17646 166675
rect 18510 165875 18566 166675
rect 19430 165875 19486 166675
rect 20442 165875 20498 166675
rect 21362 165875 21418 166675
rect 22282 165875 22338 166675
rect 23294 165875 23350 166675
rect 24214 165875 24270 166675
rect 25134 165875 25190 166675
rect 26146 165875 26202 166675
rect 27066 165875 27122 166675
rect 27986 165875 28042 166675
rect 28998 165875 29054 166675
rect 29918 165875 29974 166675
rect 30838 165875 30894 166675
rect 31850 165875 31906 166675
rect 32770 165875 32826 166675
rect 33690 165875 33746 166675
rect 34702 165875 34758 166675
rect 35622 165875 35678 166675
rect 36542 165875 36598 166675
rect 37554 165875 37610 166675
rect 38474 165875 38530 166675
rect 39394 165875 39450 166675
rect 40406 165875 40462 166675
rect 41326 165875 41382 166675
rect 42246 165875 42302 166675
rect 43258 165875 43314 166675
rect 44178 165875 44234 166675
rect 45098 165875 45154 166675
rect 46110 165875 46166 166675
rect 47030 165875 47086 166675
rect 47950 165875 48006 166675
rect 48962 165875 49018 166675
rect 49882 165875 49938 166675
rect 50802 165875 50858 166675
rect 51814 165875 51870 166675
rect 52734 165875 52790 166675
rect 53654 165875 53710 166675
rect 54666 165875 54722 166675
rect 55586 165875 55642 166675
rect 56506 165875 56562 166675
rect 57518 165875 57574 166675
rect 58438 165875 58494 166675
rect 59358 165875 59414 166675
rect 60370 165875 60426 166675
rect 61290 165875 61346 166675
rect 62210 165875 62266 166675
rect 63222 165875 63278 166675
rect 64142 165875 64198 166675
rect 65062 165875 65118 166675
rect 66074 165875 66130 166675
rect 66994 165875 67050 166675
rect 67914 165875 67970 166675
rect 68926 165875 68982 166675
rect 69846 165875 69902 166675
rect 70766 165875 70822 166675
rect 71778 165875 71834 166675
rect 72698 165875 72754 166675
rect 73618 165875 73674 166675
rect 74630 165875 74686 166675
rect 75550 165875 75606 166675
rect 76470 165875 76526 166675
rect 77482 165875 77538 166675
rect 78402 165875 78458 166675
rect 79322 165875 79378 166675
rect 80334 165875 80390 166675
rect 81254 165875 81310 166675
rect 82174 165875 82230 166675
rect 83186 165875 83242 166675
rect 84106 165875 84162 166675
rect 85026 165875 85082 166675
rect 86038 165875 86094 166675
rect 86958 165875 87014 166675
rect 87878 165875 87934 166675
rect 88890 165875 88946 166675
rect 89810 165875 89866 166675
rect 90730 165875 90786 166675
rect 91742 165875 91798 166675
rect 92662 165875 92718 166675
rect 93582 165875 93638 166675
rect 94594 165875 94650 166675
rect 95514 165875 95570 166675
rect 96434 165875 96490 166675
rect 97446 165875 97502 166675
rect 98366 165875 98422 166675
rect 99286 165875 99342 166675
rect 100298 165875 100354 166675
rect 101218 165875 101274 166675
rect 102138 165875 102194 166675
rect 103150 165875 103206 166675
rect 104070 165875 104126 166675
rect 104990 165875 105046 166675
rect 106002 165875 106058 166675
rect 106922 165875 106978 166675
rect 107842 165875 107898 166675
rect 108854 165875 108910 166675
rect 109774 165875 109830 166675
rect 110694 165875 110750 166675
rect 111706 165875 111762 166675
rect 112626 165875 112682 166675
rect 113546 165875 113602 166675
rect 114558 165875 114614 166675
rect 115478 165875 115534 166675
rect 116398 165875 116454 166675
rect 117410 165875 117466 166675
rect 118330 165875 118386 166675
rect 119250 165875 119306 166675
rect 120262 165875 120318 166675
rect 121182 165875 121238 166675
rect 122102 165875 122158 166675
rect 123114 165875 123170 166675
rect 124034 165875 124090 166675
rect 124954 165875 125010 166675
rect 125966 165875 126022 166675
rect 126886 165875 126942 166675
rect 127806 165875 127862 166675
rect 128818 165875 128874 166675
rect 129738 165875 129794 166675
rect 130658 165875 130714 166675
rect 131670 165875 131726 166675
rect 132590 165875 132646 166675
rect 133510 165875 133566 166675
rect 134522 165875 134578 166675
rect 135442 165875 135498 166675
rect 136362 165875 136418 166675
rect 137374 165875 137430 166675
rect 138294 165875 138350 166675
rect 139214 165875 139270 166675
rect 140226 165875 140282 166675
rect 141146 165875 141202 166675
rect 142066 165875 142122 166675
rect 143078 165875 143134 166675
rect 143998 165875 144054 166675
rect 144918 165875 144974 166675
rect 145930 165875 145986 166675
rect 146850 165875 146906 166675
rect 147770 165875 147826 166675
rect 148782 165875 148838 166675
rect 149702 165875 149758 166675
rect 150622 165875 150678 166675
rect 151634 165875 151690 166675
rect 152554 165875 152610 166675
rect 153474 165875 153530 166675
rect 154486 165875 154542 166675
rect 155406 165875 155462 166675
rect 156326 165875 156382 166675
rect 157338 165875 157394 166675
rect 158258 165875 158314 166675
rect 159178 165875 159234 166675
rect 160190 165875 160246 166675
rect 161110 165875 161166 166675
rect 162030 165875 162086 166675
rect 163042 165875 163098 166675
rect 163962 165875 164018 166675
rect 110 0 166 800
rect 386 0 442 800
rect 662 0 718 800
rect 938 0 994 800
rect 1214 0 1270 800
rect 1582 0 1638 800
rect 1858 0 1914 800
rect 2134 0 2190 800
rect 2410 0 2466 800
rect 2778 0 2834 800
rect 3054 0 3110 800
rect 3330 0 3386 800
rect 3606 0 3662 800
rect 3974 0 4030 800
rect 4250 0 4306 800
rect 4526 0 4582 800
rect 4802 0 4858 800
rect 5170 0 5226 800
rect 5446 0 5502 800
rect 5722 0 5778 800
rect 5998 0 6054 800
rect 6366 0 6422 800
rect 6642 0 6698 800
rect 6918 0 6974 800
rect 7194 0 7250 800
rect 7470 0 7526 800
rect 7838 0 7894 800
rect 8114 0 8170 800
rect 8390 0 8446 800
rect 8666 0 8722 800
rect 9034 0 9090 800
rect 9310 0 9366 800
rect 9586 0 9642 800
rect 9862 0 9918 800
rect 10230 0 10286 800
rect 10506 0 10562 800
rect 10782 0 10838 800
rect 11058 0 11114 800
rect 11426 0 11482 800
rect 11702 0 11758 800
rect 11978 0 12034 800
rect 12254 0 12310 800
rect 12622 0 12678 800
rect 12898 0 12954 800
rect 13174 0 13230 800
rect 13450 0 13506 800
rect 13818 0 13874 800
rect 14094 0 14150 800
rect 14370 0 14426 800
rect 14646 0 14702 800
rect 14922 0 14978 800
rect 15290 0 15346 800
rect 15566 0 15622 800
rect 15842 0 15898 800
rect 16118 0 16174 800
rect 16486 0 16542 800
rect 16762 0 16818 800
rect 17038 0 17094 800
rect 17314 0 17370 800
rect 17682 0 17738 800
rect 17958 0 18014 800
rect 18234 0 18290 800
rect 18510 0 18566 800
rect 18878 0 18934 800
rect 19154 0 19210 800
rect 19430 0 19486 800
rect 19706 0 19762 800
rect 20074 0 20130 800
rect 20350 0 20406 800
rect 20626 0 20682 800
rect 20902 0 20958 800
rect 21178 0 21234 800
rect 21546 0 21602 800
rect 21822 0 21878 800
rect 22098 0 22154 800
rect 22374 0 22430 800
rect 22742 0 22798 800
rect 23018 0 23074 800
rect 23294 0 23350 800
rect 23570 0 23626 800
rect 23938 0 23994 800
rect 24214 0 24270 800
rect 24490 0 24546 800
rect 24766 0 24822 800
rect 25134 0 25190 800
rect 25410 0 25466 800
rect 25686 0 25742 800
rect 25962 0 26018 800
rect 26330 0 26386 800
rect 26606 0 26662 800
rect 26882 0 26938 800
rect 27158 0 27214 800
rect 27526 0 27582 800
rect 27802 0 27858 800
rect 28078 0 28134 800
rect 28354 0 28410 800
rect 28630 0 28686 800
rect 28998 0 29054 800
rect 29274 0 29330 800
rect 29550 0 29606 800
rect 29826 0 29882 800
rect 30194 0 30250 800
rect 30470 0 30526 800
rect 30746 0 30802 800
rect 31022 0 31078 800
rect 31390 0 31446 800
rect 31666 0 31722 800
rect 31942 0 31998 800
rect 32218 0 32274 800
rect 32586 0 32642 800
rect 32862 0 32918 800
rect 33138 0 33194 800
rect 33414 0 33470 800
rect 33782 0 33838 800
rect 34058 0 34114 800
rect 34334 0 34390 800
rect 34610 0 34666 800
rect 34886 0 34942 800
rect 35254 0 35310 800
rect 35530 0 35586 800
rect 35806 0 35862 800
rect 36082 0 36138 800
rect 36450 0 36506 800
rect 36726 0 36782 800
rect 37002 0 37058 800
rect 37278 0 37334 800
rect 37646 0 37702 800
rect 37922 0 37978 800
rect 38198 0 38254 800
rect 38474 0 38530 800
rect 38842 0 38898 800
rect 39118 0 39174 800
rect 39394 0 39450 800
rect 39670 0 39726 800
rect 40038 0 40094 800
rect 40314 0 40370 800
rect 40590 0 40646 800
rect 40866 0 40922 800
rect 41234 0 41290 800
rect 41510 0 41566 800
rect 41786 0 41842 800
rect 42062 0 42118 800
rect 42338 0 42394 800
rect 42706 0 42762 800
rect 42982 0 43038 800
rect 43258 0 43314 800
rect 43534 0 43590 800
rect 43902 0 43958 800
rect 44178 0 44234 800
rect 44454 0 44510 800
rect 44730 0 44786 800
rect 45098 0 45154 800
rect 45374 0 45430 800
rect 45650 0 45706 800
rect 45926 0 45982 800
rect 46294 0 46350 800
rect 46570 0 46626 800
rect 46846 0 46902 800
rect 47122 0 47178 800
rect 47490 0 47546 800
rect 47766 0 47822 800
rect 48042 0 48098 800
rect 48318 0 48374 800
rect 48594 0 48650 800
rect 48962 0 49018 800
rect 49238 0 49294 800
rect 49514 0 49570 800
rect 49790 0 49846 800
rect 50158 0 50214 800
rect 50434 0 50490 800
rect 50710 0 50766 800
rect 50986 0 51042 800
rect 51354 0 51410 800
rect 51630 0 51686 800
rect 51906 0 51962 800
rect 52182 0 52238 800
rect 52550 0 52606 800
rect 52826 0 52882 800
rect 53102 0 53158 800
rect 53378 0 53434 800
rect 53746 0 53802 800
rect 54022 0 54078 800
rect 54298 0 54354 800
rect 54574 0 54630 800
rect 54942 0 54998 800
rect 55218 0 55274 800
rect 55494 0 55550 800
rect 55770 0 55826 800
rect 56046 0 56102 800
rect 56414 0 56470 800
rect 56690 0 56746 800
rect 56966 0 57022 800
rect 57242 0 57298 800
rect 57610 0 57666 800
rect 57886 0 57942 800
rect 58162 0 58218 800
rect 58438 0 58494 800
rect 58806 0 58862 800
rect 59082 0 59138 800
rect 59358 0 59414 800
rect 59634 0 59690 800
rect 60002 0 60058 800
rect 60278 0 60334 800
rect 60554 0 60610 800
rect 60830 0 60886 800
rect 61198 0 61254 800
rect 61474 0 61530 800
rect 61750 0 61806 800
rect 62026 0 62082 800
rect 62302 0 62358 800
rect 62670 0 62726 800
rect 62946 0 63002 800
rect 63222 0 63278 800
rect 63498 0 63554 800
rect 63866 0 63922 800
rect 64142 0 64198 800
rect 64418 0 64474 800
rect 64694 0 64750 800
rect 65062 0 65118 800
rect 65338 0 65394 800
rect 65614 0 65670 800
rect 65890 0 65946 800
rect 66258 0 66314 800
rect 66534 0 66590 800
rect 66810 0 66866 800
rect 67086 0 67142 800
rect 67454 0 67510 800
rect 67730 0 67786 800
rect 68006 0 68062 800
rect 68282 0 68338 800
rect 68650 0 68706 800
rect 68926 0 68982 800
rect 69202 0 69258 800
rect 69478 0 69534 800
rect 69754 0 69810 800
rect 70122 0 70178 800
rect 70398 0 70454 800
rect 70674 0 70730 800
rect 70950 0 71006 800
rect 71318 0 71374 800
rect 71594 0 71650 800
rect 71870 0 71926 800
rect 72146 0 72202 800
rect 72514 0 72570 800
rect 72790 0 72846 800
rect 73066 0 73122 800
rect 73342 0 73398 800
rect 73710 0 73766 800
rect 73986 0 74042 800
rect 74262 0 74318 800
rect 74538 0 74594 800
rect 74906 0 74962 800
rect 75182 0 75238 800
rect 75458 0 75514 800
rect 75734 0 75790 800
rect 76010 0 76066 800
rect 76378 0 76434 800
rect 76654 0 76710 800
rect 76930 0 76986 800
rect 77206 0 77262 800
rect 77574 0 77630 800
rect 77850 0 77906 800
rect 78126 0 78182 800
rect 78402 0 78458 800
rect 78770 0 78826 800
rect 79046 0 79102 800
rect 79322 0 79378 800
rect 79598 0 79654 800
rect 79966 0 80022 800
rect 80242 0 80298 800
rect 80518 0 80574 800
rect 80794 0 80850 800
rect 81162 0 81218 800
rect 81438 0 81494 800
rect 81714 0 81770 800
rect 81990 0 82046 800
rect 82358 0 82414 800
rect 82634 0 82690 800
rect 82910 0 82966 800
rect 83186 0 83242 800
rect 83462 0 83518 800
rect 83830 0 83886 800
rect 84106 0 84162 800
rect 84382 0 84438 800
rect 84658 0 84714 800
rect 85026 0 85082 800
rect 85302 0 85358 800
rect 85578 0 85634 800
rect 85854 0 85910 800
rect 86222 0 86278 800
rect 86498 0 86554 800
rect 86774 0 86830 800
rect 87050 0 87106 800
rect 87418 0 87474 800
rect 87694 0 87750 800
rect 87970 0 88026 800
rect 88246 0 88302 800
rect 88614 0 88670 800
rect 88890 0 88946 800
rect 89166 0 89222 800
rect 89442 0 89498 800
rect 89718 0 89774 800
rect 90086 0 90142 800
rect 90362 0 90418 800
rect 90638 0 90694 800
rect 90914 0 90970 800
rect 91282 0 91338 800
rect 91558 0 91614 800
rect 91834 0 91890 800
rect 92110 0 92166 800
rect 92478 0 92534 800
rect 92754 0 92810 800
rect 93030 0 93086 800
rect 93306 0 93362 800
rect 93674 0 93730 800
rect 93950 0 94006 800
rect 94226 0 94282 800
rect 94502 0 94558 800
rect 94870 0 94926 800
rect 95146 0 95202 800
rect 95422 0 95478 800
rect 95698 0 95754 800
rect 96066 0 96122 800
rect 96342 0 96398 800
rect 96618 0 96674 800
rect 96894 0 96950 800
rect 97170 0 97226 800
rect 97538 0 97594 800
rect 97814 0 97870 800
rect 98090 0 98146 800
rect 98366 0 98422 800
rect 98734 0 98790 800
rect 99010 0 99066 800
rect 99286 0 99342 800
rect 99562 0 99618 800
rect 99930 0 99986 800
rect 100206 0 100262 800
rect 100482 0 100538 800
rect 100758 0 100814 800
rect 101126 0 101182 800
rect 101402 0 101458 800
rect 101678 0 101734 800
rect 101954 0 102010 800
rect 102322 0 102378 800
rect 102598 0 102654 800
rect 102874 0 102930 800
rect 103150 0 103206 800
rect 103426 0 103482 800
rect 103794 0 103850 800
rect 104070 0 104126 800
rect 104346 0 104402 800
rect 104622 0 104678 800
rect 104990 0 105046 800
rect 105266 0 105322 800
rect 105542 0 105598 800
rect 105818 0 105874 800
rect 106186 0 106242 800
rect 106462 0 106518 800
rect 106738 0 106794 800
rect 107014 0 107070 800
rect 107382 0 107438 800
rect 107658 0 107714 800
rect 107934 0 107990 800
rect 108210 0 108266 800
rect 108578 0 108634 800
rect 108854 0 108910 800
rect 109130 0 109186 800
rect 109406 0 109462 800
rect 109774 0 109830 800
rect 110050 0 110106 800
rect 110326 0 110382 800
rect 110602 0 110658 800
rect 110878 0 110934 800
rect 111246 0 111302 800
rect 111522 0 111578 800
rect 111798 0 111854 800
rect 112074 0 112130 800
rect 112442 0 112498 800
rect 112718 0 112774 800
rect 112994 0 113050 800
rect 113270 0 113326 800
rect 113638 0 113694 800
rect 113914 0 113970 800
rect 114190 0 114246 800
rect 114466 0 114522 800
rect 114834 0 114890 800
rect 115110 0 115166 800
rect 115386 0 115442 800
rect 115662 0 115718 800
rect 116030 0 116086 800
rect 116306 0 116362 800
rect 116582 0 116638 800
rect 116858 0 116914 800
rect 117134 0 117190 800
rect 117502 0 117558 800
rect 117778 0 117834 800
rect 118054 0 118110 800
rect 118330 0 118386 800
rect 118698 0 118754 800
rect 118974 0 119030 800
rect 119250 0 119306 800
rect 119526 0 119582 800
rect 119894 0 119950 800
rect 120170 0 120226 800
rect 120446 0 120502 800
rect 120722 0 120778 800
rect 121090 0 121146 800
rect 121366 0 121422 800
rect 121642 0 121698 800
rect 121918 0 121974 800
rect 122286 0 122342 800
rect 122562 0 122618 800
rect 122838 0 122894 800
rect 123114 0 123170 800
rect 123482 0 123538 800
rect 123758 0 123814 800
rect 124034 0 124090 800
rect 124310 0 124366 800
rect 124586 0 124642 800
rect 124954 0 125010 800
rect 125230 0 125286 800
rect 125506 0 125562 800
rect 125782 0 125838 800
rect 126150 0 126206 800
rect 126426 0 126482 800
rect 126702 0 126758 800
rect 126978 0 127034 800
rect 127346 0 127402 800
rect 127622 0 127678 800
rect 127898 0 127954 800
rect 128174 0 128230 800
rect 128542 0 128598 800
rect 128818 0 128874 800
rect 129094 0 129150 800
rect 129370 0 129426 800
rect 129738 0 129794 800
rect 130014 0 130070 800
rect 130290 0 130346 800
rect 130566 0 130622 800
rect 130842 0 130898 800
rect 131210 0 131266 800
rect 131486 0 131542 800
rect 131762 0 131818 800
rect 132038 0 132094 800
rect 132406 0 132462 800
rect 132682 0 132738 800
rect 132958 0 133014 800
rect 133234 0 133290 800
rect 133602 0 133658 800
rect 133878 0 133934 800
rect 134154 0 134210 800
rect 134430 0 134486 800
rect 134798 0 134854 800
rect 135074 0 135130 800
rect 135350 0 135406 800
rect 135626 0 135682 800
rect 135994 0 136050 800
rect 136270 0 136326 800
rect 136546 0 136602 800
rect 136822 0 136878 800
rect 137190 0 137246 800
rect 137466 0 137522 800
rect 137742 0 137798 800
rect 138018 0 138074 800
rect 138294 0 138350 800
rect 138662 0 138718 800
rect 138938 0 138994 800
rect 139214 0 139270 800
rect 139490 0 139546 800
rect 139858 0 139914 800
rect 140134 0 140190 800
rect 140410 0 140466 800
rect 140686 0 140742 800
rect 141054 0 141110 800
rect 141330 0 141386 800
rect 141606 0 141662 800
rect 141882 0 141938 800
rect 142250 0 142306 800
rect 142526 0 142582 800
rect 142802 0 142858 800
rect 143078 0 143134 800
rect 143446 0 143502 800
rect 143722 0 143778 800
rect 143998 0 144054 800
rect 144274 0 144330 800
rect 144550 0 144606 800
rect 144918 0 144974 800
rect 145194 0 145250 800
rect 145470 0 145526 800
rect 145746 0 145802 800
rect 146114 0 146170 800
rect 146390 0 146446 800
rect 146666 0 146722 800
rect 146942 0 146998 800
rect 147310 0 147366 800
rect 147586 0 147642 800
rect 147862 0 147918 800
rect 148138 0 148194 800
rect 148506 0 148562 800
rect 148782 0 148838 800
rect 149058 0 149114 800
rect 149334 0 149390 800
rect 149702 0 149758 800
rect 149978 0 150034 800
rect 150254 0 150310 800
rect 150530 0 150586 800
rect 150898 0 150954 800
rect 151174 0 151230 800
rect 151450 0 151506 800
rect 151726 0 151782 800
rect 152002 0 152058 800
rect 152370 0 152426 800
rect 152646 0 152702 800
rect 152922 0 152978 800
rect 153198 0 153254 800
rect 153566 0 153622 800
rect 153842 0 153898 800
rect 154118 0 154174 800
rect 154394 0 154450 800
rect 154762 0 154818 800
rect 155038 0 155094 800
rect 155314 0 155370 800
rect 155590 0 155646 800
rect 155958 0 156014 800
rect 156234 0 156290 800
rect 156510 0 156566 800
rect 156786 0 156842 800
rect 157154 0 157210 800
rect 157430 0 157486 800
rect 157706 0 157762 800
rect 157982 0 158038 800
rect 158258 0 158314 800
rect 158626 0 158682 800
rect 158902 0 158958 800
rect 159178 0 159234 800
rect 159454 0 159510 800
rect 159822 0 159878 800
rect 160098 0 160154 800
rect 160374 0 160430 800
rect 160650 0 160706 800
rect 161018 0 161074 800
rect 161294 0 161350 800
rect 161570 0 161626 800
rect 161846 0 161902 800
rect 162214 0 162270 800
rect 162490 0 162546 800
rect 162766 0 162822 800
rect 163042 0 163098 800
rect 163410 0 163466 800
rect 163686 0 163742 800
rect 163962 0 164018 800
rect 164238 0 164294 800
<< obsm2 >>
rect 112 165819 422 165875
rect 590 165819 1342 165875
rect 1510 165819 2262 165875
rect 2430 165819 3274 165875
rect 3442 165819 4194 165875
rect 4362 165819 5114 165875
rect 5282 165819 6126 165875
rect 6294 165819 7046 165875
rect 7214 165819 7966 165875
rect 8134 165819 8978 165875
rect 9146 165819 9898 165875
rect 10066 165819 10818 165875
rect 10986 165819 11830 165875
rect 11998 165819 12750 165875
rect 12918 165819 13670 165875
rect 13838 165819 14682 165875
rect 14850 165819 15602 165875
rect 15770 165819 16522 165875
rect 16690 165819 17534 165875
rect 17702 165819 18454 165875
rect 18622 165819 19374 165875
rect 19542 165819 20386 165875
rect 20554 165819 21306 165875
rect 21474 165819 22226 165875
rect 22394 165819 23238 165875
rect 23406 165819 24158 165875
rect 24326 165819 25078 165875
rect 25246 165819 26090 165875
rect 26258 165819 27010 165875
rect 27178 165819 27930 165875
rect 28098 165819 28942 165875
rect 29110 165819 29862 165875
rect 30030 165819 30782 165875
rect 30950 165819 31794 165875
rect 31962 165819 32714 165875
rect 32882 165819 33634 165875
rect 33802 165819 34646 165875
rect 34814 165819 35566 165875
rect 35734 165819 36486 165875
rect 36654 165819 37498 165875
rect 37666 165819 38418 165875
rect 38586 165819 39338 165875
rect 39506 165819 40350 165875
rect 40518 165819 41270 165875
rect 41438 165819 42190 165875
rect 42358 165819 43202 165875
rect 43370 165819 44122 165875
rect 44290 165819 45042 165875
rect 45210 165819 46054 165875
rect 46222 165819 46974 165875
rect 47142 165819 47894 165875
rect 48062 165819 48906 165875
rect 49074 165819 49826 165875
rect 49994 165819 50746 165875
rect 50914 165819 51758 165875
rect 51926 165819 52678 165875
rect 52846 165819 53598 165875
rect 53766 165819 54610 165875
rect 54778 165819 55530 165875
rect 55698 165819 56450 165875
rect 56618 165819 57462 165875
rect 57630 165819 58382 165875
rect 58550 165819 59302 165875
rect 59470 165819 60314 165875
rect 60482 165819 61234 165875
rect 61402 165819 62154 165875
rect 62322 165819 63166 165875
rect 63334 165819 64086 165875
rect 64254 165819 65006 165875
rect 65174 165819 66018 165875
rect 66186 165819 66938 165875
rect 67106 165819 67858 165875
rect 68026 165819 68870 165875
rect 69038 165819 69790 165875
rect 69958 165819 70710 165875
rect 70878 165819 71722 165875
rect 71890 165819 72642 165875
rect 72810 165819 73562 165875
rect 73730 165819 74574 165875
rect 74742 165819 75494 165875
rect 75662 165819 76414 165875
rect 76582 165819 77426 165875
rect 77594 165819 78346 165875
rect 78514 165819 79266 165875
rect 79434 165819 80278 165875
rect 80446 165819 81198 165875
rect 81366 165819 82118 165875
rect 82286 165819 83130 165875
rect 83298 165819 84050 165875
rect 84218 165819 84970 165875
rect 85138 165819 85982 165875
rect 86150 165819 86902 165875
rect 87070 165819 87822 165875
rect 87990 165819 88834 165875
rect 89002 165819 89754 165875
rect 89922 165819 90674 165875
rect 90842 165819 91686 165875
rect 91854 165819 92606 165875
rect 92774 165819 93526 165875
rect 93694 165819 94538 165875
rect 94706 165819 95458 165875
rect 95626 165819 96378 165875
rect 96546 165819 97390 165875
rect 97558 165819 98310 165875
rect 98478 165819 99230 165875
rect 99398 165819 100242 165875
rect 100410 165819 101162 165875
rect 101330 165819 102082 165875
rect 102250 165819 103094 165875
rect 103262 165819 104014 165875
rect 104182 165819 104934 165875
rect 105102 165819 105946 165875
rect 106114 165819 106866 165875
rect 107034 165819 107786 165875
rect 107954 165819 108798 165875
rect 108966 165819 109718 165875
rect 109886 165819 110638 165875
rect 110806 165819 111650 165875
rect 111818 165819 112570 165875
rect 112738 165819 113490 165875
rect 113658 165819 114502 165875
rect 114670 165819 115422 165875
rect 115590 165819 116342 165875
rect 116510 165819 117354 165875
rect 117522 165819 118274 165875
rect 118442 165819 119194 165875
rect 119362 165819 120206 165875
rect 120374 165819 121126 165875
rect 121294 165819 122046 165875
rect 122214 165819 123058 165875
rect 123226 165819 123978 165875
rect 124146 165819 124898 165875
rect 125066 165819 125910 165875
rect 126078 165819 126830 165875
rect 126998 165819 127750 165875
rect 127918 165819 128762 165875
rect 128930 165819 129682 165875
rect 129850 165819 130602 165875
rect 130770 165819 131614 165875
rect 131782 165819 132534 165875
rect 132702 165819 133454 165875
rect 133622 165819 134466 165875
rect 134634 165819 135386 165875
rect 135554 165819 136306 165875
rect 136474 165819 137318 165875
rect 137486 165819 138238 165875
rect 138406 165819 139158 165875
rect 139326 165819 140170 165875
rect 140338 165819 141090 165875
rect 141258 165819 142010 165875
rect 142178 165819 143022 165875
rect 143190 165819 143942 165875
rect 144110 165819 144862 165875
rect 145030 165819 145874 165875
rect 146042 165819 146794 165875
rect 146962 165819 147714 165875
rect 147882 165819 148726 165875
rect 148894 165819 149646 165875
rect 149814 165819 150566 165875
rect 150734 165819 151578 165875
rect 151746 165819 152498 165875
rect 152666 165819 153418 165875
rect 153586 165819 154430 165875
rect 154598 165819 155350 165875
rect 155518 165819 156270 165875
rect 156438 165819 157282 165875
rect 157450 165819 158202 165875
rect 158370 165819 159122 165875
rect 159290 165819 160134 165875
rect 160302 165819 161054 165875
rect 161222 165819 161974 165875
rect 162142 165819 162986 165875
rect 163154 165819 163906 165875
rect 164074 165819 164478 165875
rect 112 856 164478 165819
rect 222 478 330 856
rect 498 478 606 856
rect 774 478 882 856
rect 1050 478 1158 856
rect 1326 478 1526 856
rect 1694 478 1802 856
rect 1970 478 2078 856
rect 2246 478 2354 856
rect 2522 478 2722 856
rect 2890 478 2998 856
rect 3166 478 3274 856
rect 3442 478 3550 856
rect 3718 478 3918 856
rect 4086 478 4194 856
rect 4362 478 4470 856
rect 4638 478 4746 856
rect 4914 478 5114 856
rect 5282 478 5390 856
rect 5558 478 5666 856
rect 5834 478 5942 856
rect 6110 478 6310 856
rect 6478 478 6586 856
rect 6754 478 6862 856
rect 7030 478 7138 856
rect 7306 478 7414 856
rect 7582 478 7782 856
rect 7950 478 8058 856
rect 8226 478 8334 856
rect 8502 478 8610 856
rect 8778 478 8978 856
rect 9146 478 9254 856
rect 9422 478 9530 856
rect 9698 478 9806 856
rect 9974 478 10174 856
rect 10342 478 10450 856
rect 10618 478 10726 856
rect 10894 478 11002 856
rect 11170 478 11370 856
rect 11538 478 11646 856
rect 11814 478 11922 856
rect 12090 478 12198 856
rect 12366 478 12566 856
rect 12734 478 12842 856
rect 13010 478 13118 856
rect 13286 478 13394 856
rect 13562 478 13762 856
rect 13930 478 14038 856
rect 14206 478 14314 856
rect 14482 478 14590 856
rect 14758 478 14866 856
rect 15034 478 15234 856
rect 15402 478 15510 856
rect 15678 478 15786 856
rect 15954 478 16062 856
rect 16230 478 16430 856
rect 16598 478 16706 856
rect 16874 478 16982 856
rect 17150 478 17258 856
rect 17426 478 17626 856
rect 17794 478 17902 856
rect 18070 478 18178 856
rect 18346 478 18454 856
rect 18622 478 18822 856
rect 18990 478 19098 856
rect 19266 478 19374 856
rect 19542 478 19650 856
rect 19818 478 20018 856
rect 20186 478 20294 856
rect 20462 478 20570 856
rect 20738 478 20846 856
rect 21014 478 21122 856
rect 21290 478 21490 856
rect 21658 478 21766 856
rect 21934 478 22042 856
rect 22210 478 22318 856
rect 22486 478 22686 856
rect 22854 478 22962 856
rect 23130 478 23238 856
rect 23406 478 23514 856
rect 23682 478 23882 856
rect 24050 478 24158 856
rect 24326 478 24434 856
rect 24602 478 24710 856
rect 24878 478 25078 856
rect 25246 478 25354 856
rect 25522 478 25630 856
rect 25798 478 25906 856
rect 26074 478 26274 856
rect 26442 478 26550 856
rect 26718 478 26826 856
rect 26994 478 27102 856
rect 27270 478 27470 856
rect 27638 478 27746 856
rect 27914 478 28022 856
rect 28190 478 28298 856
rect 28466 478 28574 856
rect 28742 478 28942 856
rect 29110 478 29218 856
rect 29386 478 29494 856
rect 29662 478 29770 856
rect 29938 478 30138 856
rect 30306 478 30414 856
rect 30582 478 30690 856
rect 30858 478 30966 856
rect 31134 478 31334 856
rect 31502 478 31610 856
rect 31778 478 31886 856
rect 32054 478 32162 856
rect 32330 478 32530 856
rect 32698 478 32806 856
rect 32974 478 33082 856
rect 33250 478 33358 856
rect 33526 478 33726 856
rect 33894 478 34002 856
rect 34170 478 34278 856
rect 34446 478 34554 856
rect 34722 478 34830 856
rect 34998 478 35198 856
rect 35366 478 35474 856
rect 35642 478 35750 856
rect 35918 478 36026 856
rect 36194 478 36394 856
rect 36562 478 36670 856
rect 36838 478 36946 856
rect 37114 478 37222 856
rect 37390 478 37590 856
rect 37758 478 37866 856
rect 38034 478 38142 856
rect 38310 478 38418 856
rect 38586 478 38786 856
rect 38954 478 39062 856
rect 39230 478 39338 856
rect 39506 478 39614 856
rect 39782 478 39982 856
rect 40150 478 40258 856
rect 40426 478 40534 856
rect 40702 478 40810 856
rect 40978 478 41178 856
rect 41346 478 41454 856
rect 41622 478 41730 856
rect 41898 478 42006 856
rect 42174 478 42282 856
rect 42450 478 42650 856
rect 42818 478 42926 856
rect 43094 478 43202 856
rect 43370 478 43478 856
rect 43646 478 43846 856
rect 44014 478 44122 856
rect 44290 478 44398 856
rect 44566 478 44674 856
rect 44842 478 45042 856
rect 45210 478 45318 856
rect 45486 478 45594 856
rect 45762 478 45870 856
rect 46038 478 46238 856
rect 46406 478 46514 856
rect 46682 478 46790 856
rect 46958 478 47066 856
rect 47234 478 47434 856
rect 47602 478 47710 856
rect 47878 478 47986 856
rect 48154 478 48262 856
rect 48430 478 48538 856
rect 48706 478 48906 856
rect 49074 478 49182 856
rect 49350 478 49458 856
rect 49626 478 49734 856
rect 49902 478 50102 856
rect 50270 478 50378 856
rect 50546 478 50654 856
rect 50822 478 50930 856
rect 51098 478 51298 856
rect 51466 478 51574 856
rect 51742 478 51850 856
rect 52018 478 52126 856
rect 52294 478 52494 856
rect 52662 478 52770 856
rect 52938 478 53046 856
rect 53214 478 53322 856
rect 53490 478 53690 856
rect 53858 478 53966 856
rect 54134 478 54242 856
rect 54410 478 54518 856
rect 54686 478 54886 856
rect 55054 478 55162 856
rect 55330 478 55438 856
rect 55606 478 55714 856
rect 55882 478 55990 856
rect 56158 478 56358 856
rect 56526 478 56634 856
rect 56802 478 56910 856
rect 57078 478 57186 856
rect 57354 478 57554 856
rect 57722 478 57830 856
rect 57998 478 58106 856
rect 58274 478 58382 856
rect 58550 478 58750 856
rect 58918 478 59026 856
rect 59194 478 59302 856
rect 59470 478 59578 856
rect 59746 478 59946 856
rect 60114 478 60222 856
rect 60390 478 60498 856
rect 60666 478 60774 856
rect 60942 478 61142 856
rect 61310 478 61418 856
rect 61586 478 61694 856
rect 61862 478 61970 856
rect 62138 478 62246 856
rect 62414 478 62614 856
rect 62782 478 62890 856
rect 63058 478 63166 856
rect 63334 478 63442 856
rect 63610 478 63810 856
rect 63978 478 64086 856
rect 64254 478 64362 856
rect 64530 478 64638 856
rect 64806 478 65006 856
rect 65174 478 65282 856
rect 65450 478 65558 856
rect 65726 478 65834 856
rect 66002 478 66202 856
rect 66370 478 66478 856
rect 66646 478 66754 856
rect 66922 478 67030 856
rect 67198 478 67398 856
rect 67566 478 67674 856
rect 67842 478 67950 856
rect 68118 478 68226 856
rect 68394 478 68594 856
rect 68762 478 68870 856
rect 69038 478 69146 856
rect 69314 478 69422 856
rect 69590 478 69698 856
rect 69866 478 70066 856
rect 70234 478 70342 856
rect 70510 478 70618 856
rect 70786 478 70894 856
rect 71062 478 71262 856
rect 71430 478 71538 856
rect 71706 478 71814 856
rect 71982 478 72090 856
rect 72258 478 72458 856
rect 72626 478 72734 856
rect 72902 478 73010 856
rect 73178 478 73286 856
rect 73454 478 73654 856
rect 73822 478 73930 856
rect 74098 478 74206 856
rect 74374 478 74482 856
rect 74650 478 74850 856
rect 75018 478 75126 856
rect 75294 478 75402 856
rect 75570 478 75678 856
rect 75846 478 75954 856
rect 76122 478 76322 856
rect 76490 478 76598 856
rect 76766 478 76874 856
rect 77042 478 77150 856
rect 77318 478 77518 856
rect 77686 478 77794 856
rect 77962 478 78070 856
rect 78238 478 78346 856
rect 78514 478 78714 856
rect 78882 478 78990 856
rect 79158 478 79266 856
rect 79434 478 79542 856
rect 79710 478 79910 856
rect 80078 478 80186 856
rect 80354 478 80462 856
rect 80630 478 80738 856
rect 80906 478 81106 856
rect 81274 478 81382 856
rect 81550 478 81658 856
rect 81826 478 81934 856
rect 82102 478 82302 856
rect 82470 478 82578 856
rect 82746 478 82854 856
rect 83022 478 83130 856
rect 83298 478 83406 856
rect 83574 478 83774 856
rect 83942 478 84050 856
rect 84218 478 84326 856
rect 84494 478 84602 856
rect 84770 478 84970 856
rect 85138 478 85246 856
rect 85414 478 85522 856
rect 85690 478 85798 856
rect 85966 478 86166 856
rect 86334 478 86442 856
rect 86610 478 86718 856
rect 86886 478 86994 856
rect 87162 478 87362 856
rect 87530 478 87638 856
rect 87806 478 87914 856
rect 88082 478 88190 856
rect 88358 478 88558 856
rect 88726 478 88834 856
rect 89002 478 89110 856
rect 89278 478 89386 856
rect 89554 478 89662 856
rect 89830 478 90030 856
rect 90198 478 90306 856
rect 90474 478 90582 856
rect 90750 478 90858 856
rect 91026 478 91226 856
rect 91394 478 91502 856
rect 91670 478 91778 856
rect 91946 478 92054 856
rect 92222 478 92422 856
rect 92590 478 92698 856
rect 92866 478 92974 856
rect 93142 478 93250 856
rect 93418 478 93618 856
rect 93786 478 93894 856
rect 94062 478 94170 856
rect 94338 478 94446 856
rect 94614 478 94814 856
rect 94982 478 95090 856
rect 95258 478 95366 856
rect 95534 478 95642 856
rect 95810 478 96010 856
rect 96178 478 96286 856
rect 96454 478 96562 856
rect 96730 478 96838 856
rect 97006 478 97114 856
rect 97282 478 97482 856
rect 97650 478 97758 856
rect 97926 478 98034 856
rect 98202 478 98310 856
rect 98478 478 98678 856
rect 98846 478 98954 856
rect 99122 478 99230 856
rect 99398 478 99506 856
rect 99674 478 99874 856
rect 100042 478 100150 856
rect 100318 478 100426 856
rect 100594 478 100702 856
rect 100870 478 101070 856
rect 101238 478 101346 856
rect 101514 478 101622 856
rect 101790 478 101898 856
rect 102066 478 102266 856
rect 102434 478 102542 856
rect 102710 478 102818 856
rect 102986 478 103094 856
rect 103262 478 103370 856
rect 103538 478 103738 856
rect 103906 478 104014 856
rect 104182 478 104290 856
rect 104458 478 104566 856
rect 104734 478 104934 856
rect 105102 478 105210 856
rect 105378 478 105486 856
rect 105654 478 105762 856
rect 105930 478 106130 856
rect 106298 478 106406 856
rect 106574 478 106682 856
rect 106850 478 106958 856
rect 107126 478 107326 856
rect 107494 478 107602 856
rect 107770 478 107878 856
rect 108046 478 108154 856
rect 108322 478 108522 856
rect 108690 478 108798 856
rect 108966 478 109074 856
rect 109242 478 109350 856
rect 109518 478 109718 856
rect 109886 478 109994 856
rect 110162 478 110270 856
rect 110438 478 110546 856
rect 110714 478 110822 856
rect 110990 478 111190 856
rect 111358 478 111466 856
rect 111634 478 111742 856
rect 111910 478 112018 856
rect 112186 478 112386 856
rect 112554 478 112662 856
rect 112830 478 112938 856
rect 113106 478 113214 856
rect 113382 478 113582 856
rect 113750 478 113858 856
rect 114026 478 114134 856
rect 114302 478 114410 856
rect 114578 478 114778 856
rect 114946 478 115054 856
rect 115222 478 115330 856
rect 115498 478 115606 856
rect 115774 478 115974 856
rect 116142 478 116250 856
rect 116418 478 116526 856
rect 116694 478 116802 856
rect 116970 478 117078 856
rect 117246 478 117446 856
rect 117614 478 117722 856
rect 117890 478 117998 856
rect 118166 478 118274 856
rect 118442 478 118642 856
rect 118810 478 118918 856
rect 119086 478 119194 856
rect 119362 478 119470 856
rect 119638 478 119838 856
rect 120006 478 120114 856
rect 120282 478 120390 856
rect 120558 478 120666 856
rect 120834 478 121034 856
rect 121202 478 121310 856
rect 121478 478 121586 856
rect 121754 478 121862 856
rect 122030 478 122230 856
rect 122398 478 122506 856
rect 122674 478 122782 856
rect 122950 478 123058 856
rect 123226 478 123426 856
rect 123594 478 123702 856
rect 123870 478 123978 856
rect 124146 478 124254 856
rect 124422 478 124530 856
rect 124698 478 124898 856
rect 125066 478 125174 856
rect 125342 478 125450 856
rect 125618 478 125726 856
rect 125894 478 126094 856
rect 126262 478 126370 856
rect 126538 478 126646 856
rect 126814 478 126922 856
rect 127090 478 127290 856
rect 127458 478 127566 856
rect 127734 478 127842 856
rect 128010 478 128118 856
rect 128286 478 128486 856
rect 128654 478 128762 856
rect 128930 478 129038 856
rect 129206 478 129314 856
rect 129482 478 129682 856
rect 129850 478 129958 856
rect 130126 478 130234 856
rect 130402 478 130510 856
rect 130678 478 130786 856
rect 130954 478 131154 856
rect 131322 478 131430 856
rect 131598 478 131706 856
rect 131874 478 131982 856
rect 132150 478 132350 856
rect 132518 478 132626 856
rect 132794 478 132902 856
rect 133070 478 133178 856
rect 133346 478 133546 856
rect 133714 478 133822 856
rect 133990 478 134098 856
rect 134266 478 134374 856
rect 134542 478 134742 856
rect 134910 478 135018 856
rect 135186 478 135294 856
rect 135462 478 135570 856
rect 135738 478 135938 856
rect 136106 478 136214 856
rect 136382 478 136490 856
rect 136658 478 136766 856
rect 136934 478 137134 856
rect 137302 478 137410 856
rect 137578 478 137686 856
rect 137854 478 137962 856
rect 138130 478 138238 856
rect 138406 478 138606 856
rect 138774 478 138882 856
rect 139050 478 139158 856
rect 139326 478 139434 856
rect 139602 478 139802 856
rect 139970 478 140078 856
rect 140246 478 140354 856
rect 140522 478 140630 856
rect 140798 478 140998 856
rect 141166 478 141274 856
rect 141442 478 141550 856
rect 141718 478 141826 856
rect 141994 478 142194 856
rect 142362 478 142470 856
rect 142638 478 142746 856
rect 142914 478 143022 856
rect 143190 478 143390 856
rect 143558 478 143666 856
rect 143834 478 143942 856
rect 144110 478 144218 856
rect 144386 478 144494 856
rect 144662 478 144862 856
rect 145030 478 145138 856
rect 145306 478 145414 856
rect 145582 478 145690 856
rect 145858 478 146058 856
rect 146226 478 146334 856
rect 146502 478 146610 856
rect 146778 478 146886 856
rect 147054 478 147254 856
rect 147422 478 147530 856
rect 147698 478 147806 856
rect 147974 478 148082 856
rect 148250 478 148450 856
rect 148618 478 148726 856
rect 148894 478 149002 856
rect 149170 478 149278 856
rect 149446 478 149646 856
rect 149814 478 149922 856
rect 150090 478 150198 856
rect 150366 478 150474 856
rect 150642 478 150842 856
rect 151010 478 151118 856
rect 151286 478 151394 856
rect 151562 478 151670 856
rect 151838 478 151946 856
rect 152114 478 152314 856
rect 152482 478 152590 856
rect 152758 478 152866 856
rect 153034 478 153142 856
rect 153310 478 153510 856
rect 153678 478 153786 856
rect 153954 478 154062 856
rect 154230 478 154338 856
rect 154506 478 154706 856
rect 154874 478 154982 856
rect 155150 478 155258 856
rect 155426 478 155534 856
rect 155702 478 155902 856
rect 156070 478 156178 856
rect 156346 478 156454 856
rect 156622 478 156730 856
rect 156898 478 157098 856
rect 157266 478 157374 856
rect 157542 478 157650 856
rect 157818 478 157926 856
rect 158094 478 158202 856
rect 158370 478 158570 856
rect 158738 478 158846 856
rect 159014 478 159122 856
rect 159290 478 159398 856
rect 159566 478 159766 856
rect 159934 478 160042 856
rect 160210 478 160318 856
rect 160486 478 160594 856
rect 160762 478 160962 856
rect 161130 478 161238 856
rect 161406 478 161514 856
rect 161682 478 161790 856
rect 161958 478 162158 856
rect 162326 478 162434 856
rect 162602 478 162710 856
rect 162878 478 162986 856
rect 163154 478 163354 856
rect 163522 478 163630 856
rect 163798 478 163906 856
rect 164074 478 164182 856
rect 164350 478 164478 856
<< metal3 >>
rect 0 165248 800 165368
rect 163731 165248 164531 165368
rect 0 162528 800 162648
rect 163731 162528 164531 162648
rect 0 159808 800 159928
rect 163731 159808 164531 159928
rect 0 157088 800 157208
rect 163731 157088 164531 157208
rect 0 154504 800 154624
rect 163731 154504 164531 154624
rect 0 151784 800 151904
rect 163731 151784 164531 151904
rect 0 149064 800 149184
rect 163731 149064 164531 149184
rect 0 146344 800 146464
rect 163731 146344 164531 146464
rect 0 143760 800 143880
rect 163731 143760 164531 143880
rect 0 141040 800 141160
rect 163731 141040 164531 141160
rect 0 138320 800 138440
rect 163731 138320 164531 138440
rect 0 135600 800 135720
rect 163731 135600 164531 135720
rect 0 132880 800 133000
rect 163731 132880 164531 133000
rect 0 130296 800 130416
rect 163731 130296 164531 130416
rect 0 127576 800 127696
rect 163731 127576 164531 127696
rect 0 124856 800 124976
rect 163731 124856 164531 124976
rect 0 122136 800 122256
rect 163731 122136 164531 122256
rect 0 119552 800 119672
rect 163731 119552 164531 119672
rect 0 116832 800 116952
rect 163731 116832 164531 116952
rect 0 114112 800 114232
rect 163731 114112 164531 114232
rect 0 111392 800 111512
rect 163731 111392 164531 111512
rect 0 108672 800 108792
rect 163731 108672 164531 108792
rect 0 106088 800 106208
rect 163731 106088 164531 106208
rect 0 103368 800 103488
rect 163731 103368 164531 103488
rect 0 100648 800 100768
rect 163731 100648 164531 100768
rect 0 97928 800 98048
rect 163731 97928 164531 98048
rect 0 95344 800 95464
rect 163731 95344 164531 95464
rect 0 92624 800 92744
rect 163731 92624 164531 92744
rect 0 89904 800 90024
rect 163731 89904 164531 90024
rect 0 87184 800 87304
rect 163731 87184 164531 87304
rect 0 84600 800 84720
rect 163731 84600 164531 84720
rect 0 81880 800 82000
rect 163731 81880 164531 82000
rect 0 79160 800 79280
rect 163731 79160 164531 79280
rect 0 76440 800 76560
rect 163731 76440 164531 76560
rect 0 73720 800 73840
rect 163731 73720 164531 73840
rect 0 71136 800 71256
rect 163731 71136 164531 71256
rect 0 68416 800 68536
rect 163731 68416 164531 68536
rect 0 65696 800 65816
rect 163731 65696 164531 65816
rect 0 62976 800 63096
rect 163731 62976 164531 63096
rect 0 60392 800 60512
rect 163731 60392 164531 60512
rect 0 57672 800 57792
rect 163731 57672 164531 57792
rect 0 54952 800 55072
rect 163731 54952 164531 55072
rect 0 52232 800 52352
rect 163731 52232 164531 52352
rect 0 49512 800 49632
rect 163731 49512 164531 49632
rect 0 46928 800 47048
rect 163731 46928 164531 47048
rect 0 44208 800 44328
rect 163731 44208 164531 44328
rect 0 41488 800 41608
rect 163731 41488 164531 41608
rect 0 38768 800 38888
rect 163731 38768 164531 38888
rect 0 36184 800 36304
rect 163731 36184 164531 36304
rect 0 33464 800 33584
rect 163731 33464 164531 33584
rect 0 30744 800 30864
rect 163731 30744 164531 30864
rect 0 28024 800 28144
rect 163731 28024 164531 28144
rect 0 25304 800 25424
rect 163731 25304 164531 25424
rect 0 22720 800 22840
rect 163731 22720 164531 22840
rect 0 20000 800 20120
rect 163731 20000 164531 20120
rect 0 17280 800 17400
rect 163731 17280 164531 17400
rect 0 14560 800 14680
rect 163731 14560 164531 14680
rect 0 11976 800 12096
rect 163731 11976 164531 12096
rect 0 9256 800 9376
rect 163731 9256 164531 9376
rect 0 6536 800 6656
rect 163731 6536 164531 6656
rect 0 3816 800 3936
rect 163731 3816 164531 3936
rect 0 1232 800 1352
rect 163731 1232 164531 1352
<< obsm3 >>
rect 880 165168 163651 165341
rect 800 162728 164483 165168
rect 880 162448 163651 162728
rect 800 160008 164483 162448
rect 880 159728 163651 160008
rect 800 157288 164483 159728
rect 880 157008 163651 157288
rect 800 154704 164483 157008
rect 880 154424 163651 154704
rect 800 151984 164483 154424
rect 880 151704 163651 151984
rect 800 149264 164483 151704
rect 880 148984 163651 149264
rect 800 146544 164483 148984
rect 880 146264 163651 146544
rect 800 143960 164483 146264
rect 880 143680 163651 143960
rect 800 141240 164483 143680
rect 880 140960 163651 141240
rect 800 138520 164483 140960
rect 880 138240 163651 138520
rect 800 135800 164483 138240
rect 880 135520 163651 135800
rect 800 133080 164483 135520
rect 880 132800 163651 133080
rect 800 130496 164483 132800
rect 880 130216 163651 130496
rect 800 127776 164483 130216
rect 880 127496 163651 127776
rect 800 125056 164483 127496
rect 880 124776 163651 125056
rect 800 122336 164483 124776
rect 880 122056 163651 122336
rect 800 119752 164483 122056
rect 880 119472 163651 119752
rect 800 117032 164483 119472
rect 880 116752 163651 117032
rect 800 114312 164483 116752
rect 880 114032 163651 114312
rect 800 111592 164483 114032
rect 880 111312 163651 111592
rect 800 108872 164483 111312
rect 880 108592 163651 108872
rect 800 106288 164483 108592
rect 880 106008 163651 106288
rect 800 103568 164483 106008
rect 880 103288 163651 103568
rect 800 100848 164483 103288
rect 880 100568 163651 100848
rect 800 98128 164483 100568
rect 880 97848 163651 98128
rect 800 95544 164483 97848
rect 880 95264 163651 95544
rect 800 92824 164483 95264
rect 880 92544 163651 92824
rect 800 90104 164483 92544
rect 880 89824 163651 90104
rect 800 87384 164483 89824
rect 880 87104 163651 87384
rect 800 84800 164483 87104
rect 880 84520 163651 84800
rect 800 82080 164483 84520
rect 880 81800 163651 82080
rect 800 79360 164483 81800
rect 880 79080 163651 79360
rect 800 76640 164483 79080
rect 880 76360 163651 76640
rect 800 73920 164483 76360
rect 880 73640 163651 73920
rect 800 71336 164483 73640
rect 880 71056 163651 71336
rect 800 68616 164483 71056
rect 880 68336 163651 68616
rect 800 65896 164483 68336
rect 880 65616 163651 65896
rect 800 63176 164483 65616
rect 880 62896 163651 63176
rect 800 60592 164483 62896
rect 880 60312 163651 60592
rect 800 57872 164483 60312
rect 880 57592 163651 57872
rect 800 55152 164483 57592
rect 880 54872 163651 55152
rect 800 52432 164483 54872
rect 880 52152 163651 52432
rect 800 49712 164483 52152
rect 880 49432 163651 49712
rect 800 47128 164483 49432
rect 880 46848 163651 47128
rect 800 44408 164483 46848
rect 880 44128 163651 44408
rect 800 41688 164483 44128
rect 880 41408 163651 41688
rect 800 38968 164483 41408
rect 880 38688 163651 38968
rect 800 36384 164483 38688
rect 880 36104 163651 36384
rect 800 33664 164483 36104
rect 880 33384 163651 33664
rect 800 30944 164483 33384
rect 880 30664 163651 30944
rect 800 28224 164483 30664
rect 880 27944 163651 28224
rect 800 25504 164483 27944
rect 880 25224 163651 25504
rect 800 22920 164483 25224
rect 880 22640 163651 22920
rect 800 20200 164483 22640
rect 880 19920 163651 20200
rect 800 17480 164483 19920
rect 880 17200 163651 17480
rect 800 14760 164483 17200
rect 880 14480 163651 14760
rect 800 12176 164483 14480
rect 880 11896 163651 12176
rect 800 9456 164483 11896
rect 880 9176 163651 9456
rect 800 6736 164483 9176
rect 880 6456 163651 6736
rect 800 4016 164483 6456
rect 880 3736 163651 4016
rect 800 1432 164483 3736
rect 880 1152 163651 1432
rect 800 444 164483 1152
<< metal4 >>
rect 4208 2128 4528 164336
rect 19568 2128 19888 164336
rect 34928 2128 35248 164336
rect 50288 2128 50608 164336
rect 65648 2128 65968 164336
rect 81008 2128 81328 164336
rect 96368 2128 96688 164336
rect 111728 2128 112048 164336
rect 127088 2128 127408 164336
rect 142448 2128 142768 164336
rect 157808 2128 158128 164336
<< obsm4 >>
rect 5027 2048 19488 164117
rect 19968 2048 34848 164117
rect 35328 2048 50208 164117
rect 50688 2048 65568 164117
rect 66048 2048 80928 164117
rect 81408 2048 96288 164117
rect 96768 2048 111648 164117
rect 112128 2048 127008 164117
rect 127488 2048 142368 164117
rect 142848 2048 157728 164117
rect 158208 2048 164253 164117
rect 5027 443 164253 2048
<< labels >>
rlabel metal3 s 0 6536 800 6656 6 i_dout0[0]
port 1 nsew signal input
rlabel metal2 s 134522 165875 134578 166675 6 i_dout0[10]
port 2 nsew signal input
rlabel metal3 s 163731 81880 164531 82000 6 i_dout0[11]
port 3 nsew signal input
rlabel metal2 s 137374 165875 137430 166675 6 i_dout0[12]
port 4 nsew signal input
rlabel metal3 s 0 79160 800 79280 6 i_dout0[13]
port 5 nsew signal input
rlabel metal3 s 0 81880 800 82000 6 i_dout0[14]
port 6 nsew signal input
rlabel metal3 s 163731 100648 164531 100768 6 i_dout0[15]
port 7 nsew signal input
rlabel metal2 s 157430 0 157486 800 6 i_dout0[16]
port 8 nsew signal input
rlabel metal3 s 0 100648 800 100768 6 i_dout0[17]
port 9 nsew signal input
rlabel metal2 s 157982 0 158038 800 6 i_dout0[18]
port 10 nsew signal input
rlabel metal2 s 158902 0 158958 800 6 i_dout0[19]
port 11 nsew signal input
rlabel metal3 s 163731 14560 164531 14680 6 i_dout0[1]
port 12 nsew signal input
rlabel metal3 s 0 111392 800 111512 6 i_dout0[20]
port 13 nsew signal input
rlabel metal3 s 0 116832 800 116952 6 i_dout0[21]
port 14 nsew signal input
rlabel metal2 s 160374 0 160430 800 6 i_dout0[22]
port 15 nsew signal input
rlabel metal2 s 150622 165875 150678 166675 6 i_dout0[23]
port 16 nsew signal input
rlabel metal3 s 0 130296 800 130416 6 i_dout0[24]
port 17 nsew signal input
rlabel metal2 s 153474 165875 153530 166675 6 i_dout0[25]
port 18 nsew signal input
rlabel metal3 s 163731 146344 164531 146464 6 i_dout0[26]
port 19 nsew signal input
rlabel metal2 s 156326 165875 156382 166675 6 i_dout0[27]
port 20 nsew signal input
rlabel metal2 s 158258 165875 158314 166675 6 i_dout0[28]
port 21 nsew signal input
rlabel metal2 s 163410 0 163466 800 6 i_dout0[29]
port 22 nsew signal input
rlabel metal2 s 149978 0 150034 800 6 i_dout0[2]
port 23 nsew signal input
rlabel metal2 s 163042 165875 163098 166675 6 i_dout0[30]
port 24 nsew signal input
rlabel metal3 s 0 162528 800 162648 6 i_dout0[31]
port 25 nsew signal input
rlabel metal2 s 116398 165875 116454 166675 6 i_dout0[3]
port 26 nsew signal input
rlabel metal2 s 152922 0 152978 800 6 i_dout0[4]
port 27 nsew signal input
rlabel metal3 s 163731 38768 164531 38888 6 i_dout0[5]
port 28 nsew signal input
rlabel metal3 s 163731 44208 164531 44328 6 i_dout0[6]
port 29 nsew signal input
rlabel metal2 s 155038 0 155094 800 6 i_dout0[7]
port 30 nsew signal input
rlabel metal3 s 163731 57672 164531 57792 6 i_dout0[8]
port 31 nsew signal input
rlabel metal2 s 133510 165875 133566 166675 6 i_dout0[9]
port 32 nsew signal input
rlabel metal2 s 146942 0 146998 800 6 i_dout0_1[0]
port 33 nsew signal input
rlabel metal3 s 163731 73720 164531 73840 6 i_dout0_1[10]
port 34 nsew signal input
rlabel metal2 s 135442 165875 135498 166675 6 i_dout0_1[11]
port 35 nsew signal input
rlabel metal3 s 0 71136 800 71256 6 i_dout0_1[12]
port 36 nsew signal input
rlabel metal3 s 0 76440 800 76560 6 i_dout0_1[13]
port 37 nsew signal input
rlabel metal3 s 163731 95344 164531 95464 6 i_dout0_1[14]
port 38 nsew signal input
rlabel metal3 s 0 89904 800 90024 6 i_dout0_1[15]
port 39 nsew signal input
rlabel metal3 s 0 97928 800 98048 6 i_dout0_1[16]
port 40 nsew signal input
rlabel metal2 s 143998 165875 144054 166675 6 i_dout0_1[17]
port 41 nsew signal input
rlabel metal2 s 144918 165875 144974 166675 6 i_dout0_1[18]
port 42 nsew signal input
rlabel metal2 s 146850 165875 146906 166675 6 i_dout0_1[19]
port 43 nsew signal input
rlabel metal3 s 163731 11976 164531 12096 6 i_dout0_1[1]
port 44 nsew signal input
rlabel metal2 s 159178 0 159234 800 6 i_dout0_1[20]
port 45 nsew signal input
rlabel metal3 s 163731 127576 164531 127696 6 i_dout0_1[21]
port 46 nsew signal input
rlabel metal2 s 149702 165875 149758 166675 6 i_dout0_1[22]
port 47 nsew signal input
rlabel metal2 s 161018 0 161074 800 6 i_dout0_1[23]
port 48 nsew signal input
rlabel metal3 s 163731 141040 164531 141160 6 i_dout0_1[24]
port 49 nsew signal input
rlabel metal3 s 0 132880 800 133000 6 i_dout0_1[25]
port 50 nsew signal input
rlabel metal2 s 161846 0 161902 800 6 i_dout0_1[26]
port 51 nsew signal input
rlabel metal2 s 162490 0 162546 800 6 i_dout0_1[27]
port 52 nsew signal input
rlabel metal3 s 163731 151784 164531 151904 6 i_dout0_1[28]
port 53 nsew signal input
rlabel metal2 s 159178 165875 159234 166675 6 i_dout0_1[29]
port 54 nsew signal input
rlabel metal2 s 149702 0 149758 800 6 i_dout0_1[2]
port 55 nsew signal input
rlabel metal2 s 163962 0 164018 800 6 i_dout0_1[30]
port 56 nsew signal input
rlabel metal3 s 163731 159808 164531 159928 6 i_dout0_1[31]
port 57 nsew signal input
rlabel metal3 s 163731 30744 164531 30864 6 i_dout0_1[3]
port 58 nsew signal input
rlabel metal2 s 152646 0 152702 800 6 i_dout0_1[4]
port 59 nsew signal input
rlabel metal2 s 153198 0 153254 800 6 i_dout0_1[5]
port 60 nsew signal input
rlabel metal2 s 154394 0 154450 800 6 i_dout0_1[6]
port 61 nsew signal input
rlabel metal3 s 163731 52232 164531 52352 6 i_dout0_1[7]
port 62 nsew signal input
rlabel metal2 s 130658 165875 130714 166675 6 i_dout0_1[8]
port 63 nsew signal input
rlabel metal3 s 163731 65696 164531 65816 6 i_dout0_1[9]
port 64 nsew signal input
rlabel metal2 s 147310 0 147366 800 6 i_dout1[0]
port 65 nsew signal input
rlabel metal2 s 156510 0 156566 800 6 i_dout1[10]
port 66 nsew signal input
rlabel metal3 s 163731 84600 164531 84720 6 i_dout1[11]
port 67 nsew signal input
rlabel metal3 s 0 73720 800 73840 6 i_dout1[12]
port 68 nsew signal input
rlabel metal2 s 140226 165875 140282 166675 6 i_dout1[13]
port 69 nsew signal input
rlabel metal2 s 142066 165875 142122 166675 6 i_dout1[14]
port 70 nsew signal input
rlabel metal3 s 0 92624 800 92744 6 i_dout1[15]
port 71 nsew signal input
rlabel metal3 s 163731 106088 164531 106208 6 i_dout1[16]
port 72 nsew signal input
rlabel metal3 s 0 103368 800 103488 6 i_dout1[17]
port 73 nsew signal input
rlabel metal2 s 158258 0 158314 800 6 i_dout1[18]
port 74 nsew signal input
rlabel metal3 s 0 106088 800 106208 6 i_dout1[19]
port 75 nsew signal input
rlabel metal2 s 148506 0 148562 800 6 i_dout1[1]
port 76 nsew signal input
rlabel metal2 s 159454 0 159510 800 6 i_dout1[20]
port 77 nsew signal input
rlabel metal2 s 160098 0 160154 800 6 i_dout1[21]
port 78 nsew signal input
rlabel metal2 s 160650 0 160706 800 6 i_dout1[22]
port 79 nsew signal input
rlabel metal3 s 163731 138320 164531 138440 6 i_dout1[23]
port 80 nsew signal input
rlabel metal2 s 161570 0 161626 800 6 i_dout1[24]
port 81 nsew signal input
rlabel metal3 s 0 138320 800 138440 6 i_dout1[25]
port 82 nsew signal input
rlabel metal3 s 0 143760 800 143880 6 i_dout1[26]
port 83 nsew signal input
rlabel metal2 s 162766 0 162822 800 6 i_dout1[27]
port 84 nsew signal input
rlabel metal2 s 163042 0 163098 800 6 i_dout1[28]
port 85 nsew signal input
rlabel metal3 s 0 157088 800 157208 6 i_dout1[29]
port 86 nsew signal input
rlabel metal2 s 114558 165875 114614 166675 6 i_dout1[2]
port 87 nsew signal input
rlabel metal3 s 163731 157088 164531 157208 6 i_dout1[30]
port 88 nsew signal input
rlabel metal3 s 0 165248 800 165368 6 i_dout1[31]
port 89 nsew signal input
rlabel metal2 s 151174 0 151230 800 6 i_dout1[3]
port 90 nsew signal input
rlabel metal2 s 119250 165875 119306 166675 6 i_dout1[4]
port 91 nsew signal input
rlabel metal2 s 153842 0 153898 800 6 i_dout1[5]
port 92 nsew signal input
rlabel metal3 s 163731 46928 164531 47048 6 i_dout1[6]
port 93 nsew signal input
rlabel metal3 s 0 49512 800 49632 6 i_dout1[7]
port 94 nsew signal input
rlabel metal2 s 131670 165875 131726 166675 6 i_dout1[8]
port 95 nsew signal input
rlabel metal3 s 163731 68416 164531 68536 6 i_dout1[9]
port 96 nsew signal input
rlabel metal3 s 0 9256 800 9376 6 i_dout1_1[0]
port 97 nsew signal input
rlabel metal2 s 156234 0 156290 800 6 i_dout1_1[10]
port 98 nsew signal input
rlabel metal3 s 163731 79160 164531 79280 6 i_dout1_1[11]
port 99 nsew signal input
rlabel metal3 s 163731 89904 164531 90024 6 i_dout1_1[12]
port 100 nsew signal input
rlabel metal2 s 156786 0 156842 800 6 i_dout1_1[13]
port 101 nsew signal input
rlabel metal2 s 157154 0 157210 800 6 i_dout1_1[14]
port 102 nsew signal input
rlabel metal3 s 163731 97928 164531 98048 6 i_dout1_1[15]
port 103 nsew signal input
rlabel metal3 s 163731 103368 164531 103488 6 i_dout1_1[16]
port 104 nsew signal input
rlabel metal3 s 163731 111392 164531 111512 6 i_dout1_1[17]
port 105 nsew signal input
rlabel metal3 s 163731 119552 164531 119672 6 i_dout1_1[18]
port 106 nsew signal input
rlabel metal3 s 163731 122136 164531 122256 6 i_dout1_1[19]
port 107 nsew signal input
rlabel metal2 s 148138 0 148194 800 6 i_dout1_1[1]
port 108 nsew signal input
rlabel metal3 s 163731 124856 164531 124976 6 i_dout1_1[20]
port 109 nsew signal input
rlabel metal2 s 159822 0 159878 800 6 i_dout1_1[21]
port 110 nsew signal input
rlabel metal3 s 0 122136 800 122256 6 i_dout1_1[22]
port 111 nsew signal input
rlabel metal3 s 0 124856 800 124976 6 i_dout1_1[23]
port 112 nsew signal input
rlabel metal2 s 151634 165875 151690 166675 6 i_dout1_1[24]
port 113 nsew signal input
rlabel metal3 s 0 135600 800 135720 6 i_dout1_1[25]
port 114 nsew signal input
rlabel metal2 s 155406 165875 155462 166675 6 i_dout1_1[26]
port 115 nsew signal input
rlabel metal3 s 163731 149064 164531 149184 6 i_dout1_1[27]
port 116 nsew signal input
rlabel metal3 s 0 151784 800 151904 6 i_dout1_1[28]
port 117 nsew signal input
rlabel metal2 s 160190 165875 160246 166675 6 i_dout1_1[29]
port 118 nsew signal input
rlabel metal3 s 0 20000 800 20120 6 i_dout1_1[2]
port 119 nsew signal input
rlabel metal2 s 162030 165875 162086 166675 6 i_dout1_1[30]
port 120 nsew signal input
rlabel metal3 s 163731 162528 164531 162648 6 i_dout1_1[31]
port 121 nsew signal input
rlabel metal3 s 0 25304 800 25424 6 i_dout1_1[3]
port 122 nsew signal input
rlabel metal3 s 0 30744 800 30864 6 i_dout1_1[4]
port 123 nsew signal input
rlabel metal2 s 153566 0 153622 800 6 i_dout1_1[5]
port 124 nsew signal input
rlabel metal2 s 124954 165875 125010 166675 6 i_dout1_1[6]
port 125 nsew signal input
rlabel metal3 s 0 46928 800 47048 6 i_dout1_1[7]
port 126 nsew signal input
rlabel metal3 s 0 57672 800 57792 6 i_dout1_1[8]
port 127 nsew signal input
rlabel metal3 s 0 62976 800 63096 6 i_dout1_1[9]
port 128 nsew signal input
rlabel metal2 s 478 165875 534 166675 6 io_in[0]
port 129 nsew signal input
rlabel metal2 s 28998 165875 29054 166675 6 io_in[10]
port 130 nsew signal input
rlabel metal2 s 31850 165875 31906 166675 6 io_in[11]
port 131 nsew signal input
rlabel metal2 s 34702 165875 34758 166675 6 io_in[12]
port 132 nsew signal input
rlabel metal2 s 37554 165875 37610 166675 6 io_in[13]
port 133 nsew signal input
rlabel metal2 s 40406 165875 40462 166675 6 io_in[14]
port 134 nsew signal input
rlabel metal2 s 43258 165875 43314 166675 6 io_in[15]
port 135 nsew signal input
rlabel metal2 s 46110 165875 46166 166675 6 io_in[16]
port 136 nsew signal input
rlabel metal2 s 48962 165875 49018 166675 6 io_in[17]
port 137 nsew signal input
rlabel metal2 s 51814 165875 51870 166675 6 io_in[18]
port 138 nsew signal input
rlabel metal2 s 54666 165875 54722 166675 6 io_in[19]
port 139 nsew signal input
rlabel metal2 s 3330 165875 3386 166675 6 io_in[1]
port 140 nsew signal input
rlabel metal2 s 57518 165875 57574 166675 6 io_in[20]
port 141 nsew signal input
rlabel metal2 s 60370 165875 60426 166675 6 io_in[21]
port 142 nsew signal input
rlabel metal2 s 63222 165875 63278 166675 6 io_in[22]
port 143 nsew signal input
rlabel metal2 s 66074 165875 66130 166675 6 io_in[23]
port 144 nsew signal input
rlabel metal2 s 68926 165875 68982 166675 6 io_in[24]
port 145 nsew signal input
rlabel metal2 s 71778 165875 71834 166675 6 io_in[25]
port 146 nsew signal input
rlabel metal2 s 74630 165875 74686 166675 6 io_in[26]
port 147 nsew signal input
rlabel metal2 s 77482 165875 77538 166675 6 io_in[27]
port 148 nsew signal input
rlabel metal2 s 80334 165875 80390 166675 6 io_in[28]
port 149 nsew signal input
rlabel metal2 s 83186 165875 83242 166675 6 io_in[29]
port 150 nsew signal input
rlabel metal2 s 6182 165875 6238 166675 6 io_in[2]
port 151 nsew signal input
rlabel metal2 s 86038 165875 86094 166675 6 io_in[30]
port 152 nsew signal input
rlabel metal2 s 88890 165875 88946 166675 6 io_in[31]
port 153 nsew signal input
rlabel metal2 s 91742 165875 91798 166675 6 io_in[32]
port 154 nsew signal input
rlabel metal2 s 94594 165875 94650 166675 6 io_in[33]
port 155 nsew signal input
rlabel metal2 s 97446 165875 97502 166675 6 io_in[34]
port 156 nsew signal input
rlabel metal2 s 100298 165875 100354 166675 6 io_in[35]
port 157 nsew signal input
rlabel metal2 s 103150 165875 103206 166675 6 io_in[36]
port 158 nsew signal input
rlabel metal2 s 106002 165875 106058 166675 6 io_in[37]
port 159 nsew signal input
rlabel metal2 s 9034 165875 9090 166675 6 io_in[3]
port 160 nsew signal input
rlabel metal2 s 11886 165875 11942 166675 6 io_in[4]
port 161 nsew signal input
rlabel metal2 s 14738 165875 14794 166675 6 io_in[5]
port 162 nsew signal input
rlabel metal2 s 17590 165875 17646 166675 6 io_in[6]
port 163 nsew signal input
rlabel metal2 s 20442 165875 20498 166675 6 io_in[7]
port 164 nsew signal input
rlabel metal2 s 23294 165875 23350 166675 6 io_in[8]
port 165 nsew signal input
rlabel metal2 s 26146 165875 26202 166675 6 io_in[9]
port 166 nsew signal input
rlabel metal2 s 1398 165875 1454 166675 6 io_oeb[0]
port 167 nsew signal output
rlabel metal2 s 29918 165875 29974 166675 6 io_oeb[10]
port 168 nsew signal output
rlabel metal2 s 32770 165875 32826 166675 6 io_oeb[11]
port 169 nsew signal output
rlabel metal2 s 35622 165875 35678 166675 6 io_oeb[12]
port 170 nsew signal output
rlabel metal2 s 38474 165875 38530 166675 6 io_oeb[13]
port 171 nsew signal output
rlabel metal2 s 41326 165875 41382 166675 6 io_oeb[14]
port 172 nsew signal output
rlabel metal2 s 44178 165875 44234 166675 6 io_oeb[15]
port 173 nsew signal output
rlabel metal2 s 47030 165875 47086 166675 6 io_oeb[16]
port 174 nsew signal output
rlabel metal2 s 49882 165875 49938 166675 6 io_oeb[17]
port 175 nsew signal output
rlabel metal2 s 52734 165875 52790 166675 6 io_oeb[18]
port 176 nsew signal output
rlabel metal2 s 55586 165875 55642 166675 6 io_oeb[19]
port 177 nsew signal output
rlabel metal2 s 4250 165875 4306 166675 6 io_oeb[1]
port 178 nsew signal output
rlabel metal2 s 58438 165875 58494 166675 6 io_oeb[20]
port 179 nsew signal output
rlabel metal2 s 61290 165875 61346 166675 6 io_oeb[21]
port 180 nsew signal output
rlabel metal2 s 64142 165875 64198 166675 6 io_oeb[22]
port 181 nsew signal output
rlabel metal2 s 66994 165875 67050 166675 6 io_oeb[23]
port 182 nsew signal output
rlabel metal2 s 69846 165875 69902 166675 6 io_oeb[24]
port 183 nsew signal output
rlabel metal2 s 72698 165875 72754 166675 6 io_oeb[25]
port 184 nsew signal output
rlabel metal2 s 75550 165875 75606 166675 6 io_oeb[26]
port 185 nsew signal output
rlabel metal2 s 78402 165875 78458 166675 6 io_oeb[27]
port 186 nsew signal output
rlabel metal2 s 81254 165875 81310 166675 6 io_oeb[28]
port 187 nsew signal output
rlabel metal2 s 84106 165875 84162 166675 6 io_oeb[29]
port 188 nsew signal output
rlabel metal2 s 7102 165875 7158 166675 6 io_oeb[2]
port 189 nsew signal output
rlabel metal2 s 86958 165875 87014 166675 6 io_oeb[30]
port 190 nsew signal output
rlabel metal2 s 89810 165875 89866 166675 6 io_oeb[31]
port 191 nsew signal output
rlabel metal2 s 92662 165875 92718 166675 6 io_oeb[32]
port 192 nsew signal output
rlabel metal2 s 95514 165875 95570 166675 6 io_oeb[33]
port 193 nsew signal output
rlabel metal2 s 98366 165875 98422 166675 6 io_oeb[34]
port 194 nsew signal output
rlabel metal2 s 101218 165875 101274 166675 6 io_oeb[35]
port 195 nsew signal output
rlabel metal2 s 104070 165875 104126 166675 6 io_oeb[36]
port 196 nsew signal output
rlabel metal2 s 106922 165875 106978 166675 6 io_oeb[37]
port 197 nsew signal output
rlabel metal2 s 9954 165875 10010 166675 6 io_oeb[3]
port 198 nsew signal output
rlabel metal2 s 12806 165875 12862 166675 6 io_oeb[4]
port 199 nsew signal output
rlabel metal2 s 15658 165875 15714 166675 6 io_oeb[5]
port 200 nsew signal output
rlabel metal2 s 18510 165875 18566 166675 6 io_oeb[6]
port 201 nsew signal output
rlabel metal2 s 21362 165875 21418 166675 6 io_oeb[7]
port 202 nsew signal output
rlabel metal2 s 24214 165875 24270 166675 6 io_oeb[8]
port 203 nsew signal output
rlabel metal2 s 27066 165875 27122 166675 6 io_oeb[9]
port 204 nsew signal output
rlabel metal2 s 2318 165875 2374 166675 6 io_out[0]
port 205 nsew signal output
rlabel metal2 s 30838 165875 30894 166675 6 io_out[10]
port 206 nsew signal output
rlabel metal2 s 33690 165875 33746 166675 6 io_out[11]
port 207 nsew signal output
rlabel metal2 s 36542 165875 36598 166675 6 io_out[12]
port 208 nsew signal output
rlabel metal2 s 39394 165875 39450 166675 6 io_out[13]
port 209 nsew signal output
rlabel metal2 s 42246 165875 42302 166675 6 io_out[14]
port 210 nsew signal output
rlabel metal2 s 45098 165875 45154 166675 6 io_out[15]
port 211 nsew signal output
rlabel metal2 s 47950 165875 48006 166675 6 io_out[16]
port 212 nsew signal output
rlabel metal2 s 50802 165875 50858 166675 6 io_out[17]
port 213 nsew signal output
rlabel metal2 s 53654 165875 53710 166675 6 io_out[18]
port 214 nsew signal output
rlabel metal2 s 56506 165875 56562 166675 6 io_out[19]
port 215 nsew signal output
rlabel metal2 s 5170 165875 5226 166675 6 io_out[1]
port 216 nsew signal output
rlabel metal2 s 59358 165875 59414 166675 6 io_out[20]
port 217 nsew signal output
rlabel metal2 s 62210 165875 62266 166675 6 io_out[21]
port 218 nsew signal output
rlabel metal2 s 65062 165875 65118 166675 6 io_out[22]
port 219 nsew signal output
rlabel metal2 s 67914 165875 67970 166675 6 io_out[23]
port 220 nsew signal output
rlabel metal2 s 70766 165875 70822 166675 6 io_out[24]
port 221 nsew signal output
rlabel metal2 s 73618 165875 73674 166675 6 io_out[25]
port 222 nsew signal output
rlabel metal2 s 76470 165875 76526 166675 6 io_out[26]
port 223 nsew signal output
rlabel metal2 s 79322 165875 79378 166675 6 io_out[27]
port 224 nsew signal output
rlabel metal2 s 82174 165875 82230 166675 6 io_out[28]
port 225 nsew signal output
rlabel metal2 s 85026 165875 85082 166675 6 io_out[29]
port 226 nsew signal output
rlabel metal2 s 8022 165875 8078 166675 6 io_out[2]
port 227 nsew signal output
rlabel metal2 s 87878 165875 87934 166675 6 io_out[30]
port 228 nsew signal output
rlabel metal2 s 90730 165875 90786 166675 6 io_out[31]
port 229 nsew signal output
rlabel metal2 s 93582 165875 93638 166675 6 io_out[32]
port 230 nsew signal output
rlabel metal2 s 96434 165875 96490 166675 6 io_out[33]
port 231 nsew signal output
rlabel metal2 s 99286 165875 99342 166675 6 io_out[34]
port 232 nsew signal output
rlabel metal2 s 102138 165875 102194 166675 6 io_out[35]
port 233 nsew signal output
rlabel metal2 s 104990 165875 105046 166675 6 io_out[36]
port 234 nsew signal output
rlabel metal2 s 107842 165875 107898 166675 6 io_out[37]
port 235 nsew signal output
rlabel metal2 s 10874 165875 10930 166675 6 io_out[3]
port 236 nsew signal output
rlabel metal2 s 13726 165875 13782 166675 6 io_out[4]
port 237 nsew signal output
rlabel metal2 s 16578 165875 16634 166675 6 io_out[5]
port 238 nsew signal output
rlabel metal2 s 19430 165875 19486 166675 6 io_out[6]
port 239 nsew signal output
rlabel metal2 s 22282 165875 22338 166675 6 io_out[7]
port 240 nsew signal output
rlabel metal2 s 25134 165875 25190 166675 6 io_out[8]
port 241 nsew signal output
rlabel metal2 s 27986 165875 28042 166675 6 io_out[9]
port 242 nsew signal output
rlabel metal2 s 146114 0 146170 800 6 irq[0]
port 243 nsew signal output
rlabel metal2 s 146390 0 146446 800 6 irq[1]
port 244 nsew signal output
rlabel metal2 s 146666 0 146722 800 6 irq[2]
port 245 nsew signal output
rlabel metal2 s 31666 0 31722 800 6 la_data_in[0]
port 246 nsew signal input
rlabel metal2 s 121090 0 121146 800 6 la_data_in[100]
port 247 nsew signal input
rlabel metal2 s 121918 0 121974 800 6 la_data_in[101]
port 248 nsew signal input
rlabel metal2 s 122838 0 122894 800 6 la_data_in[102]
port 249 nsew signal input
rlabel metal2 s 123758 0 123814 800 6 la_data_in[103]
port 250 nsew signal input
rlabel metal2 s 124586 0 124642 800 6 la_data_in[104]
port 251 nsew signal input
rlabel metal2 s 125506 0 125562 800 6 la_data_in[105]
port 252 nsew signal input
rlabel metal2 s 126426 0 126482 800 6 la_data_in[106]
port 253 nsew signal input
rlabel metal2 s 127346 0 127402 800 6 la_data_in[107]
port 254 nsew signal input
rlabel metal2 s 128174 0 128230 800 6 la_data_in[108]
port 255 nsew signal input
rlabel metal2 s 129094 0 129150 800 6 la_data_in[109]
port 256 nsew signal input
rlabel metal2 s 40590 0 40646 800 6 la_data_in[10]
port 257 nsew signal input
rlabel metal2 s 130014 0 130070 800 6 la_data_in[110]
port 258 nsew signal input
rlabel metal2 s 130842 0 130898 800 6 la_data_in[111]
port 259 nsew signal input
rlabel metal2 s 131762 0 131818 800 6 la_data_in[112]
port 260 nsew signal input
rlabel metal2 s 132682 0 132738 800 6 la_data_in[113]
port 261 nsew signal input
rlabel metal2 s 133602 0 133658 800 6 la_data_in[114]
port 262 nsew signal input
rlabel metal2 s 134430 0 134486 800 6 la_data_in[115]
port 263 nsew signal input
rlabel metal2 s 135350 0 135406 800 6 la_data_in[116]
port 264 nsew signal input
rlabel metal2 s 136270 0 136326 800 6 la_data_in[117]
port 265 nsew signal input
rlabel metal2 s 137190 0 137246 800 6 la_data_in[118]
port 266 nsew signal input
rlabel metal2 s 138018 0 138074 800 6 la_data_in[119]
port 267 nsew signal input
rlabel metal2 s 41510 0 41566 800 6 la_data_in[11]
port 268 nsew signal input
rlabel metal2 s 138938 0 138994 800 6 la_data_in[120]
port 269 nsew signal input
rlabel metal2 s 139858 0 139914 800 6 la_data_in[121]
port 270 nsew signal input
rlabel metal2 s 140686 0 140742 800 6 la_data_in[122]
port 271 nsew signal input
rlabel metal2 s 141606 0 141662 800 6 la_data_in[123]
port 272 nsew signal input
rlabel metal2 s 142526 0 142582 800 6 la_data_in[124]
port 273 nsew signal input
rlabel metal2 s 143446 0 143502 800 6 la_data_in[125]
port 274 nsew signal input
rlabel metal2 s 144274 0 144330 800 6 la_data_in[126]
port 275 nsew signal input
rlabel metal2 s 145194 0 145250 800 6 la_data_in[127]
port 276 nsew signal input
rlabel metal2 s 42338 0 42394 800 6 la_data_in[12]
port 277 nsew signal input
rlabel metal2 s 43258 0 43314 800 6 la_data_in[13]
port 278 nsew signal input
rlabel metal2 s 44178 0 44234 800 6 la_data_in[14]
port 279 nsew signal input
rlabel metal2 s 45098 0 45154 800 6 la_data_in[15]
port 280 nsew signal input
rlabel metal2 s 45926 0 45982 800 6 la_data_in[16]
port 281 nsew signal input
rlabel metal2 s 46846 0 46902 800 6 la_data_in[17]
port 282 nsew signal input
rlabel metal2 s 47766 0 47822 800 6 la_data_in[18]
port 283 nsew signal input
rlabel metal2 s 48594 0 48650 800 6 la_data_in[19]
port 284 nsew signal input
rlabel metal2 s 32586 0 32642 800 6 la_data_in[1]
port 285 nsew signal input
rlabel metal2 s 49514 0 49570 800 6 la_data_in[20]
port 286 nsew signal input
rlabel metal2 s 50434 0 50490 800 6 la_data_in[21]
port 287 nsew signal input
rlabel metal2 s 51354 0 51410 800 6 la_data_in[22]
port 288 nsew signal input
rlabel metal2 s 52182 0 52238 800 6 la_data_in[23]
port 289 nsew signal input
rlabel metal2 s 53102 0 53158 800 6 la_data_in[24]
port 290 nsew signal input
rlabel metal2 s 54022 0 54078 800 6 la_data_in[25]
port 291 nsew signal input
rlabel metal2 s 54942 0 54998 800 6 la_data_in[26]
port 292 nsew signal input
rlabel metal2 s 55770 0 55826 800 6 la_data_in[27]
port 293 nsew signal input
rlabel metal2 s 56690 0 56746 800 6 la_data_in[28]
port 294 nsew signal input
rlabel metal2 s 57610 0 57666 800 6 la_data_in[29]
port 295 nsew signal input
rlabel metal2 s 33414 0 33470 800 6 la_data_in[2]
port 296 nsew signal input
rlabel metal2 s 58438 0 58494 800 6 la_data_in[30]
port 297 nsew signal input
rlabel metal2 s 59358 0 59414 800 6 la_data_in[31]
port 298 nsew signal input
rlabel metal2 s 60278 0 60334 800 6 la_data_in[32]
port 299 nsew signal input
rlabel metal2 s 61198 0 61254 800 6 la_data_in[33]
port 300 nsew signal input
rlabel metal2 s 62026 0 62082 800 6 la_data_in[34]
port 301 nsew signal input
rlabel metal2 s 62946 0 63002 800 6 la_data_in[35]
port 302 nsew signal input
rlabel metal2 s 63866 0 63922 800 6 la_data_in[36]
port 303 nsew signal input
rlabel metal2 s 64694 0 64750 800 6 la_data_in[37]
port 304 nsew signal input
rlabel metal2 s 65614 0 65670 800 6 la_data_in[38]
port 305 nsew signal input
rlabel metal2 s 66534 0 66590 800 6 la_data_in[39]
port 306 nsew signal input
rlabel metal2 s 34334 0 34390 800 6 la_data_in[3]
port 307 nsew signal input
rlabel metal2 s 67454 0 67510 800 6 la_data_in[40]
port 308 nsew signal input
rlabel metal2 s 68282 0 68338 800 6 la_data_in[41]
port 309 nsew signal input
rlabel metal2 s 69202 0 69258 800 6 la_data_in[42]
port 310 nsew signal input
rlabel metal2 s 70122 0 70178 800 6 la_data_in[43]
port 311 nsew signal input
rlabel metal2 s 70950 0 71006 800 6 la_data_in[44]
port 312 nsew signal input
rlabel metal2 s 71870 0 71926 800 6 la_data_in[45]
port 313 nsew signal input
rlabel metal2 s 72790 0 72846 800 6 la_data_in[46]
port 314 nsew signal input
rlabel metal2 s 73710 0 73766 800 6 la_data_in[47]
port 315 nsew signal input
rlabel metal2 s 74538 0 74594 800 6 la_data_in[48]
port 316 nsew signal input
rlabel metal2 s 75458 0 75514 800 6 la_data_in[49]
port 317 nsew signal input
rlabel metal2 s 35254 0 35310 800 6 la_data_in[4]
port 318 nsew signal input
rlabel metal2 s 76378 0 76434 800 6 la_data_in[50]
port 319 nsew signal input
rlabel metal2 s 77206 0 77262 800 6 la_data_in[51]
port 320 nsew signal input
rlabel metal2 s 78126 0 78182 800 6 la_data_in[52]
port 321 nsew signal input
rlabel metal2 s 79046 0 79102 800 6 la_data_in[53]
port 322 nsew signal input
rlabel metal2 s 79966 0 80022 800 6 la_data_in[54]
port 323 nsew signal input
rlabel metal2 s 80794 0 80850 800 6 la_data_in[55]
port 324 nsew signal input
rlabel metal2 s 81714 0 81770 800 6 la_data_in[56]
port 325 nsew signal input
rlabel metal2 s 82634 0 82690 800 6 la_data_in[57]
port 326 nsew signal input
rlabel metal2 s 83462 0 83518 800 6 la_data_in[58]
port 327 nsew signal input
rlabel metal2 s 84382 0 84438 800 6 la_data_in[59]
port 328 nsew signal input
rlabel metal2 s 36082 0 36138 800 6 la_data_in[5]
port 329 nsew signal input
rlabel metal2 s 85302 0 85358 800 6 la_data_in[60]
port 330 nsew signal input
rlabel metal2 s 86222 0 86278 800 6 la_data_in[61]
port 331 nsew signal input
rlabel metal2 s 87050 0 87106 800 6 la_data_in[62]
port 332 nsew signal input
rlabel metal2 s 87970 0 88026 800 6 la_data_in[63]
port 333 nsew signal input
rlabel metal2 s 88890 0 88946 800 6 la_data_in[64]
port 334 nsew signal input
rlabel metal2 s 89718 0 89774 800 6 la_data_in[65]
port 335 nsew signal input
rlabel metal2 s 90638 0 90694 800 6 la_data_in[66]
port 336 nsew signal input
rlabel metal2 s 91558 0 91614 800 6 la_data_in[67]
port 337 nsew signal input
rlabel metal2 s 92478 0 92534 800 6 la_data_in[68]
port 338 nsew signal input
rlabel metal2 s 93306 0 93362 800 6 la_data_in[69]
port 339 nsew signal input
rlabel metal2 s 37002 0 37058 800 6 la_data_in[6]
port 340 nsew signal input
rlabel metal2 s 94226 0 94282 800 6 la_data_in[70]
port 341 nsew signal input
rlabel metal2 s 95146 0 95202 800 6 la_data_in[71]
port 342 nsew signal input
rlabel metal2 s 96066 0 96122 800 6 la_data_in[72]
port 343 nsew signal input
rlabel metal2 s 96894 0 96950 800 6 la_data_in[73]
port 344 nsew signal input
rlabel metal2 s 97814 0 97870 800 6 la_data_in[74]
port 345 nsew signal input
rlabel metal2 s 98734 0 98790 800 6 la_data_in[75]
port 346 nsew signal input
rlabel metal2 s 99562 0 99618 800 6 la_data_in[76]
port 347 nsew signal input
rlabel metal2 s 100482 0 100538 800 6 la_data_in[77]
port 348 nsew signal input
rlabel metal2 s 101402 0 101458 800 6 la_data_in[78]
port 349 nsew signal input
rlabel metal2 s 102322 0 102378 800 6 la_data_in[79]
port 350 nsew signal input
rlabel metal2 s 37922 0 37978 800 6 la_data_in[7]
port 351 nsew signal input
rlabel metal2 s 103150 0 103206 800 6 la_data_in[80]
port 352 nsew signal input
rlabel metal2 s 104070 0 104126 800 6 la_data_in[81]
port 353 nsew signal input
rlabel metal2 s 104990 0 105046 800 6 la_data_in[82]
port 354 nsew signal input
rlabel metal2 s 105818 0 105874 800 6 la_data_in[83]
port 355 nsew signal input
rlabel metal2 s 106738 0 106794 800 6 la_data_in[84]
port 356 nsew signal input
rlabel metal2 s 107658 0 107714 800 6 la_data_in[85]
port 357 nsew signal input
rlabel metal2 s 108578 0 108634 800 6 la_data_in[86]
port 358 nsew signal input
rlabel metal2 s 109406 0 109462 800 6 la_data_in[87]
port 359 nsew signal input
rlabel metal2 s 110326 0 110382 800 6 la_data_in[88]
port 360 nsew signal input
rlabel metal2 s 111246 0 111302 800 6 la_data_in[89]
port 361 nsew signal input
rlabel metal2 s 38842 0 38898 800 6 la_data_in[8]
port 362 nsew signal input
rlabel metal2 s 112074 0 112130 800 6 la_data_in[90]
port 363 nsew signal input
rlabel metal2 s 112994 0 113050 800 6 la_data_in[91]
port 364 nsew signal input
rlabel metal2 s 113914 0 113970 800 6 la_data_in[92]
port 365 nsew signal input
rlabel metal2 s 114834 0 114890 800 6 la_data_in[93]
port 366 nsew signal input
rlabel metal2 s 115662 0 115718 800 6 la_data_in[94]
port 367 nsew signal input
rlabel metal2 s 116582 0 116638 800 6 la_data_in[95]
port 368 nsew signal input
rlabel metal2 s 117502 0 117558 800 6 la_data_in[96]
port 369 nsew signal input
rlabel metal2 s 118330 0 118386 800 6 la_data_in[97]
port 370 nsew signal input
rlabel metal2 s 119250 0 119306 800 6 la_data_in[98]
port 371 nsew signal input
rlabel metal2 s 120170 0 120226 800 6 la_data_in[99]
port 372 nsew signal input
rlabel metal2 s 39670 0 39726 800 6 la_data_in[9]
port 373 nsew signal input
rlabel metal2 s 31942 0 31998 800 6 la_data_out[0]
port 374 nsew signal output
rlabel metal2 s 121366 0 121422 800 6 la_data_out[100]
port 375 nsew signal output
rlabel metal2 s 122286 0 122342 800 6 la_data_out[101]
port 376 nsew signal output
rlabel metal2 s 123114 0 123170 800 6 la_data_out[102]
port 377 nsew signal output
rlabel metal2 s 124034 0 124090 800 6 la_data_out[103]
port 378 nsew signal output
rlabel metal2 s 124954 0 125010 800 6 la_data_out[104]
port 379 nsew signal output
rlabel metal2 s 125782 0 125838 800 6 la_data_out[105]
port 380 nsew signal output
rlabel metal2 s 126702 0 126758 800 6 la_data_out[106]
port 381 nsew signal output
rlabel metal2 s 127622 0 127678 800 6 la_data_out[107]
port 382 nsew signal output
rlabel metal2 s 128542 0 128598 800 6 la_data_out[108]
port 383 nsew signal output
rlabel metal2 s 129370 0 129426 800 6 la_data_out[109]
port 384 nsew signal output
rlabel metal2 s 40866 0 40922 800 6 la_data_out[10]
port 385 nsew signal output
rlabel metal2 s 130290 0 130346 800 6 la_data_out[110]
port 386 nsew signal output
rlabel metal2 s 131210 0 131266 800 6 la_data_out[111]
port 387 nsew signal output
rlabel metal2 s 132038 0 132094 800 6 la_data_out[112]
port 388 nsew signal output
rlabel metal2 s 132958 0 133014 800 6 la_data_out[113]
port 389 nsew signal output
rlabel metal2 s 133878 0 133934 800 6 la_data_out[114]
port 390 nsew signal output
rlabel metal2 s 134798 0 134854 800 6 la_data_out[115]
port 391 nsew signal output
rlabel metal2 s 135626 0 135682 800 6 la_data_out[116]
port 392 nsew signal output
rlabel metal2 s 136546 0 136602 800 6 la_data_out[117]
port 393 nsew signal output
rlabel metal2 s 137466 0 137522 800 6 la_data_out[118]
port 394 nsew signal output
rlabel metal2 s 138294 0 138350 800 6 la_data_out[119]
port 395 nsew signal output
rlabel metal2 s 41786 0 41842 800 6 la_data_out[11]
port 396 nsew signal output
rlabel metal2 s 139214 0 139270 800 6 la_data_out[120]
port 397 nsew signal output
rlabel metal2 s 140134 0 140190 800 6 la_data_out[121]
port 398 nsew signal output
rlabel metal2 s 141054 0 141110 800 6 la_data_out[122]
port 399 nsew signal output
rlabel metal2 s 141882 0 141938 800 6 la_data_out[123]
port 400 nsew signal output
rlabel metal2 s 142802 0 142858 800 6 la_data_out[124]
port 401 nsew signal output
rlabel metal2 s 143722 0 143778 800 6 la_data_out[125]
port 402 nsew signal output
rlabel metal2 s 144550 0 144606 800 6 la_data_out[126]
port 403 nsew signal output
rlabel metal2 s 145470 0 145526 800 6 la_data_out[127]
port 404 nsew signal output
rlabel metal2 s 42706 0 42762 800 6 la_data_out[12]
port 405 nsew signal output
rlabel metal2 s 43534 0 43590 800 6 la_data_out[13]
port 406 nsew signal output
rlabel metal2 s 44454 0 44510 800 6 la_data_out[14]
port 407 nsew signal output
rlabel metal2 s 45374 0 45430 800 6 la_data_out[15]
port 408 nsew signal output
rlabel metal2 s 46294 0 46350 800 6 la_data_out[16]
port 409 nsew signal output
rlabel metal2 s 47122 0 47178 800 6 la_data_out[17]
port 410 nsew signal output
rlabel metal2 s 48042 0 48098 800 6 la_data_out[18]
port 411 nsew signal output
rlabel metal2 s 48962 0 49018 800 6 la_data_out[19]
port 412 nsew signal output
rlabel metal2 s 32862 0 32918 800 6 la_data_out[1]
port 413 nsew signal output
rlabel metal2 s 49790 0 49846 800 6 la_data_out[20]
port 414 nsew signal output
rlabel metal2 s 50710 0 50766 800 6 la_data_out[21]
port 415 nsew signal output
rlabel metal2 s 51630 0 51686 800 6 la_data_out[22]
port 416 nsew signal output
rlabel metal2 s 52550 0 52606 800 6 la_data_out[23]
port 417 nsew signal output
rlabel metal2 s 53378 0 53434 800 6 la_data_out[24]
port 418 nsew signal output
rlabel metal2 s 54298 0 54354 800 6 la_data_out[25]
port 419 nsew signal output
rlabel metal2 s 55218 0 55274 800 6 la_data_out[26]
port 420 nsew signal output
rlabel metal2 s 56046 0 56102 800 6 la_data_out[27]
port 421 nsew signal output
rlabel metal2 s 56966 0 57022 800 6 la_data_out[28]
port 422 nsew signal output
rlabel metal2 s 57886 0 57942 800 6 la_data_out[29]
port 423 nsew signal output
rlabel metal2 s 33782 0 33838 800 6 la_data_out[2]
port 424 nsew signal output
rlabel metal2 s 58806 0 58862 800 6 la_data_out[30]
port 425 nsew signal output
rlabel metal2 s 59634 0 59690 800 6 la_data_out[31]
port 426 nsew signal output
rlabel metal2 s 60554 0 60610 800 6 la_data_out[32]
port 427 nsew signal output
rlabel metal2 s 61474 0 61530 800 6 la_data_out[33]
port 428 nsew signal output
rlabel metal2 s 62302 0 62358 800 6 la_data_out[34]
port 429 nsew signal output
rlabel metal2 s 63222 0 63278 800 6 la_data_out[35]
port 430 nsew signal output
rlabel metal2 s 64142 0 64198 800 6 la_data_out[36]
port 431 nsew signal output
rlabel metal2 s 65062 0 65118 800 6 la_data_out[37]
port 432 nsew signal output
rlabel metal2 s 65890 0 65946 800 6 la_data_out[38]
port 433 nsew signal output
rlabel metal2 s 66810 0 66866 800 6 la_data_out[39]
port 434 nsew signal output
rlabel metal2 s 34610 0 34666 800 6 la_data_out[3]
port 435 nsew signal output
rlabel metal2 s 67730 0 67786 800 6 la_data_out[40]
port 436 nsew signal output
rlabel metal2 s 68650 0 68706 800 6 la_data_out[41]
port 437 nsew signal output
rlabel metal2 s 69478 0 69534 800 6 la_data_out[42]
port 438 nsew signal output
rlabel metal2 s 70398 0 70454 800 6 la_data_out[43]
port 439 nsew signal output
rlabel metal2 s 71318 0 71374 800 6 la_data_out[44]
port 440 nsew signal output
rlabel metal2 s 72146 0 72202 800 6 la_data_out[45]
port 441 nsew signal output
rlabel metal2 s 73066 0 73122 800 6 la_data_out[46]
port 442 nsew signal output
rlabel metal2 s 73986 0 74042 800 6 la_data_out[47]
port 443 nsew signal output
rlabel metal2 s 74906 0 74962 800 6 la_data_out[48]
port 444 nsew signal output
rlabel metal2 s 75734 0 75790 800 6 la_data_out[49]
port 445 nsew signal output
rlabel metal2 s 35530 0 35586 800 6 la_data_out[4]
port 446 nsew signal output
rlabel metal2 s 76654 0 76710 800 6 la_data_out[50]
port 447 nsew signal output
rlabel metal2 s 77574 0 77630 800 6 la_data_out[51]
port 448 nsew signal output
rlabel metal2 s 78402 0 78458 800 6 la_data_out[52]
port 449 nsew signal output
rlabel metal2 s 79322 0 79378 800 6 la_data_out[53]
port 450 nsew signal output
rlabel metal2 s 80242 0 80298 800 6 la_data_out[54]
port 451 nsew signal output
rlabel metal2 s 81162 0 81218 800 6 la_data_out[55]
port 452 nsew signal output
rlabel metal2 s 81990 0 82046 800 6 la_data_out[56]
port 453 nsew signal output
rlabel metal2 s 82910 0 82966 800 6 la_data_out[57]
port 454 nsew signal output
rlabel metal2 s 83830 0 83886 800 6 la_data_out[58]
port 455 nsew signal output
rlabel metal2 s 84658 0 84714 800 6 la_data_out[59]
port 456 nsew signal output
rlabel metal2 s 36450 0 36506 800 6 la_data_out[5]
port 457 nsew signal output
rlabel metal2 s 85578 0 85634 800 6 la_data_out[60]
port 458 nsew signal output
rlabel metal2 s 86498 0 86554 800 6 la_data_out[61]
port 459 nsew signal output
rlabel metal2 s 87418 0 87474 800 6 la_data_out[62]
port 460 nsew signal output
rlabel metal2 s 88246 0 88302 800 6 la_data_out[63]
port 461 nsew signal output
rlabel metal2 s 89166 0 89222 800 6 la_data_out[64]
port 462 nsew signal output
rlabel metal2 s 90086 0 90142 800 6 la_data_out[65]
port 463 nsew signal output
rlabel metal2 s 90914 0 90970 800 6 la_data_out[66]
port 464 nsew signal output
rlabel metal2 s 91834 0 91890 800 6 la_data_out[67]
port 465 nsew signal output
rlabel metal2 s 92754 0 92810 800 6 la_data_out[68]
port 466 nsew signal output
rlabel metal2 s 93674 0 93730 800 6 la_data_out[69]
port 467 nsew signal output
rlabel metal2 s 37278 0 37334 800 6 la_data_out[6]
port 468 nsew signal output
rlabel metal2 s 94502 0 94558 800 6 la_data_out[70]
port 469 nsew signal output
rlabel metal2 s 95422 0 95478 800 6 la_data_out[71]
port 470 nsew signal output
rlabel metal2 s 96342 0 96398 800 6 la_data_out[72]
port 471 nsew signal output
rlabel metal2 s 97170 0 97226 800 6 la_data_out[73]
port 472 nsew signal output
rlabel metal2 s 98090 0 98146 800 6 la_data_out[74]
port 473 nsew signal output
rlabel metal2 s 99010 0 99066 800 6 la_data_out[75]
port 474 nsew signal output
rlabel metal2 s 99930 0 99986 800 6 la_data_out[76]
port 475 nsew signal output
rlabel metal2 s 100758 0 100814 800 6 la_data_out[77]
port 476 nsew signal output
rlabel metal2 s 101678 0 101734 800 6 la_data_out[78]
port 477 nsew signal output
rlabel metal2 s 102598 0 102654 800 6 la_data_out[79]
port 478 nsew signal output
rlabel metal2 s 38198 0 38254 800 6 la_data_out[7]
port 479 nsew signal output
rlabel metal2 s 103426 0 103482 800 6 la_data_out[80]
port 480 nsew signal output
rlabel metal2 s 104346 0 104402 800 6 la_data_out[81]
port 481 nsew signal output
rlabel metal2 s 105266 0 105322 800 6 la_data_out[82]
port 482 nsew signal output
rlabel metal2 s 106186 0 106242 800 6 la_data_out[83]
port 483 nsew signal output
rlabel metal2 s 107014 0 107070 800 6 la_data_out[84]
port 484 nsew signal output
rlabel metal2 s 107934 0 107990 800 6 la_data_out[85]
port 485 nsew signal output
rlabel metal2 s 108854 0 108910 800 6 la_data_out[86]
port 486 nsew signal output
rlabel metal2 s 109774 0 109830 800 6 la_data_out[87]
port 487 nsew signal output
rlabel metal2 s 110602 0 110658 800 6 la_data_out[88]
port 488 nsew signal output
rlabel metal2 s 111522 0 111578 800 6 la_data_out[89]
port 489 nsew signal output
rlabel metal2 s 39118 0 39174 800 6 la_data_out[8]
port 490 nsew signal output
rlabel metal2 s 112442 0 112498 800 6 la_data_out[90]
port 491 nsew signal output
rlabel metal2 s 113270 0 113326 800 6 la_data_out[91]
port 492 nsew signal output
rlabel metal2 s 114190 0 114246 800 6 la_data_out[92]
port 493 nsew signal output
rlabel metal2 s 115110 0 115166 800 6 la_data_out[93]
port 494 nsew signal output
rlabel metal2 s 116030 0 116086 800 6 la_data_out[94]
port 495 nsew signal output
rlabel metal2 s 116858 0 116914 800 6 la_data_out[95]
port 496 nsew signal output
rlabel metal2 s 117778 0 117834 800 6 la_data_out[96]
port 497 nsew signal output
rlabel metal2 s 118698 0 118754 800 6 la_data_out[97]
port 498 nsew signal output
rlabel metal2 s 119526 0 119582 800 6 la_data_out[98]
port 499 nsew signal output
rlabel metal2 s 120446 0 120502 800 6 la_data_out[99]
port 500 nsew signal output
rlabel metal2 s 40038 0 40094 800 6 la_data_out[9]
port 501 nsew signal output
rlabel metal2 s 32218 0 32274 800 6 la_oenb[0]
port 502 nsew signal input
rlabel metal2 s 121642 0 121698 800 6 la_oenb[100]
port 503 nsew signal input
rlabel metal2 s 122562 0 122618 800 6 la_oenb[101]
port 504 nsew signal input
rlabel metal2 s 123482 0 123538 800 6 la_oenb[102]
port 505 nsew signal input
rlabel metal2 s 124310 0 124366 800 6 la_oenb[103]
port 506 nsew signal input
rlabel metal2 s 125230 0 125286 800 6 la_oenb[104]
port 507 nsew signal input
rlabel metal2 s 126150 0 126206 800 6 la_oenb[105]
port 508 nsew signal input
rlabel metal2 s 126978 0 127034 800 6 la_oenb[106]
port 509 nsew signal input
rlabel metal2 s 127898 0 127954 800 6 la_oenb[107]
port 510 nsew signal input
rlabel metal2 s 128818 0 128874 800 6 la_oenb[108]
port 511 nsew signal input
rlabel metal2 s 129738 0 129794 800 6 la_oenb[109]
port 512 nsew signal input
rlabel metal2 s 41234 0 41290 800 6 la_oenb[10]
port 513 nsew signal input
rlabel metal2 s 130566 0 130622 800 6 la_oenb[110]
port 514 nsew signal input
rlabel metal2 s 131486 0 131542 800 6 la_oenb[111]
port 515 nsew signal input
rlabel metal2 s 132406 0 132462 800 6 la_oenb[112]
port 516 nsew signal input
rlabel metal2 s 133234 0 133290 800 6 la_oenb[113]
port 517 nsew signal input
rlabel metal2 s 134154 0 134210 800 6 la_oenb[114]
port 518 nsew signal input
rlabel metal2 s 135074 0 135130 800 6 la_oenb[115]
port 519 nsew signal input
rlabel metal2 s 135994 0 136050 800 6 la_oenb[116]
port 520 nsew signal input
rlabel metal2 s 136822 0 136878 800 6 la_oenb[117]
port 521 nsew signal input
rlabel metal2 s 137742 0 137798 800 6 la_oenb[118]
port 522 nsew signal input
rlabel metal2 s 138662 0 138718 800 6 la_oenb[119]
port 523 nsew signal input
rlabel metal2 s 42062 0 42118 800 6 la_oenb[11]
port 524 nsew signal input
rlabel metal2 s 139490 0 139546 800 6 la_oenb[120]
port 525 nsew signal input
rlabel metal2 s 140410 0 140466 800 6 la_oenb[121]
port 526 nsew signal input
rlabel metal2 s 141330 0 141386 800 6 la_oenb[122]
port 527 nsew signal input
rlabel metal2 s 142250 0 142306 800 6 la_oenb[123]
port 528 nsew signal input
rlabel metal2 s 143078 0 143134 800 6 la_oenb[124]
port 529 nsew signal input
rlabel metal2 s 143998 0 144054 800 6 la_oenb[125]
port 530 nsew signal input
rlabel metal2 s 144918 0 144974 800 6 la_oenb[126]
port 531 nsew signal input
rlabel metal2 s 145746 0 145802 800 6 la_oenb[127]
port 532 nsew signal input
rlabel metal2 s 42982 0 43038 800 6 la_oenb[12]
port 533 nsew signal input
rlabel metal2 s 43902 0 43958 800 6 la_oenb[13]
port 534 nsew signal input
rlabel metal2 s 44730 0 44786 800 6 la_oenb[14]
port 535 nsew signal input
rlabel metal2 s 45650 0 45706 800 6 la_oenb[15]
port 536 nsew signal input
rlabel metal2 s 46570 0 46626 800 6 la_oenb[16]
port 537 nsew signal input
rlabel metal2 s 47490 0 47546 800 6 la_oenb[17]
port 538 nsew signal input
rlabel metal2 s 48318 0 48374 800 6 la_oenb[18]
port 539 nsew signal input
rlabel metal2 s 49238 0 49294 800 6 la_oenb[19]
port 540 nsew signal input
rlabel metal2 s 33138 0 33194 800 6 la_oenb[1]
port 541 nsew signal input
rlabel metal2 s 50158 0 50214 800 6 la_oenb[20]
port 542 nsew signal input
rlabel metal2 s 50986 0 51042 800 6 la_oenb[21]
port 543 nsew signal input
rlabel metal2 s 51906 0 51962 800 6 la_oenb[22]
port 544 nsew signal input
rlabel metal2 s 52826 0 52882 800 6 la_oenb[23]
port 545 nsew signal input
rlabel metal2 s 53746 0 53802 800 6 la_oenb[24]
port 546 nsew signal input
rlabel metal2 s 54574 0 54630 800 6 la_oenb[25]
port 547 nsew signal input
rlabel metal2 s 55494 0 55550 800 6 la_oenb[26]
port 548 nsew signal input
rlabel metal2 s 56414 0 56470 800 6 la_oenb[27]
port 549 nsew signal input
rlabel metal2 s 57242 0 57298 800 6 la_oenb[28]
port 550 nsew signal input
rlabel metal2 s 58162 0 58218 800 6 la_oenb[29]
port 551 nsew signal input
rlabel metal2 s 34058 0 34114 800 6 la_oenb[2]
port 552 nsew signal input
rlabel metal2 s 59082 0 59138 800 6 la_oenb[30]
port 553 nsew signal input
rlabel metal2 s 60002 0 60058 800 6 la_oenb[31]
port 554 nsew signal input
rlabel metal2 s 60830 0 60886 800 6 la_oenb[32]
port 555 nsew signal input
rlabel metal2 s 61750 0 61806 800 6 la_oenb[33]
port 556 nsew signal input
rlabel metal2 s 62670 0 62726 800 6 la_oenb[34]
port 557 nsew signal input
rlabel metal2 s 63498 0 63554 800 6 la_oenb[35]
port 558 nsew signal input
rlabel metal2 s 64418 0 64474 800 6 la_oenb[36]
port 559 nsew signal input
rlabel metal2 s 65338 0 65394 800 6 la_oenb[37]
port 560 nsew signal input
rlabel metal2 s 66258 0 66314 800 6 la_oenb[38]
port 561 nsew signal input
rlabel metal2 s 67086 0 67142 800 6 la_oenb[39]
port 562 nsew signal input
rlabel metal2 s 34886 0 34942 800 6 la_oenb[3]
port 563 nsew signal input
rlabel metal2 s 68006 0 68062 800 6 la_oenb[40]
port 564 nsew signal input
rlabel metal2 s 68926 0 68982 800 6 la_oenb[41]
port 565 nsew signal input
rlabel metal2 s 69754 0 69810 800 6 la_oenb[42]
port 566 nsew signal input
rlabel metal2 s 70674 0 70730 800 6 la_oenb[43]
port 567 nsew signal input
rlabel metal2 s 71594 0 71650 800 6 la_oenb[44]
port 568 nsew signal input
rlabel metal2 s 72514 0 72570 800 6 la_oenb[45]
port 569 nsew signal input
rlabel metal2 s 73342 0 73398 800 6 la_oenb[46]
port 570 nsew signal input
rlabel metal2 s 74262 0 74318 800 6 la_oenb[47]
port 571 nsew signal input
rlabel metal2 s 75182 0 75238 800 6 la_oenb[48]
port 572 nsew signal input
rlabel metal2 s 76010 0 76066 800 6 la_oenb[49]
port 573 nsew signal input
rlabel metal2 s 35806 0 35862 800 6 la_oenb[4]
port 574 nsew signal input
rlabel metal2 s 76930 0 76986 800 6 la_oenb[50]
port 575 nsew signal input
rlabel metal2 s 77850 0 77906 800 6 la_oenb[51]
port 576 nsew signal input
rlabel metal2 s 78770 0 78826 800 6 la_oenb[52]
port 577 nsew signal input
rlabel metal2 s 79598 0 79654 800 6 la_oenb[53]
port 578 nsew signal input
rlabel metal2 s 80518 0 80574 800 6 la_oenb[54]
port 579 nsew signal input
rlabel metal2 s 81438 0 81494 800 6 la_oenb[55]
port 580 nsew signal input
rlabel metal2 s 82358 0 82414 800 6 la_oenb[56]
port 581 nsew signal input
rlabel metal2 s 83186 0 83242 800 6 la_oenb[57]
port 582 nsew signal input
rlabel metal2 s 84106 0 84162 800 6 la_oenb[58]
port 583 nsew signal input
rlabel metal2 s 85026 0 85082 800 6 la_oenb[59]
port 584 nsew signal input
rlabel metal2 s 36726 0 36782 800 6 la_oenb[5]
port 585 nsew signal input
rlabel metal2 s 85854 0 85910 800 6 la_oenb[60]
port 586 nsew signal input
rlabel metal2 s 86774 0 86830 800 6 la_oenb[61]
port 587 nsew signal input
rlabel metal2 s 87694 0 87750 800 6 la_oenb[62]
port 588 nsew signal input
rlabel metal2 s 88614 0 88670 800 6 la_oenb[63]
port 589 nsew signal input
rlabel metal2 s 89442 0 89498 800 6 la_oenb[64]
port 590 nsew signal input
rlabel metal2 s 90362 0 90418 800 6 la_oenb[65]
port 591 nsew signal input
rlabel metal2 s 91282 0 91338 800 6 la_oenb[66]
port 592 nsew signal input
rlabel metal2 s 92110 0 92166 800 6 la_oenb[67]
port 593 nsew signal input
rlabel metal2 s 93030 0 93086 800 6 la_oenb[68]
port 594 nsew signal input
rlabel metal2 s 93950 0 94006 800 6 la_oenb[69]
port 595 nsew signal input
rlabel metal2 s 37646 0 37702 800 6 la_oenb[6]
port 596 nsew signal input
rlabel metal2 s 94870 0 94926 800 6 la_oenb[70]
port 597 nsew signal input
rlabel metal2 s 95698 0 95754 800 6 la_oenb[71]
port 598 nsew signal input
rlabel metal2 s 96618 0 96674 800 6 la_oenb[72]
port 599 nsew signal input
rlabel metal2 s 97538 0 97594 800 6 la_oenb[73]
port 600 nsew signal input
rlabel metal2 s 98366 0 98422 800 6 la_oenb[74]
port 601 nsew signal input
rlabel metal2 s 99286 0 99342 800 6 la_oenb[75]
port 602 nsew signal input
rlabel metal2 s 100206 0 100262 800 6 la_oenb[76]
port 603 nsew signal input
rlabel metal2 s 101126 0 101182 800 6 la_oenb[77]
port 604 nsew signal input
rlabel metal2 s 101954 0 102010 800 6 la_oenb[78]
port 605 nsew signal input
rlabel metal2 s 102874 0 102930 800 6 la_oenb[79]
port 606 nsew signal input
rlabel metal2 s 38474 0 38530 800 6 la_oenb[7]
port 607 nsew signal input
rlabel metal2 s 103794 0 103850 800 6 la_oenb[80]
port 608 nsew signal input
rlabel metal2 s 104622 0 104678 800 6 la_oenb[81]
port 609 nsew signal input
rlabel metal2 s 105542 0 105598 800 6 la_oenb[82]
port 610 nsew signal input
rlabel metal2 s 106462 0 106518 800 6 la_oenb[83]
port 611 nsew signal input
rlabel metal2 s 107382 0 107438 800 6 la_oenb[84]
port 612 nsew signal input
rlabel metal2 s 108210 0 108266 800 6 la_oenb[85]
port 613 nsew signal input
rlabel metal2 s 109130 0 109186 800 6 la_oenb[86]
port 614 nsew signal input
rlabel metal2 s 110050 0 110106 800 6 la_oenb[87]
port 615 nsew signal input
rlabel metal2 s 110878 0 110934 800 6 la_oenb[88]
port 616 nsew signal input
rlabel metal2 s 111798 0 111854 800 6 la_oenb[89]
port 617 nsew signal input
rlabel metal2 s 39394 0 39450 800 6 la_oenb[8]
port 618 nsew signal input
rlabel metal2 s 112718 0 112774 800 6 la_oenb[90]
port 619 nsew signal input
rlabel metal2 s 113638 0 113694 800 6 la_oenb[91]
port 620 nsew signal input
rlabel metal2 s 114466 0 114522 800 6 la_oenb[92]
port 621 nsew signal input
rlabel metal2 s 115386 0 115442 800 6 la_oenb[93]
port 622 nsew signal input
rlabel metal2 s 116306 0 116362 800 6 la_oenb[94]
port 623 nsew signal input
rlabel metal2 s 117134 0 117190 800 6 la_oenb[95]
port 624 nsew signal input
rlabel metal2 s 118054 0 118110 800 6 la_oenb[96]
port 625 nsew signal input
rlabel metal2 s 118974 0 119030 800 6 la_oenb[97]
port 626 nsew signal input
rlabel metal2 s 119894 0 119950 800 6 la_oenb[98]
port 627 nsew signal input
rlabel metal2 s 120722 0 120778 800 6 la_oenb[99]
port 628 nsew signal input
rlabel metal2 s 40314 0 40370 800 6 la_oenb[9]
port 629 nsew signal input
rlabel metal2 s 147586 0 147642 800 6 o_addr1[0]
port 630 nsew signal output
rlabel metal3 s 0 14560 800 14680 6 o_addr1[1]
port 631 nsew signal output
rlabel metal2 s 115478 165875 115534 166675 6 o_addr1[2]
port 632 nsew signal output
rlabel metal3 s 0 28024 800 28144 6 o_addr1[3]
port 633 nsew signal output
rlabel metal3 s 163731 36184 164531 36304 6 o_addr1[4]
port 634 nsew signal output
rlabel metal3 s 163731 41488 164531 41608 6 o_addr1[5]
port 635 nsew signal output
rlabel metal2 s 126886 165875 126942 166675 6 o_addr1[6]
port 636 nsew signal output
rlabel metal3 s 0 52232 800 52352 6 o_addr1[7]
port 637 nsew signal output
rlabel metal3 s 163731 60392 164531 60512 6 o_addr1[8]
port 638 nsew signal output
rlabel metal2 s 110694 165875 110750 166675 6 o_addr1_1[0]
port 639 nsew signal output
rlabel metal2 s 148782 0 148838 800 6 o_addr1_1[1]
port 640 nsew signal output
rlabel metal2 s 150254 0 150310 800 6 o_addr1_1[2]
port 641 nsew signal output
rlabel metal2 s 151450 0 151506 800 6 o_addr1_1[3]
port 642 nsew signal output
rlabel metal2 s 120262 165875 120318 166675 6 o_addr1_1[4]
port 643 nsew signal output
rlabel metal3 s 0 41488 800 41608 6 o_addr1_1[5]
port 644 nsew signal output
rlabel metal2 s 125966 165875 126022 166675 6 o_addr1_1[6]
port 645 nsew signal output
rlabel metal2 s 128818 165875 128874 166675 6 o_addr1_1[7]
port 646 nsew signal output
rlabel metal2 s 132590 165875 132646 166675 6 o_addr1_1[8]
port 647 nsew signal output
rlabel metal3 s 163731 1232 164531 1352 6 o_csb0
port 648 nsew signal output
rlabel metal2 s 108854 165875 108910 166675 6 o_csb0_1
port 649 nsew signal output
rlabel metal3 s 0 1232 800 1352 6 o_csb1
port 650 nsew signal output
rlabel metal3 s 0 3816 800 3936 6 o_csb1_1
port 651 nsew signal output
rlabel metal2 s 111706 165875 111762 166675 6 o_din0[0]
port 652 nsew signal output
rlabel metal3 s 0 68416 800 68536 6 o_din0[10]
port 653 nsew signal output
rlabel metal2 s 136362 165875 136418 166675 6 o_din0[11]
port 654 nsew signal output
rlabel metal2 s 139214 165875 139270 166675 6 o_din0[12]
port 655 nsew signal output
rlabel metal3 s 163731 92624 164531 92744 6 o_din0[13]
port 656 nsew signal output
rlabel metal3 s 0 87184 800 87304 6 o_din0[14]
port 657 nsew signal output
rlabel metal3 s 0 95344 800 95464 6 o_din0[15]
port 658 nsew signal output
rlabel metal2 s 157706 0 157762 800 6 o_din0[16]
port 659 nsew signal output
rlabel metal3 s 163731 116832 164531 116952 6 o_din0[17]
port 660 nsew signal output
rlabel metal2 s 158626 0 158682 800 6 o_din0[18]
port 661 nsew signal output
rlabel metal2 s 147770 165875 147826 166675 6 o_din0[19]
port 662 nsew signal output
rlabel metal3 s 163731 17280 164531 17400 6 o_din0[1]
port 663 nsew signal output
rlabel metal2 s 148782 165875 148838 166675 6 o_din0[20]
port 664 nsew signal output
rlabel metal3 s 163731 130296 164531 130416 6 o_din0[21]
port 665 nsew signal output
rlabel metal3 s 163731 135600 164531 135720 6 o_din0[22]
port 666 nsew signal output
rlabel metal3 s 0 127576 800 127696 6 o_din0[23]
port 667 nsew signal output
rlabel metal2 s 152554 165875 152610 166675 6 o_din0[24]
port 668 nsew signal output
rlabel metal3 s 0 141040 800 141160 6 o_din0[25]
port 669 nsew signal output
rlabel metal3 s 0 146344 800 146464 6 o_din0[26]
port 670 nsew signal output
rlabel metal3 s 0 149064 800 149184 6 o_din0[27]
port 671 nsew signal output
rlabel metal3 s 163731 154504 164531 154624 6 o_din0[28]
port 672 nsew signal output
rlabel metal2 s 163686 0 163742 800 6 o_din0[29]
port 673 nsew signal output
rlabel metal2 s 150530 0 150586 800 6 o_din0[2]
port 674 nsew signal output
rlabel metal2 s 164238 0 164294 800 6 o_din0[30]
port 675 nsew signal output
rlabel metal3 s 163731 165248 164531 165368 6 o_din0[31]
port 676 nsew signal output
rlabel metal3 s 163731 33464 164531 33584 6 o_din0[3]
port 677 nsew signal output
rlabel metal3 s 0 33464 800 33584 6 o_din0[4]
port 678 nsew signal output
rlabel metal2 s 122102 165875 122158 166675 6 o_din0[5]
port 679 nsew signal output
rlabel metal2 s 127806 165875 127862 166675 6 o_din0[6]
port 680 nsew signal output
rlabel metal3 s 0 54952 800 55072 6 o_din0[7]
port 681 nsew signal output
rlabel metal2 s 155958 0 156014 800 6 o_din0[8]
port 682 nsew signal output
rlabel metal3 s 163731 71136 164531 71256 6 o_din0[9]
port 683 nsew signal output
rlabel metal2 s 147862 0 147918 800 6 o_din0_1[0]
port 684 nsew signal output
rlabel metal3 s 163731 76440 164531 76560 6 o_din0_1[10]
port 685 nsew signal output
rlabel metal3 s 163731 87184 164531 87304 6 o_din0_1[11]
port 686 nsew signal output
rlabel metal2 s 138294 165875 138350 166675 6 o_din0_1[12]
port 687 nsew signal output
rlabel metal2 s 141146 165875 141202 166675 6 o_din0_1[13]
port 688 nsew signal output
rlabel metal3 s 0 84600 800 84720 6 o_din0_1[14]
port 689 nsew signal output
rlabel metal2 s 143078 165875 143134 166675 6 o_din0_1[15]
port 690 nsew signal output
rlabel metal3 s 163731 108672 164531 108792 6 o_din0_1[16]
port 691 nsew signal output
rlabel metal3 s 163731 114112 164531 114232 6 o_din0_1[17]
port 692 nsew signal output
rlabel metal2 s 145930 165875 145986 166675 6 o_din0_1[18]
port 693 nsew signal output
rlabel metal3 s 0 108672 800 108792 6 o_din0_1[19]
port 694 nsew signal output
rlabel metal3 s 0 17280 800 17400 6 o_din0_1[1]
port 695 nsew signal output
rlabel metal3 s 0 114112 800 114232 6 o_din0_1[20]
port 696 nsew signal output
rlabel metal3 s 0 119552 800 119672 6 o_din0_1[21]
port 697 nsew signal output
rlabel metal3 s 163731 132880 164531 133000 6 o_din0_1[22]
port 698 nsew signal output
rlabel metal2 s 161294 0 161350 800 6 o_din0_1[23]
port 699 nsew signal output
rlabel metal3 s 163731 143760 164531 143880 6 o_din0_1[24]
port 700 nsew signal output
rlabel metal2 s 154486 165875 154542 166675 6 o_din0_1[25]
port 701 nsew signal output
rlabel metal2 s 162214 0 162270 800 6 o_din0_1[26]
port 702 nsew signal output
rlabel metal2 s 157338 165875 157394 166675 6 o_din0_1[27]
port 703 nsew signal output
rlabel metal3 s 0 154504 800 154624 6 o_din0_1[28]
port 704 nsew signal output
rlabel metal2 s 161110 165875 161166 166675 6 o_din0_1[29]
port 705 nsew signal output
rlabel metal3 s 163731 22720 164531 22840 6 o_din0_1[2]
port 706 nsew signal output
rlabel metal3 s 0 159808 800 159928 6 o_din0_1[30]
port 707 nsew signal output
rlabel metal2 s 163962 165875 164018 166675 6 o_din0_1[31]
port 708 nsew signal output
rlabel metal2 s 151726 0 151782 800 6 o_din0_1[3]
port 709 nsew signal output
rlabel metal2 s 121182 165875 121238 166675 6 o_din0_1[4]
port 710 nsew signal output
rlabel metal2 s 154118 0 154174 800 6 o_din0_1[5]
port 711 nsew signal output
rlabel metal3 s 0 44208 800 44328 6 o_din0_1[6]
port 712 nsew signal output
rlabel metal2 s 129738 165875 129794 166675 6 o_din0_1[7]
port 713 nsew signal output
rlabel metal2 s 155590 0 155646 800 6 o_din0_1[8]
port 714 nsew signal output
rlabel metal3 s 0 65696 800 65816 6 o_din0_1[9]
port 715 nsew signal output
rlabel metal3 s 163731 6536 164531 6656 6 o_waddr0[0]
port 716 nsew signal output
rlabel metal3 s 163731 20000 164531 20120 6 o_waddr0[1]
port 717 nsew signal output
rlabel metal3 s 163731 25304 164531 25424 6 o_waddr0[2]
port 718 nsew signal output
rlabel metal2 s 152002 0 152058 800 6 o_waddr0[3]
port 719 nsew signal output
rlabel metal3 s 0 38768 800 38888 6 o_waddr0[4]
port 720 nsew signal output
rlabel metal2 s 124034 165875 124090 166675 6 o_waddr0[5]
port 721 nsew signal output
rlabel metal2 s 154762 0 154818 800 6 o_waddr0[6]
port 722 nsew signal output
rlabel metal3 s 163731 54952 164531 55072 6 o_waddr0[7]
port 723 nsew signal output
rlabel metal3 s 0 60392 800 60512 6 o_waddr0[8]
port 724 nsew signal output
rlabel metal3 s 0 11976 800 12096 6 o_waddr0_1[0]
port 725 nsew signal output
rlabel metal2 s 113546 165875 113602 166675 6 o_waddr0_1[1]
port 726 nsew signal output
rlabel metal2 s 150898 0 150954 800 6 o_waddr0_1[2]
port 727 nsew signal output
rlabel metal2 s 117410 165875 117466 166675 6 o_waddr0_1[3]
port 728 nsew signal output
rlabel metal3 s 0 36184 800 36304 6 o_waddr0_1[4]
port 729 nsew signal output
rlabel metal2 s 123114 165875 123170 166675 6 o_waddr0_1[5]
port 730 nsew signal output
rlabel metal3 s 163731 49512 164531 49632 6 o_waddr0_1[6]
port 731 nsew signal output
rlabel metal2 s 155314 0 155370 800 6 o_waddr0_1[7]
port 732 nsew signal output
rlabel metal3 s 163731 62976 164531 63096 6 o_waddr0_1[8]
port 733 nsew signal output
rlabel metal2 s 109774 165875 109830 166675 6 o_web0
port 734 nsew signal output
rlabel metal3 s 163731 3816 164531 3936 6 o_web0_1
port 735 nsew signal output
rlabel metal3 s 163731 9256 164531 9376 6 o_wmask0[0]
port 736 nsew signal output
rlabel metal2 s 149334 0 149390 800 6 o_wmask0[1]
port 737 nsew signal output
rlabel metal3 s 163731 28024 164531 28144 6 o_wmask0[2]
port 738 nsew signal output
rlabel metal2 s 152370 0 152426 800 6 o_wmask0[3]
port 739 nsew signal output
rlabel metal2 s 112626 165875 112682 166675 6 o_wmask0_1[0]
port 740 nsew signal output
rlabel metal2 s 149058 0 149114 800 6 o_wmask0_1[1]
port 741 nsew signal output
rlabel metal3 s 0 22720 800 22840 6 o_wmask0_1[2]
port 742 nsew signal output
rlabel metal2 s 118330 165875 118386 166675 6 o_wmask0_1[3]
port 743 nsew signal output
rlabel metal4 s 4208 2128 4528 164336 6 vccd1
port 744 nsew power input
rlabel metal4 s 34928 2128 35248 164336 6 vccd1
port 744 nsew power input
rlabel metal4 s 65648 2128 65968 164336 6 vccd1
port 744 nsew power input
rlabel metal4 s 96368 2128 96688 164336 6 vccd1
port 744 nsew power input
rlabel metal4 s 127088 2128 127408 164336 6 vccd1
port 744 nsew power input
rlabel metal4 s 157808 2128 158128 164336 6 vccd1
port 744 nsew power input
rlabel metal4 s 19568 2128 19888 164336 6 vssd1
port 745 nsew ground input
rlabel metal4 s 50288 2128 50608 164336 6 vssd1
port 745 nsew ground input
rlabel metal4 s 81008 2128 81328 164336 6 vssd1
port 745 nsew ground input
rlabel metal4 s 111728 2128 112048 164336 6 vssd1
port 745 nsew ground input
rlabel metal4 s 142448 2128 142768 164336 6 vssd1
port 745 nsew ground input
rlabel metal2 s 110 0 166 800 6 wb_clk_i
port 746 nsew signal input
rlabel metal2 s 386 0 442 800 6 wb_rst_i
port 747 nsew signal input
rlabel metal2 s 662 0 718 800 6 wbs_ack_o
port 748 nsew signal output
rlabel metal2 s 1858 0 1914 800 6 wbs_adr_i[0]
port 749 nsew signal input
rlabel metal2 s 11978 0 12034 800 6 wbs_adr_i[10]
port 750 nsew signal input
rlabel metal2 s 12898 0 12954 800 6 wbs_adr_i[11]
port 751 nsew signal input
rlabel metal2 s 13818 0 13874 800 6 wbs_adr_i[12]
port 752 nsew signal input
rlabel metal2 s 14646 0 14702 800 6 wbs_adr_i[13]
port 753 nsew signal input
rlabel metal2 s 15566 0 15622 800 6 wbs_adr_i[14]
port 754 nsew signal input
rlabel metal2 s 16486 0 16542 800 6 wbs_adr_i[15]
port 755 nsew signal input
rlabel metal2 s 17314 0 17370 800 6 wbs_adr_i[16]
port 756 nsew signal input
rlabel metal2 s 18234 0 18290 800 6 wbs_adr_i[17]
port 757 nsew signal input
rlabel metal2 s 19154 0 19210 800 6 wbs_adr_i[18]
port 758 nsew signal input
rlabel metal2 s 20074 0 20130 800 6 wbs_adr_i[19]
port 759 nsew signal input
rlabel metal2 s 3054 0 3110 800 6 wbs_adr_i[1]
port 760 nsew signal input
rlabel metal2 s 20902 0 20958 800 6 wbs_adr_i[20]
port 761 nsew signal input
rlabel metal2 s 21822 0 21878 800 6 wbs_adr_i[21]
port 762 nsew signal input
rlabel metal2 s 22742 0 22798 800 6 wbs_adr_i[22]
port 763 nsew signal input
rlabel metal2 s 23570 0 23626 800 6 wbs_adr_i[23]
port 764 nsew signal input
rlabel metal2 s 24490 0 24546 800 6 wbs_adr_i[24]
port 765 nsew signal input
rlabel metal2 s 25410 0 25466 800 6 wbs_adr_i[25]
port 766 nsew signal input
rlabel metal2 s 26330 0 26386 800 6 wbs_adr_i[26]
port 767 nsew signal input
rlabel metal2 s 27158 0 27214 800 6 wbs_adr_i[27]
port 768 nsew signal input
rlabel metal2 s 28078 0 28134 800 6 wbs_adr_i[28]
port 769 nsew signal input
rlabel metal2 s 28998 0 29054 800 6 wbs_adr_i[29]
port 770 nsew signal input
rlabel metal2 s 4250 0 4306 800 6 wbs_adr_i[2]
port 771 nsew signal input
rlabel metal2 s 29826 0 29882 800 6 wbs_adr_i[30]
port 772 nsew signal input
rlabel metal2 s 30746 0 30802 800 6 wbs_adr_i[31]
port 773 nsew signal input
rlabel metal2 s 5446 0 5502 800 6 wbs_adr_i[3]
port 774 nsew signal input
rlabel metal2 s 6642 0 6698 800 6 wbs_adr_i[4]
port 775 nsew signal input
rlabel metal2 s 7470 0 7526 800 6 wbs_adr_i[5]
port 776 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 wbs_adr_i[6]
port 777 nsew signal input
rlabel metal2 s 9310 0 9366 800 6 wbs_adr_i[7]
port 778 nsew signal input
rlabel metal2 s 10230 0 10286 800 6 wbs_adr_i[8]
port 779 nsew signal input
rlabel metal2 s 11058 0 11114 800 6 wbs_adr_i[9]
port 780 nsew signal input
rlabel metal2 s 938 0 994 800 6 wbs_cyc_i
port 781 nsew signal input
rlabel metal2 s 2134 0 2190 800 6 wbs_dat_i[0]
port 782 nsew signal input
rlabel metal2 s 12254 0 12310 800 6 wbs_dat_i[10]
port 783 nsew signal input
rlabel metal2 s 13174 0 13230 800 6 wbs_dat_i[11]
port 784 nsew signal input
rlabel metal2 s 14094 0 14150 800 6 wbs_dat_i[12]
port 785 nsew signal input
rlabel metal2 s 14922 0 14978 800 6 wbs_dat_i[13]
port 786 nsew signal input
rlabel metal2 s 15842 0 15898 800 6 wbs_dat_i[14]
port 787 nsew signal input
rlabel metal2 s 16762 0 16818 800 6 wbs_dat_i[15]
port 788 nsew signal input
rlabel metal2 s 17682 0 17738 800 6 wbs_dat_i[16]
port 789 nsew signal input
rlabel metal2 s 18510 0 18566 800 6 wbs_dat_i[17]
port 790 nsew signal input
rlabel metal2 s 19430 0 19486 800 6 wbs_dat_i[18]
port 791 nsew signal input
rlabel metal2 s 20350 0 20406 800 6 wbs_dat_i[19]
port 792 nsew signal input
rlabel metal2 s 3330 0 3386 800 6 wbs_dat_i[1]
port 793 nsew signal input
rlabel metal2 s 21178 0 21234 800 6 wbs_dat_i[20]
port 794 nsew signal input
rlabel metal2 s 22098 0 22154 800 6 wbs_dat_i[21]
port 795 nsew signal input
rlabel metal2 s 23018 0 23074 800 6 wbs_dat_i[22]
port 796 nsew signal input
rlabel metal2 s 23938 0 23994 800 6 wbs_dat_i[23]
port 797 nsew signal input
rlabel metal2 s 24766 0 24822 800 6 wbs_dat_i[24]
port 798 nsew signal input
rlabel metal2 s 25686 0 25742 800 6 wbs_dat_i[25]
port 799 nsew signal input
rlabel metal2 s 26606 0 26662 800 6 wbs_dat_i[26]
port 800 nsew signal input
rlabel metal2 s 27526 0 27582 800 6 wbs_dat_i[27]
port 801 nsew signal input
rlabel metal2 s 28354 0 28410 800 6 wbs_dat_i[28]
port 802 nsew signal input
rlabel metal2 s 29274 0 29330 800 6 wbs_dat_i[29]
port 803 nsew signal input
rlabel metal2 s 4526 0 4582 800 6 wbs_dat_i[2]
port 804 nsew signal input
rlabel metal2 s 30194 0 30250 800 6 wbs_dat_i[30]
port 805 nsew signal input
rlabel metal2 s 31022 0 31078 800 6 wbs_dat_i[31]
port 806 nsew signal input
rlabel metal2 s 5722 0 5778 800 6 wbs_dat_i[3]
port 807 nsew signal input
rlabel metal2 s 6918 0 6974 800 6 wbs_dat_i[4]
port 808 nsew signal input
rlabel metal2 s 7838 0 7894 800 6 wbs_dat_i[5]
port 809 nsew signal input
rlabel metal2 s 8666 0 8722 800 6 wbs_dat_i[6]
port 810 nsew signal input
rlabel metal2 s 9586 0 9642 800 6 wbs_dat_i[7]
port 811 nsew signal input
rlabel metal2 s 10506 0 10562 800 6 wbs_dat_i[8]
port 812 nsew signal input
rlabel metal2 s 11426 0 11482 800 6 wbs_dat_i[9]
port 813 nsew signal input
rlabel metal2 s 2410 0 2466 800 6 wbs_dat_o[0]
port 814 nsew signal output
rlabel metal2 s 12622 0 12678 800 6 wbs_dat_o[10]
port 815 nsew signal output
rlabel metal2 s 13450 0 13506 800 6 wbs_dat_o[11]
port 816 nsew signal output
rlabel metal2 s 14370 0 14426 800 6 wbs_dat_o[12]
port 817 nsew signal output
rlabel metal2 s 15290 0 15346 800 6 wbs_dat_o[13]
port 818 nsew signal output
rlabel metal2 s 16118 0 16174 800 6 wbs_dat_o[14]
port 819 nsew signal output
rlabel metal2 s 17038 0 17094 800 6 wbs_dat_o[15]
port 820 nsew signal output
rlabel metal2 s 17958 0 18014 800 6 wbs_dat_o[16]
port 821 nsew signal output
rlabel metal2 s 18878 0 18934 800 6 wbs_dat_o[17]
port 822 nsew signal output
rlabel metal2 s 19706 0 19762 800 6 wbs_dat_o[18]
port 823 nsew signal output
rlabel metal2 s 20626 0 20682 800 6 wbs_dat_o[19]
port 824 nsew signal output
rlabel metal2 s 3606 0 3662 800 6 wbs_dat_o[1]
port 825 nsew signal output
rlabel metal2 s 21546 0 21602 800 6 wbs_dat_o[20]
port 826 nsew signal output
rlabel metal2 s 22374 0 22430 800 6 wbs_dat_o[21]
port 827 nsew signal output
rlabel metal2 s 23294 0 23350 800 6 wbs_dat_o[22]
port 828 nsew signal output
rlabel metal2 s 24214 0 24270 800 6 wbs_dat_o[23]
port 829 nsew signal output
rlabel metal2 s 25134 0 25190 800 6 wbs_dat_o[24]
port 830 nsew signal output
rlabel metal2 s 25962 0 26018 800 6 wbs_dat_o[25]
port 831 nsew signal output
rlabel metal2 s 26882 0 26938 800 6 wbs_dat_o[26]
port 832 nsew signal output
rlabel metal2 s 27802 0 27858 800 6 wbs_dat_o[27]
port 833 nsew signal output
rlabel metal2 s 28630 0 28686 800 6 wbs_dat_o[28]
port 834 nsew signal output
rlabel metal2 s 29550 0 29606 800 6 wbs_dat_o[29]
port 835 nsew signal output
rlabel metal2 s 4802 0 4858 800 6 wbs_dat_o[2]
port 836 nsew signal output
rlabel metal2 s 30470 0 30526 800 6 wbs_dat_o[30]
port 837 nsew signal output
rlabel metal2 s 31390 0 31446 800 6 wbs_dat_o[31]
port 838 nsew signal output
rlabel metal2 s 5998 0 6054 800 6 wbs_dat_o[3]
port 839 nsew signal output
rlabel metal2 s 7194 0 7250 800 6 wbs_dat_o[4]
port 840 nsew signal output
rlabel metal2 s 8114 0 8170 800 6 wbs_dat_o[5]
port 841 nsew signal output
rlabel metal2 s 9034 0 9090 800 6 wbs_dat_o[6]
port 842 nsew signal output
rlabel metal2 s 9862 0 9918 800 6 wbs_dat_o[7]
port 843 nsew signal output
rlabel metal2 s 10782 0 10838 800 6 wbs_dat_o[8]
port 844 nsew signal output
rlabel metal2 s 11702 0 11758 800 6 wbs_dat_o[9]
port 845 nsew signal output
rlabel metal2 s 2778 0 2834 800 6 wbs_sel_i[0]
port 846 nsew signal input
rlabel metal2 s 3974 0 4030 800 6 wbs_sel_i[1]
port 847 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 wbs_sel_i[2]
port 848 nsew signal input
rlabel metal2 s 6366 0 6422 800 6 wbs_sel_i[3]
port 849 nsew signal input
rlabel metal2 s 1214 0 1270 800 6 wbs_stb_i
port 850 nsew signal input
rlabel metal2 s 1582 0 1638 800 6 wbs_we_i
port 851 nsew signal input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 164531 166675
string LEFview TRUE
string GDS_FILE /local/caravel_user_project/openlane/user_proj/runs/user_proj/results/magic/user_proj.gds
string GDS_END 79185436
string GDS_START 1368802
<< end >>

