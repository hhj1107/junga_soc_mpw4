VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_proj
  CLASS BLOCK ;
  FOREIGN user_proj ;
  ORIGIN 0.000 0.000 ;
  SIZE 823.900 BY 834.620 ;
  PIN i_dout0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 20.440 823.900 21.040 ;
    END
  END i_dout0[0]
  PIN i_dout0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.070 830.620 673.350 834.620 ;
    END
  END i_dout0[10]
  PIN i_dout0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 361.800 823.900 362.400 ;
    END
  END i_dout0[11]
  PIN i_dout0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 438.640 4.000 439.240 ;
    END
  END i_dout0[12]
  PIN i_dout0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 416.880 823.900 417.480 ;
    END
  END i_dout0[13]
  PIN i_dout0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 444.080 823.900 444.680 ;
    END
  END i_dout0[14]
  PIN i_dout0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 712.630 830.620 712.910 834.620 ;
    END
  END i_dout0[15]
  PIN i_dout0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 732.410 830.620 732.690 834.620 ;
    END
  END i_dout0[16]
  PIN i_dout0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 485.560 823.900 486.160 ;
    END
  END i_dout0[17]
  PIN i_dout0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 742.070 830.620 742.350 834.620 ;
    END
  END i_dout0[18]
  PIN i_dout0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 512.760 823.900 513.360 ;
    END
  END i_dout0[19]
  PIN i_dout0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.000 4.000 66.600 ;
    END
  END i_dout0[1]
  PIN i_dout0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 526.360 823.900 526.960 ;
    END
  END i_dout0[20]
  PIN i_dout0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 587.560 4.000 588.160 ;
    END
  END i_dout0[21]
  PIN i_dout0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 771.970 830.620 772.250 834.620 ;
    END
  END i_dout0[22]
  PIN i_dout0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 806.470 0.000 806.750 4.000 ;
    END
  END i_dout0[23]
  PIN i_dout0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 647.400 4.000 648.000 ;
    END
  END i_dout0[24]
  PIN i_dout0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 676.640 4.000 677.240 ;
    END
  END i_dout0[25]
  PIN i_dout0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 815.210 0.000 815.490 4.000 ;
    END
  END i_dout0[26]
  PIN i_dout0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 736.480 4.000 737.080 ;
    END
  END i_dout0[27]
  PIN i_dout0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 818.430 0.000 818.710 4.000 ;
    END
  END i_dout0[28]
  PIN i_dout0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 745.320 823.900 745.920 ;
    END
  END i_dout0[29]
  PIN i_dout0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 88.440 823.900 89.040 ;
    END
  END i_dout0[2]
  PIN i_dout0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 821.190 0.000 821.470 4.000 ;
    END
  END i_dout0[30]
  PIN i_dout0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 799.720 823.900 800.320 ;
    END
  END i_dout0[31]
  PIN i_dout0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 143.520 823.900 144.120 ;
    END
  END i_dout0[3]
  PIN i_dout0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.920 4.000 215.520 ;
    END
  END i_dout0[4]
  PIN i_dout0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 748.510 0.000 748.790 4.000 ;
    END
  END i_dout0[5]
  PIN i_dout0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 755.870 0.000 756.150 4.000 ;
    END
  END i_dout0[6]
  PIN i_dout0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 761.390 0.000 761.670 4.000 ;
    END
  END i_dout0[7]
  PIN i_dout0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 767.370 0.000 767.650 4.000 ;
    END
  END i_dout0[8]
  PIN i_dout0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 663.410 830.620 663.690 834.620 ;
    END
  END i_dout0[9]
  PIN i_dout0_1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 722.290 0.000 722.570 4.000 ;
    END
  END i_dout0_1[0]
  PIN i_dout0_1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 321.000 823.900 321.600 ;
    END
  END i_dout0_1[10]
  PIN i_dout0_1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 682.730 830.620 683.010 834.620 ;
    END
  END i_dout0_1[11]
  PIN i_dout0_1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 777.490 0.000 777.770 4.000 ;
    END
  END i_dout0_1[12]
  PIN i_dout0_1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 453.600 4.000 454.200 ;
    END
  END i_dout0_1[13]
  PIN i_dout0_1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 697.910 830.620 698.190 834.620 ;
    END
  END i_dout0_1[14]
  PIN i_dout0_1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 707.570 830.620 707.850 834.620 ;
    END
  END i_dout0_1[15]
  PIN i_dout0_1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 727.350 830.620 727.630 834.620 ;
    END
  END i_dout0_1[16]
  PIN i_dout0_1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 498.480 4.000 499.080 ;
    END
  END i_dout0_1[17]
  PIN i_dout0_1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 499.160 823.900 499.760 ;
    END
  END i_dout0_1[18]
  PIN i_dout0_1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 542.680 4.000 543.280 ;
    END
  END i_dout0_1[19]
  PIN i_dout0_1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 61.240 823.900 61.840 ;
    END
  END i_dout0_1[1]
  PIN i_dout0_1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 799.570 0.000 799.850 4.000 ;
    END
  END i_dout0_1[20]
  PIN i_dout0_1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 766.910 830.620 767.190 834.620 ;
    END
  END i_dout0_1[21]
  PIN i_dout0_1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 803.710 0.000 803.990 4.000 ;
    END
  END i_dout0_1[22]
  PIN i_dout0_1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 617.480 4.000 618.080 ;
    END
  END i_dout0_1[23]
  PIN i_dout0_1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 811.070 0.000 811.350 4.000 ;
    END
  END i_dout0_1[24]
  PIN i_dout0_1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 786.690 830.620 786.970 834.620 ;
    END
  END i_dout0_1[25]
  PIN i_dout0_1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 791.290 830.620 791.570 834.620 ;
    END
  END i_dout0_1[26]
  PIN i_dout0_1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 796.350 830.620 796.630 834.620 ;
    END
  END i_dout0_1[27]
  PIN i_dout0_1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 806.470 830.620 806.750 834.620 ;
    END
  END i_dout0_1[28]
  PIN i_dout0_1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 731.720 823.900 732.320 ;
    END
  END i_dout0_1[29]
  PIN i_dout0_1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 589.350 830.620 589.630 834.620 ;
    END
  END i_dout0_1[2]
  PIN i_dout0_1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 819.810 0.000 820.090 4.000 ;
    END
  END i_dout0_1[30]
  PIN i_dout0_1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 811.280 4.000 811.880 ;
    END
  END i_dout0_1[31]
  PIN i_dout0_1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 129.920 823.900 130.520 ;
    END
  END i_dout0_1[3]
  PIN i_dout0_1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 743.910 0.000 744.190 4.000 ;
    END
  END i_dout0_1[4]
  PIN i_dout0_1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 225.120 823.900 225.720 ;
    END
  END i_dout0_1[5]
  PIN i_dout0_1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 628.910 830.620 629.190 834.620 ;
    END
  END i_dout0_1[6]
  PIN i_dout0_1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.010 0.000 760.290 4.000 ;
    END
  END i_dout0_1[7]
  PIN i_dout0_1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 765.990 0.000 766.270 4.000 ;
    END
  END i_dout0_1[8]
  PIN i_dout0_1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 307.400 823.900 308.000 ;
    END
  END i_dout0_1[9]
  PIN i_dout1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 723.670 0.000 723.950 4.000 ;
    END
  END i_dout1[0]
  PIN i_dout1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 334.600 823.900 335.200 ;
    END
  END i_dout1[10]
  PIN i_dout1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 376.080 823.900 376.680 ;
    END
  END i_dout1[11]
  PIN i_dout1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 389.680 823.900 390.280 ;
    END
  END i_dout1[12]
  PIN i_dout1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 780.250 0.000 780.530 4.000 ;
    END
  END i_dout1[13]
  PIN i_dout1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 457.680 823.900 458.280 ;
    END
  END i_dout1[14]
  PIN i_dout1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 717.690 830.620 717.970 834.620 ;
    END
  END i_dout1[15]
  PIN i_dout1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 786.230 0.000 786.510 4.000 ;
    END
  END i_dout1[16]
  PIN i_dout1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 512.760 4.000 513.360 ;
    END
  END i_dout1[17]
  PIN i_dout1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 794.970 0.000 795.250 4.000 ;
    END
  END i_dout1[18]
  PIN i_dout1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 752.190 830.620 752.470 834.620 ;
    END
  END i_dout1[19]
  PIN i_dout1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 74.840 823.900 75.440 ;
    END
  END i_dout1[1]
  PIN i_dout1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 539.960 823.900 540.560 ;
    END
  END i_dout1[20]
  PIN i_dout1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 802.330 0.000 802.610 4.000 ;
    END
  END i_dout1[21]
  PIN i_dout1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 580.760 823.900 581.360 ;
    END
  END i_dout1[22]
  PIN i_dout1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 632.440 4.000 633.040 ;
    END
  END i_dout1[23]
  PIN i_dout1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 812.450 0.000 812.730 4.000 ;
    END
  END i_dout1[24]
  PIN i_dout1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 635.840 823.900 636.440 ;
    END
  END i_dout1[25]
  PIN i_dout1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 817.050 0.000 817.330 4.000 ;
    END
  END i_dout1[26]
  PIN i_dout1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 751.440 4.000 752.040 ;
    END
  END i_dout1[27]
  PIN i_dout1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 703.840 823.900 704.440 ;
    END
  END i_dout1[28]
  PIN i_dout1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 766.400 4.000 767.000 ;
    END
  END i_dout1[29]
  PIN i_dout1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.920 4.000 96.520 ;
    END
  END i_dout1[2]
  PIN i_dout1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 781.360 4.000 781.960 ;
    END
  END i_dout1[30]
  PIN i_dout1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 813.320 823.900 813.920 ;
    END
  END i_dout1[31]
  PIN i_dout1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.010 830.620 599.290 834.620 ;
    END
  END i_dout1[3]
  PIN i_dout1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 618.790 830.620 619.070 834.620 ;
    END
  END i_dout1[4]
  PIN i_dout1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 749.890 0.000 750.170 4.000 ;
    END
  END i_dout1[5]
  PIN i_dout1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 757.250 0.000 757.530 4.000 ;
    END
  END i_dout1[6]
  PIN i_dout1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 266.600 823.900 267.200 ;
    END
  END i_dout1[7]
  PIN i_dout1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 768.750 0.000 769.030 4.000 ;
    END
  END i_dout1[8]
  PIN i_dout1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 378.800 4.000 379.400 ;
    END
  END i_dout1[9]
  PIN i_dout1_1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 34.040 823.900 34.640 ;
    END
  END i_dout1_1[0]
  PIN i_dout1_1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 774.730 0.000 775.010 4.000 ;
    END
  END i_dout1_1[10]
  PIN i_dout1_1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 408.720 4.000 409.320 ;
    END
  END i_dout1_1[11]
  PIN i_dout1_1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 423.680 4.000 424.280 ;
    END
  END i_dout1_1[12]
  PIN i_dout1_1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 778.870 0.000 779.150 4.000 ;
    END
  END i_dout1_1[13]
  PIN i_dout1_1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 430.480 823.900 431.080 ;
    END
  END i_dout1_1[14]
  PIN i_dout1_1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 784.850 0.000 785.130 4.000 ;
    END
  END i_dout1_1[15]
  PIN i_dout1_1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 471.280 823.900 471.880 ;
    END
  END i_dout1_1[16]
  PIN i_dout1_1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 790.830 0.000 791.110 4.000 ;
    END
  END i_dout1_1[17]
  PIN i_dout1_1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 793.590 0.000 793.870 4.000 ;
    END
  END i_dout1_1[18]
  PIN i_dout1_1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 796.350 0.000 796.630 4.000 ;
    END
  END i_dout1_1[19]
  PIN i_dout1_1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 729.190 0.000 729.470 4.000 ;
    END
  END i_dout1_1[1]
  PIN i_dout1_1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 800.950 0.000 801.230 4.000 ;
    END
  END i_dout1_1[20]
  PIN i_dout1_1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 572.600 4.000 573.200 ;
    END
  END i_dout1_1[21]
  PIN i_dout1_1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 602.520 4.000 603.120 ;
    END
  END i_dout1_1[22]
  PIN i_dout1_1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 608.640 823.900 609.240 ;
    END
  END i_dout1_1[23]
  PIN i_dout1_1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 776.570 830.620 776.850 834.620 ;
    END
  END i_dout1_1[24]
  PIN i_dout1_1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 662.360 4.000 662.960 ;
    END
  END i_dout1_1[25]
  PIN i_dout1_1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 663.040 823.900 663.640 ;
    END
  END i_dout1_1[26]
  PIN i_dout1_1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 721.520 4.000 722.120 ;
    END
  END i_dout1_1[27]
  PIN i_dout1_1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 690.240 823.900 690.840 ;
    END
  END i_dout1_1[28]
  PIN i_dout1_1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 816.130 830.620 816.410 834.620 ;
    END
  END i_dout1_1[29]
  PIN i_dout1_1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.930 0.000 738.210 4.000 ;
    END
  END i_dout1_1[2]
  PIN i_dout1_1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 772.520 823.900 773.120 ;
    END
  END i_dout1_1[30]
  PIN i_dout1_1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 822.570 0.000 822.850 4.000 ;
    END
  END i_dout1_1[31]
  PIN i_dout1_1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 741.150 0.000 741.430 4.000 ;
    END
  END i_dout1_1[3]
  PIN i_dout1_1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 613.730 830.620 614.010 834.620 ;
    END
  END i_dout1_1[4]
  PIN i_dout1_1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 623.850 830.620 624.130 834.620 ;
    END
  END i_dout1_1[5]
  PIN i_dout1_1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 754.030 0.000 754.310 4.000 ;
    END
  END i_dout1_1[6]
  PIN i_dout1_1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 319.640 4.000 320.240 ;
    END
  END i_dout1_1[7]
  PIN i_dout1_1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 334.600 4.000 335.200 ;
    END
  END i_dout1_1[8]
  PIN i_dout1_1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 773.350 0.000 773.630 4.000 ;
    END
  END i_dout1_1[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.390 830.620 2.670 834.620 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.050 830.620 150.330 834.620 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.770 830.620 165.050 834.620 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.950 830.620 180.230 834.620 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.670 830.620 194.950 834.620 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.390 830.620 209.670 834.620 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.110 830.620 224.390 834.620 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.830 830.620 239.110 834.620 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.550 830.620 253.830 834.620 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.730 830.620 269.010 834.620 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.450 830.620 283.730 834.620 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.110 830.620 17.390 834.620 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.170 830.620 298.450 834.620 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.890 830.620 313.170 834.620 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.610 830.620 327.890 834.620 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.330 830.620 342.610 834.620 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.510 830.620 357.790 834.620 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 372.230 830.620 372.510 834.620 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.950 830.620 387.230 834.620 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 401.670 830.620 401.950 834.620 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.390 830.620 416.670 834.620 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.570 830.620 431.850 834.620 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.830 830.620 32.110 834.620 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 446.290 830.620 446.570 834.620 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.010 830.620 461.290 834.620 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 475.730 830.620 476.010 834.620 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 490.450 830.620 490.730 834.620 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.170 830.620 505.450 834.620 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 520.350 830.620 520.630 834.620 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 535.070 830.620 535.350 834.620 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 549.790 830.620 550.070 834.620 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.550 830.620 46.830 834.620 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 830.620 61.550 834.620 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.990 830.620 76.270 834.620 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.170 830.620 91.450 834.620 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.890 830.620 106.170 834.620 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.610 830.620 120.890 834.620 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 830.620 135.610 834.620 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 830.620 7.270 834.620 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.110 830.620 155.390 834.620 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.830 830.620 170.110 834.620 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.550 830.620 184.830 834.620 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.270 830.620 199.550 834.620 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.450 830.620 214.730 834.620 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.170 830.620 229.450 834.620 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.890 830.620 244.170 834.620 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.610 830.620 258.890 834.620 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.330 830.620 273.610 834.620 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.510 830.620 288.790 834.620 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.710 830.620 21.990 834.620 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.230 830.620 303.510 834.620 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.950 830.620 318.230 834.620 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.670 830.620 332.950 834.620 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.390 830.620 347.670 834.620 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.110 830.620 362.390 834.620 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.290 830.620 377.570 834.620 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.010 830.620 392.290 834.620 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 406.730 830.620 407.010 834.620 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.450 830.620 421.730 834.620 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 436.170 830.620 436.450 834.620 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.890 830.620 37.170 834.620 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.890 830.620 451.170 834.620 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.070 830.620 466.350 834.620 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 480.790 830.620 481.070 834.620 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.510 830.620 495.790 834.620 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 510.230 830.620 510.510 834.620 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.950 830.620 525.230 834.620 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 539.670 830.620 539.950 834.620 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 554.850 830.620 555.130 834.620 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 830.620 51.890 834.620 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.330 830.620 66.610 834.620 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.050 830.620 81.330 834.620 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.770 830.620 96.050 834.620 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.490 830.620 110.770 834.620 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 830.620 125.950 834.620 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.390 830.620 140.670 834.620 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.050 830.620 12.330 834.620 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.170 830.620 160.450 834.620 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.890 830.620 175.170 834.620 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.610 830.620 189.890 834.620 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.330 830.620 204.610 834.620 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 830.620 219.330 834.620 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.230 830.620 234.510 834.620 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.950 830.620 249.230 834.620 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.670 830.620 263.950 834.620 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.390 830.620 278.670 834.620 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.110 830.620 293.390 834.620 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.770 830.620 27.050 834.620 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 307.830 830.620 308.110 834.620 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.010 830.620 323.290 834.620 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.730 830.620 338.010 834.620 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.450 830.620 352.730 834.620 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.170 830.620 367.450 834.620 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 381.890 830.620 382.170 834.620 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.610 830.620 396.890 834.620 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 411.790 830.620 412.070 834.620 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 426.510 830.620 426.790 834.620 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.230 830.620 441.510 834.620 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.490 830.620 41.770 834.620 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.950 830.620 456.230 834.620 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.670 830.620 470.950 834.620 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 485.850 830.620 486.130 834.620 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 500.570 830.620 500.850 834.620 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 515.290 830.620 515.570 834.620 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 530.010 830.620 530.290 834.620 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.730 830.620 545.010 834.620 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 559.450 830.620 559.730 834.620 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.210 830.620 56.490 834.620 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.390 830.620 71.670 834.620 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.110 830.620 86.390 834.620 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.830 830.620 101.110 834.620 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.550 830.620 115.830 834.620 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.270 830.620 130.550 834.620 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.450 830.620 145.730 834.620 ;
    END
  END io_out[9]
  PIN irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 714.930 0.000 715.210 4.000 ;
    END
  END irq[0]
  PIN irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 716.310 0.000 716.590 4.000 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 717.690 0.000 717.970 4.000 ;
    END
  END irq[2]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.110 0.000 155.390 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 592.110 0.000 592.390 4.000 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 596.710 0.000 596.990 4.000 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 601.310 0.000 601.590 4.000 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.450 0.000 605.730 4.000 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 610.050 0.000 610.330 4.000 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 614.190 0.000 614.470 4.000 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 618.790 0.000 619.070 4.000 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 622.930 0.000 623.210 4.000 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.530 0.000 627.810 4.000 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 631.670 0.000 631.950 4.000 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.810 0.000 199.090 4.000 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 636.270 0.000 636.550 4.000 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 640.410 0.000 640.690 4.000 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 645.010 0.000 645.290 4.000 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 649.150 0.000 649.430 4.000 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 653.750 0.000 654.030 4.000 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 657.890 0.000 658.170 4.000 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 662.490 0.000 662.770 4.000 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 666.630 0.000 666.910 4.000 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 671.230 0.000 671.510 4.000 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 675.370 0.000 675.650 4.000 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 0.000 203.230 4.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 679.970 0.000 680.250 4.000 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 684.110 0.000 684.390 4.000 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 688.710 0.000 688.990 4.000 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 692.850 0.000 693.130 4.000 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 697.450 0.000 697.730 4.000 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 701.590 0.000 701.870 4.000 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 706.190 0.000 706.470 4.000 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 710.330 0.000 710.610 4.000 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.550 0.000 207.830 4.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.690 0.000 211.970 4.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.290 0.000 216.570 4.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.430 0.000 220.710 4.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.030 0.000 225.310 4.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.170 0.000 229.450 4.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.770 0.000 234.050 4.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.910 0.000 238.190 4.000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.250 0.000 159.530 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.510 0.000 242.790 4.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.650 0.000 246.930 4.000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.250 0.000 251.530 4.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.390 0.000 255.670 4.000 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.990 0.000 260.270 4.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.130 0.000 264.410 4.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.730 0.000 269.010 4.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.870 0.000 273.150 4.000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.470 0.000 277.750 4.000 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.610 0.000 281.890 4.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.850 0.000 164.130 4.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.210 0.000 286.490 4.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.350 0.000 290.630 4.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.950 0.000 295.230 4.000 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.090 0.000 299.370 4.000 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.690 0.000 303.970 4.000 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 307.830 0.000 308.110 4.000 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.430 0.000 312.710 4.000 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.570 0.000 316.850 4.000 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.170 0.000 321.450 4.000 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.310 0.000 325.590 4.000 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.990 0.000 168.270 4.000 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.910 0.000 330.190 4.000 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.050 0.000 334.330 4.000 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.650 0.000 338.930 4.000 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.790 0.000 343.070 4.000 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.390 0.000 347.670 4.000 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.530 0.000 351.810 4.000 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 356.130 0.000 356.410 4.000 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.270 0.000 360.550 4.000 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.870 0.000 365.150 4.000 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.010 0.000 369.290 4.000 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.590 0.000 172.870 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.610 0.000 373.890 4.000 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.210 0.000 378.490 4.000 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 382.350 0.000 382.630 4.000 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.950 0.000 387.230 4.000 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.090 0.000 391.370 4.000 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 395.690 0.000 395.970 4.000 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.830 0.000 400.110 4.000 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.430 0.000 404.710 4.000 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 408.570 0.000 408.850 4.000 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 413.170 0.000 413.450 4.000 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.730 0.000 177.010 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 417.310 0.000 417.590 4.000 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.910 0.000 422.190 4.000 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 426.050 0.000 426.330 4.000 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 430.650 0.000 430.930 4.000 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.790 0.000 435.070 4.000 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.390 0.000 439.670 4.000 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.530 0.000 443.810 4.000 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 448.130 0.000 448.410 4.000 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 452.270 0.000 452.550 4.000 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 456.870 0.000 457.150 4.000 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.330 0.000 181.610 4.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.010 0.000 461.290 4.000 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 465.610 0.000 465.890 4.000 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.750 0.000 470.030 4.000 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 474.350 0.000 474.630 4.000 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.490 0.000 478.770 4.000 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.090 0.000 483.370 4.000 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 487.230 0.000 487.510 4.000 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 491.830 0.000 492.110 4.000 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.970 0.000 496.250 4.000 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 500.570 0.000 500.850 4.000 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.470 0.000 185.750 4.000 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 504.710 0.000 504.990 4.000 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 509.310 0.000 509.590 4.000 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 513.450 0.000 513.730 4.000 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.050 0.000 518.330 4.000 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.190 0.000 522.470 4.000 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 526.790 0.000 527.070 4.000 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 530.930 0.000 531.210 4.000 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 535.530 0.000 535.810 4.000 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 539.670 0.000 539.950 4.000 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.270 0.000 544.550 4.000 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.070 0.000 190.350 4.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 548.410 0.000 548.690 4.000 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.010 0.000 553.290 4.000 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.150 0.000 557.430 4.000 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 561.750 0.000 562.030 4.000 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 565.890 0.000 566.170 4.000 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.490 0.000 570.770 4.000 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 574.630 0.000 574.910 4.000 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.230 0.000 579.510 4.000 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 583.370 0.000 583.650 4.000 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.970 0.000 588.250 4.000 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.210 0.000 194.490 4.000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.490 0.000 156.770 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.950 0.000 594.230 4.000 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 598.090 0.000 598.370 4.000 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 602.690 0.000 602.970 4.000 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 606.830 0.000 607.110 4.000 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.430 0.000 611.710 4.000 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 615.570 0.000 615.850 4.000 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 620.170 0.000 620.450 4.000 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 624.310 0.000 624.590 4.000 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 628.910 0.000 629.190 4.000 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 633.050 0.000 633.330 4.000 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.190 0.000 200.470 4.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 637.650 0.000 637.930 4.000 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 641.790 0.000 642.070 4.000 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 646.390 0.000 646.670 4.000 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.530 0.000 650.810 4.000 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 655.130 0.000 655.410 4.000 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 659.270 0.000 659.550 4.000 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 663.870 0.000 664.150 4.000 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 668.010 0.000 668.290 4.000 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 672.610 0.000 672.890 4.000 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.750 0.000 677.030 4.000 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.330 0.000 204.610 4.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 681.350 0.000 681.630 4.000 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.490 0.000 685.770 4.000 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 690.090 0.000 690.370 4.000 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 694.230 0.000 694.510 4.000 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 698.830 0.000 699.110 4.000 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.970 0.000 703.250 4.000 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 707.570 0.000 707.850 4.000 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 711.710 0.000 711.990 4.000 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.930 0.000 209.210 4.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.070 0.000 213.350 4.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.670 0.000 217.950 4.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.810 0.000 222.090 4.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.410 0.000 226.690 4.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.550 0.000 230.830 4.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.150 0.000 235.430 4.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.290 0.000 239.570 4.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.630 0.000 160.910 4.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.890 0.000 244.170 4.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.030 0.000 248.310 4.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.630 0.000 252.910 4.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.770 0.000 257.050 4.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.370 0.000 261.650 4.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.510 0.000 265.790 4.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.110 0.000 270.390 4.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.250 0.000 274.530 4.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.850 0.000 279.130 4.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.990 0.000 283.270 4.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.230 0.000 165.510 4.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.590 0.000 287.870 4.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.730 0.000 292.010 4.000 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.330 0.000 296.610 4.000 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.930 0.000 301.210 4.000 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.070 0.000 305.350 4.000 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.670 0.000 309.950 4.000 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 313.810 0.000 314.090 4.000 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.410 0.000 318.690 4.000 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.550 0.000 322.830 4.000 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.150 0.000 327.430 4.000 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.370 0.000 169.650 4.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.290 0.000 331.570 4.000 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.890 0.000 336.170 4.000 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.030 0.000 340.310 4.000 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.630 0.000 344.910 4.000 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 348.770 0.000 349.050 4.000 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 353.370 0.000 353.650 4.000 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.510 0.000 357.790 4.000 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.110 0.000 362.390 4.000 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.250 0.000 366.530 4.000 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.850 0.000 371.130 4.000 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 0.000 174.250 4.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.990 0.000 375.270 4.000 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.590 0.000 379.870 4.000 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.730 0.000 384.010 4.000 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 388.330 0.000 388.610 4.000 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.470 0.000 392.750 4.000 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.070 0.000 397.350 4.000 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 401.210 0.000 401.490 4.000 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.810 0.000 406.090 4.000 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.950 0.000 410.230 4.000 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 414.550 0.000 414.830 4.000 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.110 0.000 178.390 4.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.690 0.000 418.970 4.000 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 423.290 0.000 423.570 4.000 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 427.430 0.000 427.710 4.000 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.030 0.000 432.310 4.000 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 436.170 0.000 436.450 4.000 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 440.770 0.000 441.050 4.000 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 444.910 0.000 445.190 4.000 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.510 0.000 449.790 4.000 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 453.650 0.000 453.930 4.000 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 458.250 0.000 458.530 4.000 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.710 0.000 182.990 4.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 462.390 0.000 462.670 4.000 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.990 0.000 467.270 4.000 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 471.130 0.000 471.410 4.000 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 475.730 0.000 476.010 4.000 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.870 0.000 480.150 4.000 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.470 0.000 484.750 4.000 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 488.610 0.000 488.890 4.000 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 493.210 0.000 493.490 4.000 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 497.350 0.000 497.630 4.000 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.950 0.000 502.230 4.000 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.850 0.000 187.130 4.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 506.090 0.000 506.370 4.000 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 510.690 0.000 510.970 4.000 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 514.830 0.000 515.110 4.000 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 519.430 0.000 519.710 4.000 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 523.570 0.000 523.850 4.000 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.170 0.000 528.450 4.000 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 532.770 0.000 533.050 4.000 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 536.910 0.000 537.190 4.000 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.510 0.000 541.790 4.000 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 545.650 0.000 545.930 4.000 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.450 0.000 191.730 4.000 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 550.250 0.000 550.530 4.000 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 554.390 0.000 554.670 4.000 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 558.990 0.000 559.270 4.000 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 563.130 0.000 563.410 4.000 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 567.730 0.000 568.010 4.000 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 571.870 0.000 572.150 4.000 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.470 0.000 576.750 4.000 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 580.610 0.000 580.890 4.000 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 585.210 0.000 585.490 4.000 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 589.350 0.000 589.630 4.000 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.590 0.000 195.870 4.000 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 0.000 158.150 4.000 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 595.330 0.000 595.610 4.000 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.470 0.000 599.750 4.000 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 604.070 0.000 604.350 4.000 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.210 0.000 608.490 4.000 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 612.810 0.000 613.090 4.000 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 616.950 0.000 617.230 4.000 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 621.550 0.000 621.830 4.000 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 625.690 0.000 625.970 4.000 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 630.290 0.000 630.570 4.000 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.430 0.000 634.710 4.000 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.570 0.000 201.850 4.000 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 639.030 0.000 639.310 4.000 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 643.170 0.000 643.450 4.000 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 647.770 0.000 648.050 4.000 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 651.910 0.000 652.190 4.000 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.510 0.000 656.790 4.000 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 660.650 0.000 660.930 4.000 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 665.250 0.000 665.530 4.000 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 669.390 0.000 669.670 4.000 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.990 0.000 674.270 4.000 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 678.590 0.000 678.870 4.000 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.710 0.000 205.990 4.000 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 682.730 0.000 683.010 4.000 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 687.330 0.000 687.610 4.000 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 691.470 0.000 691.750 4.000 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 696.070 0.000 696.350 4.000 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 700.210 0.000 700.490 4.000 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 704.810 0.000 705.090 4.000 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.950 0.000 709.230 4.000 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 713.550 0.000 713.830 4.000 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.310 0.000 210.590 4.000 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.450 0.000 214.730 4.000 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 0.000 219.330 4.000 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.190 0.000 223.470 4.000 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.790 0.000 228.070 4.000 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.390 0.000 232.670 4.000 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.530 0.000 236.810 4.000 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.130 0.000 241.410 4.000 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.010 0.000 162.290 4.000 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.270 0.000 245.550 4.000 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.870 0.000 250.150 4.000 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.010 0.000 254.290 4.000 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.610 0.000 258.890 4.000 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.750 0.000 263.030 4.000 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.350 0.000 267.630 4.000 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.490 0.000 271.770 4.000 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.090 0.000 276.370 4.000 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.230 0.000 280.510 4.000 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.830 0.000 285.110 4.000 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.610 0.000 166.890 4.000 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.970 0.000 289.250 4.000 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.570 0.000 293.850 4.000 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.710 0.000 297.990 4.000 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.310 0.000 302.590 4.000 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.450 0.000 306.730 4.000 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.050 0.000 311.330 4.000 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.190 0.000 315.470 4.000 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.790 0.000 320.070 4.000 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.930 0.000 324.210 4.000 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.530 0.000 328.810 4.000 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 0.000 171.030 4.000 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.670 0.000 332.950 4.000 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.270 0.000 337.550 4.000 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.410 0.000 341.690 4.000 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.010 0.000 346.290 4.000 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 350.150 0.000 350.430 4.000 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.750 0.000 355.030 4.000 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.890 0.000 359.170 4.000 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.490 0.000 363.770 4.000 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.630 0.000 367.910 4.000 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 372.230 0.000 372.510 4.000 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.350 0.000 175.630 4.000 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.370 0.000 376.650 4.000 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.970 0.000 381.250 4.000 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 385.110 0.000 385.390 4.000 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.710 0.000 389.990 4.000 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 393.850 0.000 394.130 4.000 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.450 0.000 398.730 4.000 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.590 0.000 402.870 4.000 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 407.190 0.000 407.470 4.000 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 411.330 0.000 411.610 4.000 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.930 0.000 416.210 4.000 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.490 0.000 179.770 4.000 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.070 0.000 420.350 4.000 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 424.670 0.000 424.950 4.000 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.810 0.000 429.090 4.000 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 433.410 0.000 433.690 4.000 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 437.550 0.000 437.830 4.000 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 442.150 0.000 442.430 4.000 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 446.290 0.000 446.570 4.000 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.890 0.000 451.170 4.000 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.490 0.000 455.770 4.000 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 459.630 0.000 459.910 4.000 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.090 0.000 184.370 4.000 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 464.230 0.000 464.510 4.000 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 468.370 0.000 468.650 4.000 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.970 0.000 473.250 4.000 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 477.110 0.000 477.390 4.000 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 481.710 0.000 481.990 4.000 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 485.850 0.000 486.130 4.000 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 490.450 0.000 490.730 4.000 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 494.590 0.000 494.870 4.000 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.190 0.000 499.470 4.000 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 503.330 0.000 503.610 4.000 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.230 0.000 188.510 4.000 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.930 0.000 508.210 4.000 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.070 0.000 512.350 4.000 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 516.670 0.000 516.950 4.000 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 520.810 0.000 521.090 4.000 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 525.410 0.000 525.690 4.000 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 529.550 0.000 529.830 4.000 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.150 0.000 534.430 4.000 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 538.290 0.000 538.570 4.000 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 542.890 0.000 543.170 4.000 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.030 0.000 547.310 4.000 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.830 0.000 193.110 4.000 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 551.630 0.000 551.910 4.000 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 555.770 0.000 556.050 4.000 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.370 0.000 560.650 4.000 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.510 0.000 564.790 4.000 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 569.110 0.000 569.390 4.000 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.250 0.000 573.530 4.000 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 577.850 0.000 578.130 4.000 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.990 0.000 582.270 4.000 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.590 0.000 586.870 4.000 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 590.730 0.000 591.010 4.000 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.970 0.000 197.250 4.000 ;
    END
  END la_oenb[9]
  PIN o_addr1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.080 4.000 36.680 ;
    END
  END o_addr1[0]
  PIN o_addr1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.960 4.000 81.560 ;
    END
  END o_addr1[1]
  PIN o_addr1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.840 4.000 126.440 ;
    END
  END o_addr1[2]
  PIN o_addr1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.720 4.000 171.320 ;
    END
  END o_addr1[3]
  PIN o_addr1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 229.880 4.000 230.480 ;
    END
  END o_addr1[4]
  PIN o_addr1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 751.270 0.000 751.550 4.000 ;
    END
  END o_addr1[5]
  PIN o_addr1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 304.680 4.000 305.280 ;
    END
  END o_addr1[6]
  PIN o_addr1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 643.630 830.620 643.910 834.620 ;
    END
  END o_addr1[7]
  PIN o_addr1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 770.130 0.000 770.410 4.000 ;
    END
  END o_addr1[8]
  PIN o_addr1_1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.120 4.000 21.720 ;
    END
  END o_addr1_1[0]
  PIN o_addr1_1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 731.030 0.000 731.310 4.000 ;
    END
  END o_addr1_1[1]
  PIN o_addr1_1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.880 4.000 111.480 ;
    END
  END o_addr1_1[2]
  PIN o_addr1_1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 157.120 823.900 157.720 ;
    END
  END o_addr1_1[3]
  PIN o_addr1_1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 184.320 823.900 184.920 ;
    END
  END o_addr1_1[4]
  PIN o_addr1_1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.840 4.000 245.440 ;
    END
  END o_addr1_1[5]
  PIN o_addr1_1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 633.510 830.620 633.790 834.620 ;
    END
  END o_addr1_1[6]
  PIN o_addr1_1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 762.770 0.000 763.050 4.000 ;
    END
  END o_addr1_1[7]
  PIN o_addr1_1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 658.350 830.620 658.630 834.620 ;
    END
  END o_addr1_1[8]
  PIN o_csb0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 719.070 0.000 719.350 4.000 ;
    END
  END o_csb0
  PIN o_csb0_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 720.450 0.000 720.730 4.000 ;
    END
  END o_csb0_1
  PIN o_csb1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END o_csb1
  PIN o_csb1_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 6.840 823.900 7.440 ;
    END
  END o_csb1_1
  PIN o_din0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 725.050 0.000 725.330 4.000 ;
    END
  END o_din0[0]
  PIN o_din0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 348.200 823.900 348.800 ;
    END
  END o_din0[10]
  PIN o_din0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 687.790 830.620 688.070 834.620 ;
    END
  END o_din0[11]
  PIN o_din0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 692.850 830.620 693.130 834.620 ;
    END
  END o_din0[12]
  PIN o_din0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 782.090 0.000 782.370 4.000 ;
    END
  END o_din0[13]
  PIN o_din0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 783.470 0.000 783.750 4.000 ;
    END
  END o_din0[14]
  PIN o_din0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 722.290 830.620 722.570 834.620 ;
    END
  END o_din0[15]
  PIN o_din0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 788.990 0.000 789.270 4.000 ;
    END
  END o_din0[16]
  PIN o_din0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 737.010 830.620 737.290 834.620 ;
    END
  END o_din0[17]
  PIN o_din0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 527.720 4.000 528.320 ;
    END
  END o_din0[18]
  PIN o_din0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 797.730 0.000 798.010 4.000 ;
    END
  END o_din0[19]
  PIN o_din0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 733.790 0.000 734.070 4.000 ;
    END
  END o_din0[1]
  PIN o_din0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 761.850 830.620 762.130 834.620 ;
    END
  END o_din0[20]
  PIN o_din0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 567.160 823.900 567.760 ;
    END
  END o_din0[21]
  PIN o_din0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 594.360 823.900 594.960 ;
    END
  END o_din0[22]
  PIN o_din0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 809.690 0.000 809.970 4.000 ;
    END
  END o_din0[23]
  PIN o_din0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 781.630 830.620 781.910 834.620 ;
    END
  END o_din0[24]
  PIN o_din0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 649.440 823.900 650.040 ;
    END
  END o_din0[25]
  PIN o_din0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 706.560 4.000 707.160 ;
    END
  END o_din0[26]
  PIN o_din0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 801.410 830.620 801.690 834.620 ;
    END
  END o_din0[27]
  PIN o_din0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 811.070 830.620 811.350 834.620 ;
    END
  END o_din0[28]
  PIN o_din0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 758.920 823.900 759.520 ;
    END
  END o_din0[29]
  PIN o_din0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 102.040 823.900 102.640 ;
    END
  END o_din0[2]
  PIN o_din0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 786.120 823.900 786.720 ;
    END
  END o_din0[30]
  PIN o_din0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 826.920 823.900 827.520 ;
    END
  END o_din0[31]
  PIN o_din0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 185.000 4.000 185.600 ;
    END
  END o_din0[3]
  PIN o_din0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 746.670 0.000 746.950 4.000 ;
    END
  END o_din0[4]
  PIN o_din0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 274.760 4.000 275.360 ;
    END
  END o_din0[5]
  PIN o_din0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 238.720 823.900 239.320 ;
    END
  END o_din0[6]
  PIN o_din0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 648.230 830.620 648.510 834.620 ;
    END
  END o_din0[7]
  PIN o_din0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 348.880 4.000 349.480 ;
    END
  END o_din0[8]
  PIN o_din0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 668.010 830.620 668.290 834.620 ;
    END
  END o_din0[9]
  PIN o_din0_1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END o_din0_1[0]
  PIN o_din0_1[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 678.130 830.620 678.410 834.620 ;
    END
  END o_din0_1[10]
  PIN o_din0_1[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 776.110 0.000 776.390 4.000 ;
    END
  END o_din0_1[11]
  PIN o_din0_1[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 403.280 823.900 403.880 ;
    END
  END o_din0_1[12]
  PIN o_din0_1[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 468.560 4.000 469.160 ;
    END
  END o_din0_1[13]
  PIN o_din0_1[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.510 830.620 702.790 834.620 ;
    END
  END o_din0_1[14]
  PIN o_din0_1[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 483.520 4.000 484.120 ;
    END
  END o_din0_1[15]
  PIN o_din0_1[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 787.610 0.000 787.890 4.000 ;
    END
  END o_din0_1[16]
  PIN o_din0_1[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 792.210 0.000 792.490 4.000 ;
    END
  END o_din0_1[17]
  PIN o_din0_1[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 747.130 830.620 747.410 834.620 ;
    END
  END o_din0_1[18]
  PIN o_din0_1[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 557.640 4.000 558.240 ;
    END
  END o_din0_1[19]
  PIN o_din0_1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 732.410 0.000 732.690 4.000 ;
    END
  END o_din0_1[1]
  PIN o_din0_1[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 756.790 830.620 757.070 834.620 ;
    END
  END o_din0_1[20]
  PIN o_din0_1[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 553.560 823.900 554.160 ;
    END
  END o_din0_1[21]
  PIN o_din0_1[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 805.090 0.000 805.370 4.000 ;
    END
  END o_din0_1[22]
  PIN o_din0_1[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 808.310 0.000 808.590 4.000 ;
    END
  END o_din0_1[23]
  PIN o_din0_1[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 622.240 823.900 622.840 ;
    END
  END o_din0_1[24]
  PIN o_din0_1[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 813.830 0.000 814.110 4.000 ;
    END
  END o_din0_1[25]
  PIN o_din0_1[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 691.600 4.000 692.200 ;
    END
  END o_din0_1[26]
  PIN o_din0_1[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 676.640 823.900 677.240 ;
    END
  END o_din0_1[27]
  PIN o_din0_1[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 717.440 823.900 718.040 ;
    END
  END o_din0_1[28]
  PIN o_din0_1[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 821.190 830.620 821.470 834.620 ;
    END
  END o_din0_1[29]
  PIN o_din0_1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.950 830.620 594.230 834.620 ;
    END
  END o_din0_1[2]
  PIN o_din0_1[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 796.320 4.000 796.920 ;
    END
  END o_din0_1[30]
  PIN o_din0_1[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 826.240 4.000 826.840 ;
    END
  END o_din0_1[31]
  PIN o_din0_1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 742.530 0.000 742.810 4.000 ;
    END
  END o_din0_1[3]
  PIN o_din0_1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 745.290 0.000 745.570 4.000 ;
    END
  END o_din0_1[4]
  PIN o_din0_1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 259.800 4.000 260.400 ;
    END
  END o_din0_1[5]
  PIN o_din0_1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 758.630 0.000 758.910 4.000 ;
    END
  END o_din0_1[6]
  PIN o_din0_1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 280.200 823.900 280.800 ;
    END
  END o_din0_1[7]
  PIN o_din0_1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 771.510 0.000 771.790 4.000 ;
    END
  END o_din0_1[8]
  PIN o_din0_1[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 393.760 4.000 394.360 ;
    END
  END o_din0_1[9]
  PIN o_waddr0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 47.640 823.900 48.240 ;
    END
  END o_waddr0[0]
  PIN o_waddr0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 735.170 0.000 735.450 4.000 ;
    END
  END o_waddr0[1]
  PIN o_waddr0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 115.640 823.900 116.240 ;
    END
  END o_waddr0[2]
  PIN o_waddr0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 199.960 4.000 200.560 ;
    END
  END o_waddr0[3]
  PIN o_waddr0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 211.520 823.900 212.120 ;
    END
  END o_waddr0[4]
  PIN o_waddr0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 752.650 0.000 752.930 4.000 ;
    END
  END o_waddr0[5]
  PIN o_waddr0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 253.000 823.900 253.600 ;
    END
  END o_waddr0[6]
  PIN o_waddr0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 764.610 0.000 764.890 4.000 ;
    END
  END o_waddr0[7]
  PIN o_waddr0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 363.840 4.000 364.440 ;
    END
  END o_waddr0[8]
  PIN o_waddr0_1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 726.430 0.000 726.710 4.000 ;
    END
  END o_waddr0_1[0]
  PIN o_waddr0_1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.230 830.620 579.510 834.620 ;
    END
  END o_waddr0_1[1]
  PIN o_waddr0_1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 140.800 4.000 141.400 ;
    END
  END o_waddr0_1[2]
  PIN o_waddr0_1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 604.070 830.620 604.350 834.620 ;
    END
  END o_waddr0_1[3]
  PIN o_waddr0_1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 197.920 823.900 198.520 ;
    END
  END o_waddr0_1[4]
  PIN o_waddr0_1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 289.720 4.000 290.320 ;
    END
  END o_waddr0_1[5]
  PIN o_waddr0_1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 638.570 830.620 638.850 834.620 ;
    END
  END o_waddr0_1[6]
  PIN o_waddr0_1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 653.290 830.620 653.570 834.620 ;
    END
  END o_waddr0_1[7]
  PIN o_waddr0_1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 293.800 823.900 294.400 ;
    END
  END o_waddr0_1[8]
  PIN o_web0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.510 830.620 564.790 834.620 ;
    END
  END o_web0
  PIN o_web0_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 569.570 830.620 569.850 834.620 ;
    END
  END o_web0_1
  PIN o_wmask0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 574.630 830.620 574.910 834.620 ;
    END
  END o_wmask0[0]
  PIN o_wmask0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 584.290 830.620 584.570 834.620 ;
    END
  END o_wmask0[1]
  PIN o_wmask0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 155.760 4.000 156.360 ;
    END
  END o_wmask0[2]
  PIN o_wmask0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.900 170.720 823.900 171.320 ;
    END
  END o_wmask0[3]
  PIN o_wmask0_1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 727.810 0.000 728.090 4.000 ;
    END
  END o_wmask0_1[0]
  PIN o_wmask0_1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 736.550 0.000 736.830 4.000 ;
    END
  END o_wmask0_1[1]
  PIN o_wmask0_1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 739.770 0.000 740.050 4.000 ;
    END
  END o_wmask0_1[2]
  PIN o_wmask0_1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 609.130 830.620 609.410 834.620 ;
    END
  END o_wmask0_1[3]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 821.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 821.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 821.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 821.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 821.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 821.680 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 821.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 821.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 821.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 821.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 821.680 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.550 0.000 0.830 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.930 0.000 2.210 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 0.000 3.590 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.290 0.000 9.570 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.510 0.000 58.790 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.110 0.000 63.390 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.250 0.000 67.530 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.850 0.000 72.130 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.990 0.000 76.270 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.730 0.000 85.010 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.330 0.000 89.610 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 0.000 93.750 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.070 0.000 98.350 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.810 0.000 15.090 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.210 0.000 102.490 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.810 0.000 107.090 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.950 0.000 111.230 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.550 0.000 115.830 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.690 0.000 119.970 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.290 0.000 124.570 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.430 0.000 128.710 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.030 0.000 133.310 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.170 0.000 137.450 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.770 0.000 142.050 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 0.000 21.070 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.910 0.000 146.190 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.510 0.000 150.790 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.770 0.000 27.050 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.890 0.000 37.170 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.030 0.000 41.310 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.630 0.000 45.910 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.770 0.000 50.050 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.370 0.000 54.650 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.690 0.000 4.970 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.670 0.000 10.950 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.890 0.000 60.170 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.630 0.000 68.910 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.230 0.000 73.510 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.830 0.000 78.110 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.970 0.000 82.250 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.570 0.000 86.850 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.710 0.000 90.990 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.310 0.000 95.590 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.450 0.000 99.730 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.050 0.000 104.330 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.190 0.000 108.470 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 0.000 113.070 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.930 0.000 117.210 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.530 0.000 121.810 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 0.000 125.950 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.270 0.000 130.550 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.410 0.000 134.690 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.010 0.000 139.290 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.150 0.000 143.430 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.170 0.000 22.450 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.750 0.000 148.030 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.890 0.000 152.170 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.150 0.000 28.430 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.670 0.000 33.950 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.270 0.000 38.550 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.410 0.000 42.690 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.010 0.000 47.290 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.150 0.000 51.430 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.750 0.000 56.030 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.050 0.000 12.330 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.730 0.000 62.010 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.870 0.000 66.150 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.470 0.000 70.750 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.610 0.000 74.890 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.210 0.000 79.490 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.350 0.000 83.630 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.950 0.000 88.230 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.090 0.000 92.370 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.830 0.000 101.110 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.030 0.000 18.310 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.430 0.000 105.710 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.170 0.000 114.450 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.310 0.000 118.590 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.910 0.000 123.190 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.050 0.000 127.330 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.650 0.000 131.930 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.790 0.000 136.070 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.390 0.000 140.670 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.530 0.000 144.810 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.550 0.000 23.830 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.130 0.000 149.410 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.270 0.000 153.550 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.530 0.000 29.810 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.650 0.000 39.930 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.250 0.000 44.530 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.990 0.000 53.270 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.130 0.000 57.410 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.430 0.000 13.710 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 4.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.930 0.000 25.210 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.910 0.000 31.190 4.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.070 0.000 6.350 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.450 0.000 7.730 4.000 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 5.865 823.715 827.135 ;
      LAYER met1 ;
        RECT 0.070 2.420 823.790 827.180 ;
      LAYER met2 ;
        RECT 0.100 830.340 2.110 830.620 ;
        RECT 2.950 830.340 6.710 830.620 ;
        RECT 7.550 830.340 11.770 830.620 ;
        RECT 12.610 830.340 16.830 830.620 ;
        RECT 17.670 830.340 21.430 830.620 ;
        RECT 22.270 830.340 26.490 830.620 ;
        RECT 27.330 830.340 31.550 830.620 ;
        RECT 32.390 830.340 36.610 830.620 ;
        RECT 37.450 830.340 41.210 830.620 ;
        RECT 42.050 830.340 46.270 830.620 ;
        RECT 47.110 830.340 51.330 830.620 ;
        RECT 52.170 830.340 55.930 830.620 ;
        RECT 56.770 830.340 60.990 830.620 ;
        RECT 61.830 830.340 66.050 830.620 ;
        RECT 66.890 830.340 71.110 830.620 ;
        RECT 71.950 830.340 75.710 830.620 ;
        RECT 76.550 830.340 80.770 830.620 ;
        RECT 81.610 830.340 85.830 830.620 ;
        RECT 86.670 830.340 90.890 830.620 ;
        RECT 91.730 830.340 95.490 830.620 ;
        RECT 96.330 830.340 100.550 830.620 ;
        RECT 101.390 830.340 105.610 830.620 ;
        RECT 106.450 830.340 110.210 830.620 ;
        RECT 111.050 830.340 115.270 830.620 ;
        RECT 116.110 830.340 120.330 830.620 ;
        RECT 121.170 830.340 125.390 830.620 ;
        RECT 126.230 830.340 129.990 830.620 ;
        RECT 130.830 830.340 135.050 830.620 ;
        RECT 135.890 830.340 140.110 830.620 ;
        RECT 140.950 830.340 145.170 830.620 ;
        RECT 146.010 830.340 149.770 830.620 ;
        RECT 150.610 830.340 154.830 830.620 ;
        RECT 155.670 830.340 159.890 830.620 ;
        RECT 160.730 830.340 164.490 830.620 ;
        RECT 165.330 830.340 169.550 830.620 ;
        RECT 170.390 830.340 174.610 830.620 ;
        RECT 175.450 830.340 179.670 830.620 ;
        RECT 180.510 830.340 184.270 830.620 ;
        RECT 185.110 830.340 189.330 830.620 ;
        RECT 190.170 830.340 194.390 830.620 ;
        RECT 195.230 830.340 198.990 830.620 ;
        RECT 199.830 830.340 204.050 830.620 ;
        RECT 204.890 830.340 209.110 830.620 ;
        RECT 209.950 830.340 214.170 830.620 ;
        RECT 215.010 830.340 218.770 830.620 ;
        RECT 219.610 830.340 223.830 830.620 ;
        RECT 224.670 830.340 228.890 830.620 ;
        RECT 229.730 830.340 233.950 830.620 ;
        RECT 234.790 830.340 238.550 830.620 ;
        RECT 239.390 830.340 243.610 830.620 ;
        RECT 244.450 830.340 248.670 830.620 ;
        RECT 249.510 830.340 253.270 830.620 ;
        RECT 254.110 830.340 258.330 830.620 ;
        RECT 259.170 830.340 263.390 830.620 ;
        RECT 264.230 830.340 268.450 830.620 ;
        RECT 269.290 830.340 273.050 830.620 ;
        RECT 273.890 830.340 278.110 830.620 ;
        RECT 278.950 830.340 283.170 830.620 ;
        RECT 284.010 830.340 288.230 830.620 ;
        RECT 289.070 830.340 292.830 830.620 ;
        RECT 293.670 830.340 297.890 830.620 ;
        RECT 298.730 830.340 302.950 830.620 ;
        RECT 303.790 830.340 307.550 830.620 ;
        RECT 308.390 830.340 312.610 830.620 ;
        RECT 313.450 830.340 317.670 830.620 ;
        RECT 318.510 830.340 322.730 830.620 ;
        RECT 323.570 830.340 327.330 830.620 ;
        RECT 328.170 830.340 332.390 830.620 ;
        RECT 333.230 830.340 337.450 830.620 ;
        RECT 338.290 830.340 342.050 830.620 ;
        RECT 342.890 830.340 347.110 830.620 ;
        RECT 347.950 830.340 352.170 830.620 ;
        RECT 353.010 830.340 357.230 830.620 ;
        RECT 358.070 830.340 361.830 830.620 ;
        RECT 362.670 830.340 366.890 830.620 ;
        RECT 367.730 830.340 371.950 830.620 ;
        RECT 372.790 830.340 377.010 830.620 ;
        RECT 377.850 830.340 381.610 830.620 ;
        RECT 382.450 830.340 386.670 830.620 ;
        RECT 387.510 830.340 391.730 830.620 ;
        RECT 392.570 830.340 396.330 830.620 ;
        RECT 397.170 830.340 401.390 830.620 ;
        RECT 402.230 830.340 406.450 830.620 ;
        RECT 407.290 830.340 411.510 830.620 ;
        RECT 412.350 830.340 416.110 830.620 ;
        RECT 416.950 830.340 421.170 830.620 ;
        RECT 422.010 830.340 426.230 830.620 ;
        RECT 427.070 830.340 431.290 830.620 ;
        RECT 432.130 830.340 435.890 830.620 ;
        RECT 436.730 830.340 440.950 830.620 ;
        RECT 441.790 830.340 446.010 830.620 ;
        RECT 446.850 830.340 450.610 830.620 ;
        RECT 451.450 830.340 455.670 830.620 ;
        RECT 456.510 830.340 460.730 830.620 ;
        RECT 461.570 830.340 465.790 830.620 ;
        RECT 466.630 830.340 470.390 830.620 ;
        RECT 471.230 830.340 475.450 830.620 ;
        RECT 476.290 830.340 480.510 830.620 ;
        RECT 481.350 830.340 485.570 830.620 ;
        RECT 486.410 830.340 490.170 830.620 ;
        RECT 491.010 830.340 495.230 830.620 ;
        RECT 496.070 830.340 500.290 830.620 ;
        RECT 501.130 830.340 504.890 830.620 ;
        RECT 505.730 830.340 509.950 830.620 ;
        RECT 510.790 830.340 515.010 830.620 ;
        RECT 515.850 830.340 520.070 830.620 ;
        RECT 520.910 830.340 524.670 830.620 ;
        RECT 525.510 830.340 529.730 830.620 ;
        RECT 530.570 830.340 534.790 830.620 ;
        RECT 535.630 830.340 539.390 830.620 ;
        RECT 540.230 830.340 544.450 830.620 ;
        RECT 545.290 830.340 549.510 830.620 ;
        RECT 550.350 830.340 554.570 830.620 ;
        RECT 555.410 830.340 559.170 830.620 ;
        RECT 560.010 830.340 564.230 830.620 ;
        RECT 565.070 830.340 569.290 830.620 ;
        RECT 570.130 830.340 574.350 830.620 ;
        RECT 575.190 830.340 578.950 830.620 ;
        RECT 579.790 830.340 584.010 830.620 ;
        RECT 584.850 830.340 589.070 830.620 ;
        RECT 589.910 830.340 593.670 830.620 ;
        RECT 594.510 830.340 598.730 830.620 ;
        RECT 599.570 830.340 603.790 830.620 ;
        RECT 604.630 830.340 608.850 830.620 ;
        RECT 609.690 830.340 613.450 830.620 ;
        RECT 614.290 830.340 618.510 830.620 ;
        RECT 619.350 830.340 623.570 830.620 ;
        RECT 624.410 830.340 628.630 830.620 ;
        RECT 629.470 830.340 633.230 830.620 ;
        RECT 634.070 830.340 638.290 830.620 ;
        RECT 639.130 830.340 643.350 830.620 ;
        RECT 644.190 830.340 647.950 830.620 ;
        RECT 648.790 830.340 653.010 830.620 ;
        RECT 653.850 830.340 658.070 830.620 ;
        RECT 658.910 830.340 663.130 830.620 ;
        RECT 663.970 830.340 667.730 830.620 ;
        RECT 668.570 830.340 672.790 830.620 ;
        RECT 673.630 830.340 677.850 830.620 ;
        RECT 678.690 830.340 682.450 830.620 ;
        RECT 683.290 830.340 687.510 830.620 ;
        RECT 688.350 830.340 692.570 830.620 ;
        RECT 693.410 830.340 697.630 830.620 ;
        RECT 698.470 830.340 702.230 830.620 ;
        RECT 703.070 830.340 707.290 830.620 ;
        RECT 708.130 830.340 712.350 830.620 ;
        RECT 713.190 830.340 717.410 830.620 ;
        RECT 718.250 830.340 722.010 830.620 ;
        RECT 722.850 830.340 727.070 830.620 ;
        RECT 727.910 830.340 732.130 830.620 ;
        RECT 732.970 830.340 736.730 830.620 ;
        RECT 737.570 830.340 741.790 830.620 ;
        RECT 742.630 830.340 746.850 830.620 ;
        RECT 747.690 830.340 751.910 830.620 ;
        RECT 752.750 830.340 756.510 830.620 ;
        RECT 757.350 830.340 761.570 830.620 ;
        RECT 762.410 830.340 766.630 830.620 ;
        RECT 767.470 830.340 771.690 830.620 ;
        RECT 772.530 830.340 776.290 830.620 ;
        RECT 777.130 830.340 781.350 830.620 ;
        RECT 782.190 830.340 786.410 830.620 ;
        RECT 787.250 830.340 791.010 830.620 ;
        RECT 791.850 830.340 796.070 830.620 ;
        RECT 796.910 830.340 801.130 830.620 ;
        RECT 801.970 830.340 806.190 830.620 ;
        RECT 807.030 830.340 810.790 830.620 ;
        RECT 811.630 830.340 815.850 830.620 ;
        RECT 816.690 830.340 820.910 830.620 ;
        RECT 821.750 830.340 823.770 830.620 ;
        RECT 0.100 4.280 823.770 830.340 ;
        RECT 0.100 2.390 0.270 4.280 ;
        RECT 1.110 2.390 1.650 4.280 ;
        RECT 2.490 2.390 3.030 4.280 ;
        RECT 3.870 2.390 4.410 4.280 ;
        RECT 5.250 2.390 5.790 4.280 ;
        RECT 6.630 2.390 7.170 4.280 ;
        RECT 8.010 2.390 9.010 4.280 ;
        RECT 9.850 2.390 10.390 4.280 ;
        RECT 11.230 2.390 11.770 4.280 ;
        RECT 12.610 2.390 13.150 4.280 ;
        RECT 13.990 2.390 14.530 4.280 ;
        RECT 15.370 2.390 15.910 4.280 ;
        RECT 16.750 2.390 17.750 4.280 ;
        RECT 18.590 2.390 19.130 4.280 ;
        RECT 19.970 2.390 20.510 4.280 ;
        RECT 21.350 2.390 21.890 4.280 ;
        RECT 22.730 2.390 23.270 4.280 ;
        RECT 24.110 2.390 24.650 4.280 ;
        RECT 25.490 2.390 26.490 4.280 ;
        RECT 27.330 2.390 27.870 4.280 ;
        RECT 28.710 2.390 29.250 4.280 ;
        RECT 30.090 2.390 30.630 4.280 ;
        RECT 31.470 2.390 32.010 4.280 ;
        RECT 32.850 2.390 33.390 4.280 ;
        RECT 34.230 2.390 35.230 4.280 ;
        RECT 36.070 2.390 36.610 4.280 ;
        RECT 37.450 2.390 37.990 4.280 ;
        RECT 38.830 2.390 39.370 4.280 ;
        RECT 40.210 2.390 40.750 4.280 ;
        RECT 41.590 2.390 42.130 4.280 ;
        RECT 42.970 2.390 43.970 4.280 ;
        RECT 44.810 2.390 45.350 4.280 ;
        RECT 46.190 2.390 46.730 4.280 ;
        RECT 47.570 2.390 48.110 4.280 ;
        RECT 48.950 2.390 49.490 4.280 ;
        RECT 50.330 2.390 50.870 4.280 ;
        RECT 51.710 2.390 52.710 4.280 ;
        RECT 53.550 2.390 54.090 4.280 ;
        RECT 54.930 2.390 55.470 4.280 ;
        RECT 56.310 2.390 56.850 4.280 ;
        RECT 57.690 2.390 58.230 4.280 ;
        RECT 59.070 2.390 59.610 4.280 ;
        RECT 60.450 2.390 61.450 4.280 ;
        RECT 62.290 2.390 62.830 4.280 ;
        RECT 63.670 2.390 64.210 4.280 ;
        RECT 65.050 2.390 65.590 4.280 ;
        RECT 66.430 2.390 66.970 4.280 ;
        RECT 67.810 2.390 68.350 4.280 ;
        RECT 69.190 2.390 70.190 4.280 ;
        RECT 71.030 2.390 71.570 4.280 ;
        RECT 72.410 2.390 72.950 4.280 ;
        RECT 73.790 2.390 74.330 4.280 ;
        RECT 75.170 2.390 75.710 4.280 ;
        RECT 76.550 2.390 77.550 4.280 ;
        RECT 78.390 2.390 78.930 4.280 ;
        RECT 79.770 2.390 80.310 4.280 ;
        RECT 81.150 2.390 81.690 4.280 ;
        RECT 82.530 2.390 83.070 4.280 ;
        RECT 83.910 2.390 84.450 4.280 ;
        RECT 85.290 2.390 86.290 4.280 ;
        RECT 87.130 2.390 87.670 4.280 ;
        RECT 88.510 2.390 89.050 4.280 ;
        RECT 89.890 2.390 90.430 4.280 ;
        RECT 91.270 2.390 91.810 4.280 ;
        RECT 92.650 2.390 93.190 4.280 ;
        RECT 94.030 2.390 95.030 4.280 ;
        RECT 95.870 2.390 96.410 4.280 ;
        RECT 97.250 2.390 97.790 4.280 ;
        RECT 98.630 2.390 99.170 4.280 ;
        RECT 100.010 2.390 100.550 4.280 ;
        RECT 101.390 2.390 101.930 4.280 ;
        RECT 102.770 2.390 103.770 4.280 ;
        RECT 104.610 2.390 105.150 4.280 ;
        RECT 105.990 2.390 106.530 4.280 ;
        RECT 107.370 2.390 107.910 4.280 ;
        RECT 108.750 2.390 109.290 4.280 ;
        RECT 110.130 2.390 110.670 4.280 ;
        RECT 111.510 2.390 112.510 4.280 ;
        RECT 113.350 2.390 113.890 4.280 ;
        RECT 114.730 2.390 115.270 4.280 ;
        RECT 116.110 2.390 116.650 4.280 ;
        RECT 117.490 2.390 118.030 4.280 ;
        RECT 118.870 2.390 119.410 4.280 ;
        RECT 120.250 2.390 121.250 4.280 ;
        RECT 122.090 2.390 122.630 4.280 ;
        RECT 123.470 2.390 124.010 4.280 ;
        RECT 124.850 2.390 125.390 4.280 ;
        RECT 126.230 2.390 126.770 4.280 ;
        RECT 127.610 2.390 128.150 4.280 ;
        RECT 128.990 2.390 129.990 4.280 ;
        RECT 130.830 2.390 131.370 4.280 ;
        RECT 132.210 2.390 132.750 4.280 ;
        RECT 133.590 2.390 134.130 4.280 ;
        RECT 134.970 2.390 135.510 4.280 ;
        RECT 136.350 2.390 136.890 4.280 ;
        RECT 137.730 2.390 138.730 4.280 ;
        RECT 139.570 2.390 140.110 4.280 ;
        RECT 140.950 2.390 141.490 4.280 ;
        RECT 142.330 2.390 142.870 4.280 ;
        RECT 143.710 2.390 144.250 4.280 ;
        RECT 145.090 2.390 145.630 4.280 ;
        RECT 146.470 2.390 147.470 4.280 ;
        RECT 148.310 2.390 148.850 4.280 ;
        RECT 149.690 2.390 150.230 4.280 ;
        RECT 151.070 2.390 151.610 4.280 ;
        RECT 152.450 2.390 152.990 4.280 ;
        RECT 153.830 2.390 154.830 4.280 ;
        RECT 155.670 2.390 156.210 4.280 ;
        RECT 157.050 2.390 157.590 4.280 ;
        RECT 158.430 2.390 158.970 4.280 ;
        RECT 159.810 2.390 160.350 4.280 ;
        RECT 161.190 2.390 161.730 4.280 ;
        RECT 162.570 2.390 163.570 4.280 ;
        RECT 164.410 2.390 164.950 4.280 ;
        RECT 165.790 2.390 166.330 4.280 ;
        RECT 167.170 2.390 167.710 4.280 ;
        RECT 168.550 2.390 169.090 4.280 ;
        RECT 169.930 2.390 170.470 4.280 ;
        RECT 171.310 2.390 172.310 4.280 ;
        RECT 173.150 2.390 173.690 4.280 ;
        RECT 174.530 2.390 175.070 4.280 ;
        RECT 175.910 2.390 176.450 4.280 ;
        RECT 177.290 2.390 177.830 4.280 ;
        RECT 178.670 2.390 179.210 4.280 ;
        RECT 180.050 2.390 181.050 4.280 ;
        RECT 181.890 2.390 182.430 4.280 ;
        RECT 183.270 2.390 183.810 4.280 ;
        RECT 184.650 2.390 185.190 4.280 ;
        RECT 186.030 2.390 186.570 4.280 ;
        RECT 187.410 2.390 187.950 4.280 ;
        RECT 188.790 2.390 189.790 4.280 ;
        RECT 190.630 2.390 191.170 4.280 ;
        RECT 192.010 2.390 192.550 4.280 ;
        RECT 193.390 2.390 193.930 4.280 ;
        RECT 194.770 2.390 195.310 4.280 ;
        RECT 196.150 2.390 196.690 4.280 ;
        RECT 197.530 2.390 198.530 4.280 ;
        RECT 199.370 2.390 199.910 4.280 ;
        RECT 200.750 2.390 201.290 4.280 ;
        RECT 202.130 2.390 202.670 4.280 ;
        RECT 203.510 2.390 204.050 4.280 ;
        RECT 204.890 2.390 205.430 4.280 ;
        RECT 206.270 2.390 207.270 4.280 ;
        RECT 208.110 2.390 208.650 4.280 ;
        RECT 209.490 2.390 210.030 4.280 ;
        RECT 210.870 2.390 211.410 4.280 ;
        RECT 212.250 2.390 212.790 4.280 ;
        RECT 213.630 2.390 214.170 4.280 ;
        RECT 215.010 2.390 216.010 4.280 ;
        RECT 216.850 2.390 217.390 4.280 ;
        RECT 218.230 2.390 218.770 4.280 ;
        RECT 219.610 2.390 220.150 4.280 ;
        RECT 220.990 2.390 221.530 4.280 ;
        RECT 222.370 2.390 222.910 4.280 ;
        RECT 223.750 2.390 224.750 4.280 ;
        RECT 225.590 2.390 226.130 4.280 ;
        RECT 226.970 2.390 227.510 4.280 ;
        RECT 228.350 2.390 228.890 4.280 ;
        RECT 229.730 2.390 230.270 4.280 ;
        RECT 231.110 2.390 232.110 4.280 ;
        RECT 232.950 2.390 233.490 4.280 ;
        RECT 234.330 2.390 234.870 4.280 ;
        RECT 235.710 2.390 236.250 4.280 ;
        RECT 237.090 2.390 237.630 4.280 ;
        RECT 238.470 2.390 239.010 4.280 ;
        RECT 239.850 2.390 240.850 4.280 ;
        RECT 241.690 2.390 242.230 4.280 ;
        RECT 243.070 2.390 243.610 4.280 ;
        RECT 244.450 2.390 244.990 4.280 ;
        RECT 245.830 2.390 246.370 4.280 ;
        RECT 247.210 2.390 247.750 4.280 ;
        RECT 248.590 2.390 249.590 4.280 ;
        RECT 250.430 2.390 250.970 4.280 ;
        RECT 251.810 2.390 252.350 4.280 ;
        RECT 253.190 2.390 253.730 4.280 ;
        RECT 254.570 2.390 255.110 4.280 ;
        RECT 255.950 2.390 256.490 4.280 ;
        RECT 257.330 2.390 258.330 4.280 ;
        RECT 259.170 2.390 259.710 4.280 ;
        RECT 260.550 2.390 261.090 4.280 ;
        RECT 261.930 2.390 262.470 4.280 ;
        RECT 263.310 2.390 263.850 4.280 ;
        RECT 264.690 2.390 265.230 4.280 ;
        RECT 266.070 2.390 267.070 4.280 ;
        RECT 267.910 2.390 268.450 4.280 ;
        RECT 269.290 2.390 269.830 4.280 ;
        RECT 270.670 2.390 271.210 4.280 ;
        RECT 272.050 2.390 272.590 4.280 ;
        RECT 273.430 2.390 273.970 4.280 ;
        RECT 274.810 2.390 275.810 4.280 ;
        RECT 276.650 2.390 277.190 4.280 ;
        RECT 278.030 2.390 278.570 4.280 ;
        RECT 279.410 2.390 279.950 4.280 ;
        RECT 280.790 2.390 281.330 4.280 ;
        RECT 282.170 2.390 282.710 4.280 ;
        RECT 283.550 2.390 284.550 4.280 ;
        RECT 285.390 2.390 285.930 4.280 ;
        RECT 286.770 2.390 287.310 4.280 ;
        RECT 288.150 2.390 288.690 4.280 ;
        RECT 289.530 2.390 290.070 4.280 ;
        RECT 290.910 2.390 291.450 4.280 ;
        RECT 292.290 2.390 293.290 4.280 ;
        RECT 294.130 2.390 294.670 4.280 ;
        RECT 295.510 2.390 296.050 4.280 ;
        RECT 296.890 2.390 297.430 4.280 ;
        RECT 298.270 2.390 298.810 4.280 ;
        RECT 299.650 2.390 300.650 4.280 ;
        RECT 301.490 2.390 302.030 4.280 ;
        RECT 302.870 2.390 303.410 4.280 ;
        RECT 304.250 2.390 304.790 4.280 ;
        RECT 305.630 2.390 306.170 4.280 ;
        RECT 307.010 2.390 307.550 4.280 ;
        RECT 308.390 2.390 309.390 4.280 ;
        RECT 310.230 2.390 310.770 4.280 ;
        RECT 311.610 2.390 312.150 4.280 ;
        RECT 312.990 2.390 313.530 4.280 ;
        RECT 314.370 2.390 314.910 4.280 ;
        RECT 315.750 2.390 316.290 4.280 ;
        RECT 317.130 2.390 318.130 4.280 ;
        RECT 318.970 2.390 319.510 4.280 ;
        RECT 320.350 2.390 320.890 4.280 ;
        RECT 321.730 2.390 322.270 4.280 ;
        RECT 323.110 2.390 323.650 4.280 ;
        RECT 324.490 2.390 325.030 4.280 ;
        RECT 325.870 2.390 326.870 4.280 ;
        RECT 327.710 2.390 328.250 4.280 ;
        RECT 329.090 2.390 329.630 4.280 ;
        RECT 330.470 2.390 331.010 4.280 ;
        RECT 331.850 2.390 332.390 4.280 ;
        RECT 333.230 2.390 333.770 4.280 ;
        RECT 334.610 2.390 335.610 4.280 ;
        RECT 336.450 2.390 336.990 4.280 ;
        RECT 337.830 2.390 338.370 4.280 ;
        RECT 339.210 2.390 339.750 4.280 ;
        RECT 340.590 2.390 341.130 4.280 ;
        RECT 341.970 2.390 342.510 4.280 ;
        RECT 343.350 2.390 344.350 4.280 ;
        RECT 345.190 2.390 345.730 4.280 ;
        RECT 346.570 2.390 347.110 4.280 ;
        RECT 347.950 2.390 348.490 4.280 ;
        RECT 349.330 2.390 349.870 4.280 ;
        RECT 350.710 2.390 351.250 4.280 ;
        RECT 352.090 2.390 353.090 4.280 ;
        RECT 353.930 2.390 354.470 4.280 ;
        RECT 355.310 2.390 355.850 4.280 ;
        RECT 356.690 2.390 357.230 4.280 ;
        RECT 358.070 2.390 358.610 4.280 ;
        RECT 359.450 2.390 359.990 4.280 ;
        RECT 360.830 2.390 361.830 4.280 ;
        RECT 362.670 2.390 363.210 4.280 ;
        RECT 364.050 2.390 364.590 4.280 ;
        RECT 365.430 2.390 365.970 4.280 ;
        RECT 366.810 2.390 367.350 4.280 ;
        RECT 368.190 2.390 368.730 4.280 ;
        RECT 369.570 2.390 370.570 4.280 ;
        RECT 371.410 2.390 371.950 4.280 ;
        RECT 372.790 2.390 373.330 4.280 ;
        RECT 374.170 2.390 374.710 4.280 ;
        RECT 375.550 2.390 376.090 4.280 ;
        RECT 376.930 2.390 377.930 4.280 ;
        RECT 378.770 2.390 379.310 4.280 ;
        RECT 380.150 2.390 380.690 4.280 ;
        RECT 381.530 2.390 382.070 4.280 ;
        RECT 382.910 2.390 383.450 4.280 ;
        RECT 384.290 2.390 384.830 4.280 ;
        RECT 385.670 2.390 386.670 4.280 ;
        RECT 387.510 2.390 388.050 4.280 ;
        RECT 388.890 2.390 389.430 4.280 ;
        RECT 390.270 2.390 390.810 4.280 ;
        RECT 391.650 2.390 392.190 4.280 ;
        RECT 393.030 2.390 393.570 4.280 ;
        RECT 394.410 2.390 395.410 4.280 ;
        RECT 396.250 2.390 396.790 4.280 ;
        RECT 397.630 2.390 398.170 4.280 ;
        RECT 399.010 2.390 399.550 4.280 ;
        RECT 400.390 2.390 400.930 4.280 ;
        RECT 401.770 2.390 402.310 4.280 ;
        RECT 403.150 2.390 404.150 4.280 ;
        RECT 404.990 2.390 405.530 4.280 ;
        RECT 406.370 2.390 406.910 4.280 ;
        RECT 407.750 2.390 408.290 4.280 ;
        RECT 409.130 2.390 409.670 4.280 ;
        RECT 410.510 2.390 411.050 4.280 ;
        RECT 411.890 2.390 412.890 4.280 ;
        RECT 413.730 2.390 414.270 4.280 ;
        RECT 415.110 2.390 415.650 4.280 ;
        RECT 416.490 2.390 417.030 4.280 ;
        RECT 417.870 2.390 418.410 4.280 ;
        RECT 419.250 2.390 419.790 4.280 ;
        RECT 420.630 2.390 421.630 4.280 ;
        RECT 422.470 2.390 423.010 4.280 ;
        RECT 423.850 2.390 424.390 4.280 ;
        RECT 425.230 2.390 425.770 4.280 ;
        RECT 426.610 2.390 427.150 4.280 ;
        RECT 427.990 2.390 428.530 4.280 ;
        RECT 429.370 2.390 430.370 4.280 ;
        RECT 431.210 2.390 431.750 4.280 ;
        RECT 432.590 2.390 433.130 4.280 ;
        RECT 433.970 2.390 434.510 4.280 ;
        RECT 435.350 2.390 435.890 4.280 ;
        RECT 436.730 2.390 437.270 4.280 ;
        RECT 438.110 2.390 439.110 4.280 ;
        RECT 439.950 2.390 440.490 4.280 ;
        RECT 441.330 2.390 441.870 4.280 ;
        RECT 442.710 2.390 443.250 4.280 ;
        RECT 444.090 2.390 444.630 4.280 ;
        RECT 445.470 2.390 446.010 4.280 ;
        RECT 446.850 2.390 447.850 4.280 ;
        RECT 448.690 2.390 449.230 4.280 ;
        RECT 450.070 2.390 450.610 4.280 ;
        RECT 451.450 2.390 451.990 4.280 ;
        RECT 452.830 2.390 453.370 4.280 ;
        RECT 454.210 2.390 455.210 4.280 ;
        RECT 456.050 2.390 456.590 4.280 ;
        RECT 457.430 2.390 457.970 4.280 ;
        RECT 458.810 2.390 459.350 4.280 ;
        RECT 460.190 2.390 460.730 4.280 ;
        RECT 461.570 2.390 462.110 4.280 ;
        RECT 462.950 2.390 463.950 4.280 ;
        RECT 464.790 2.390 465.330 4.280 ;
        RECT 466.170 2.390 466.710 4.280 ;
        RECT 467.550 2.390 468.090 4.280 ;
        RECT 468.930 2.390 469.470 4.280 ;
        RECT 470.310 2.390 470.850 4.280 ;
        RECT 471.690 2.390 472.690 4.280 ;
        RECT 473.530 2.390 474.070 4.280 ;
        RECT 474.910 2.390 475.450 4.280 ;
        RECT 476.290 2.390 476.830 4.280 ;
        RECT 477.670 2.390 478.210 4.280 ;
        RECT 479.050 2.390 479.590 4.280 ;
        RECT 480.430 2.390 481.430 4.280 ;
        RECT 482.270 2.390 482.810 4.280 ;
        RECT 483.650 2.390 484.190 4.280 ;
        RECT 485.030 2.390 485.570 4.280 ;
        RECT 486.410 2.390 486.950 4.280 ;
        RECT 487.790 2.390 488.330 4.280 ;
        RECT 489.170 2.390 490.170 4.280 ;
        RECT 491.010 2.390 491.550 4.280 ;
        RECT 492.390 2.390 492.930 4.280 ;
        RECT 493.770 2.390 494.310 4.280 ;
        RECT 495.150 2.390 495.690 4.280 ;
        RECT 496.530 2.390 497.070 4.280 ;
        RECT 497.910 2.390 498.910 4.280 ;
        RECT 499.750 2.390 500.290 4.280 ;
        RECT 501.130 2.390 501.670 4.280 ;
        RECT 502.510 2.390 503.050 4.280 ;
        RECT 503.890 2.390 504.430 4.280 ;
        RECT 505.270 2.390 505.810 4.280 ;
        RECT 506.650 2.390 507.650 4.280 ;
        RECT 508.490 2.390 509.030 4.280 ;
        RECT 509.870 2.390 510.410 4.280 ;
        RECT 511.250 2.390 511.790 4.280 ;
        RECT 512.630 2.390 513.170 4.280 ;
        RECT 514.010 2.390 514.550 4.280 ;
        RECT 515.390 2.390 516.390 4.280 ;
        RECT 517.230 2.390 517.770 4.280 ;
        RECT 518.610 2.390 519.150 4.280 ;
        RECT 519.990 2.390 520.530 4.280 ;
        RECT 521.370 2.390 521.910 4.280 ;
        RECT 522.750 2.390 523.290 4.280 ;
        RECT 524.130 2.390 525.130 4.280 ;
        RECT 525.970 2.390 526.510 4.280 ;
        RECT 527.350 2.390 527.890 4.280 ;
        RECT 528.730 2.390 529.270 4.280 ;
        RECT 530.110 2.390 530.650 4.280 ;
        RECT 531.490 2.390 532.490 4.280 ;
        RECT 533.330 2.390 533.870 4.280 ;
        RECT 534.710 2.390 535.250 4.280 ;
        RECT 536.090 2.390 536.630 4.280 ;
        RECT 537.470 2.390 538.010 4.280 ;
        RECT 538.850 2.390 539.390 4.280 ;
        RECT 540.230 2.390 541.230 4.280 ;
        RECT 542.070 2.390 542.610 4.280 ;
        RECT 543.450 2.390 543.990 4.280 ;
        RECT 544.830 2.390 545.370 4.280 ;
        RECT 546.210 2.390 546.750 4.280 ;
        RECT 547.590 2.390 548.130 4.280 ;
        RECT 548.970 2.390 549.970 4.280 ;
        RECT 550.810 2.390 551.350 4.280 ;
        RECT 552.190 2.390 552.730 4.280 ;
        RECT 553.570 2.390 554.110 4.280 ;
        RECT 554.950 2.390 555.490 4.280 ;
        RECT 556.330 2.390 556.870 4.280 ;
        RECT 557.710 2.390 558.710 4.280 ;
        RECT 559.550 2.390 560.090 4.280 ;
        RECT 560.930 2.390 561.470 4.280 ;
        RECT 562.310 2.390 562.850 4.280 ;
        RECT 563.690 2.390 564.230 4.280 ;
        RECT 565.070 2.390 565.610 4.280 ;
        RECT 566.450 2.390 567.450 4.280 ;
        RECT 568.290 2.390 568.830 4.280 ;
        RECT 569.670 2.390 570.210 4.280 ;
        RECT 571.050 2.390 571.590 4.280 ;
        RECT 572.430 2.390 572.970 4.280 ;
        RECT 573.810 2.390 574.350 4.280 ;
        RECT 575.190 2.390 576.190 4.280 ;
        RECT 577.030 2.390 577.570 4.280 ;
        RECT 578.410 2.390 578.950 4.280 ;
        RECT 579.790 2.390 580.330 4.280 ;
        RECT 581.170 2.390 581.710 4.280 ;
        RECT 582.550 2.390 583.090 4.280 ;
        RECT 583.930 2.390 584.930 4.280 ;
        RECT 585.770 2.390 586.310 4.280 ;
        RECT 587.150 2.390 587.690 4.280 ;
        RECT 588.530 2.390 589.070 4.280 ;
        RECT 589.910 2.390 590.450 4.280 ;
        RECT 591.290 2.390 591.830 4.280 ;
        RECT 592.670 2.390 593.670 4.280 ;
        RECT 594.510 2.390 595.050 4.280 ;
        RECT 595.890 2.390 596.430 4.280 ;
        RECT 597.270 2.390 597.810 4.280 ;
        RECT 598.650 2.390 599.190 4.280 ;
        RECT 600.030 2.390 601.030 4.280 ;
        RECT 601.870 2.390 602.410 4.280 ;
        RECT 603.250 2.390 603.790 4.280 ;
        RECT 604.630 2.390 605.170 4.280 ;
        RECT 606.010 2.390 606.550 4.280 ;
        RECT 607.390 2.390 607.930 4.280 ;
        RECT 608.770 2.390 609.770 4.280 ;
        RECT 610.610 2.390 611.150 4.280 ;
        RECT 611.990 2.390 612.530 4.280 ;
        RECT 613.370 2.390 613.910 4.280 ;
        RECT 614.750 2.390 615.290 4.280 ;
        RECT 616.130 2.390 616.670 4.280 ;
        RECT 617.510 2.390 618.510 4.280 ;
        RECT 619.350 2.390 619.890 4.280 ;
        RECT 620.730 2.390 621.270 4.280 ;
        RECT 622.110 2.390 622.650 4.280 ;
        RECT 623.490 2.390 624.030 4.280 ;
        RECT 624.870 2.390 625.410 4.280 ;
        RECT 626.250 2.390 627.250 4.280 ;
        RECT 628.090 2.390 628.630 4.280 ;
        RECT 629.470 2.390 630.010 4.280 ;
        RECT 630.850 2.390 631.390 4.280 ;
        RECT 632.230 2.390 632.770 4.280 ;
        RECT 633.610 2.390 634.150 4.280 ;
        RECT 634.990 2.390 635.990 4.280 ;
        RECT 636.830 2.390 637.370 4.280 ;
        RECT 638.210 2.390 638.750 4.280 ;
        RECT 639.590 2.390 640.130 4.280 ;
        RECT 640.970 2.390 641.510 4.280 ;
        RECT 642.350 2.390 642.890 4.280 ;
        RECT 643.730 2.390 644.730 4.280 ;
        RECT 645.570 2.390 646.110 4.280 ;
        RECT 646.950 2.390 647.490 4.280 ;
        RECT 648.330 2.390 648.870 4.280 ;
        RECT 649.710 2.390 650.250 4.280 ;
        RECT 651.090 2.390 651.630 4.280 ;
        RECT 652.470 2.390 653.470 4.280 ;
        RECT 654.310 2.390 654.850 4.280 ;
        RECT 655.690 2.390 656.230 4.280 ;
        RECT 657.070 2.390 657.610 4.280 ;
        RECT 658.450 2.390 658.990 4.280 ;
        RECT 659.830 2.390 660.370 4.280 ;
        RECT 661.210 2.390 662.210 4.280 ;
        RECT 663.050 2.390 663.590 4.280 ;
        RECT 664.430 2.390 664.970 4.280 ;
        RECT 665.810 2.390 666.350 4.280 ;
        RECT 667.190 2.390 667.730 4.280 ;
        RECT 668.570 2.390 669.110 4.280 ;
        RECT 669.950 2.390 670.950 4.280 ;
        RECT 671.790 2.390 672.330 4.280 ;
        RECT 673.170 2.390 673.710 4.280 ;
        RECT 674.550 2.390 675.090 4.280 ;
        RECT 675.930 2.390 676.470 4.280 ;
        RECT 677.310 2.390 678.310 4.280 ;
        RECT 679.150 2.390 679.690 4.280 ;
        RECT 680.530 2.390 681.070 4.280 ;
        RECT 681.910 2.390 682.450 4.280 ;
        RECT 683.290 2.390 683.830 4.280 ;
        RECT 684.670 2.390 685.210 4.280 ;
        RECT 686.050 2.390 687.050 4.280 ;
        RECT 687.890 2.390 688.430 4.280 ;
        RECT 689.270 2.390 689.810 4.280 ;
        RECT 690.650 2.390 691.190 4.280 ;
        RECT 692.030 2.390 692.570 4.280 ;
        RECT 693.410 2.390 693.950 4.280 ;
        RECT 694.790 2.390 695.790 4.280 ;
        RECT 696.630 2.390 697.170 4.280 ;
        RECT 698.010 2.390 698.550 4.280 ;
        RECT 699.390 2.390 699.930 4.280 ;
        RECT 700.770 2.390 701.310 4.280 ;
        RECT 702.150 2.390 702.690 4.280 ;
        RECT 703.530 2.390 704.530 4.280 ;
        RECT 705.370 2.390 705.910 4.280 ;
        RECT 706.750 2.390 707.290 4.280 ;
        RECT 708.130 2.390 708.670 4.280 ;
        RECT 709.510 2.390 710.050 4.280 ;
        RECT 710.890 2.390 711.430 4.280 ;
        RECT 712.270 2.390 713.270 4.280 ;
        RECT 714.110 2.390 714.650 4.280 ;
        RECT 715.490 2.390 716.030 4.280 ;
        RECT 716.870 2.390 717.410 4.280 ;
        RECT 718.250 2.390 718.790 4.280 ;
        RECT 719.630 2.390 720.170 4.280 ;
        RECT 721.010 2.390 722.010 4.280 ;
        RECT 722.850 2.390 723.390 4.280 ;
        RECT 724.230 2.390 724.770 4.280 ;
        RECT 725.610 2.390 726.150 4.280 ;
        RECT 726.990 2.390 727.530 4.280 ;
        RECT 728.370 2.390 728.910 4.280 ;
        RECT 729.750 2.390 730.750 4.280 ;
        RECT 731.590 2.390 732.130 4.280 ;
        RECT 732.970 2.390 733.510 4.280 ;
        RECT 734.350 2.390 734.890 4.280 ;
        RECT 735.730 2.390 736.270 4.280 ;
        RECT 737.110 2.390 737.650 4.280 ;
        RECT 738.490 2.390 739.490 4.280 ;
        RECT 740.330 2.390 740.870 4.280 ;
        RECT 741.710 2.390 742.250 4.280 ;
        RECT 743.090 2.390 743.630 4.280 ;
        RECT 744.470 2.390 745.010 4.280 ;
        RECT 745.850 2.390 746.390 4.280 ;
        RECT 747.230 2.390 748.230 4.280 ;
        RECT 749.070 2.390 749.610 4.280 ;
        RECT 750.450 2.390 750.990 4.280 ;
        RECT 751.830 2.390 752.370 4.280 ;
        RECT 753.210 2.390 753.750 4.280 ;
        RECT 754.590 2.390 755.590 4.280 ;
        RECT 756.430 2.390 756.970 4.280 ;
        RECT 757.810 2.390 758.350 4.280 ;
        RECT 759.190 2.390 759.730 4.280 ;
        RECT 760.570 2.390 761.110 4.280 ;
        RECT 761.950 2.390 762.490 4.280 ;
        RECT 763.330 2.390 764.330 4.280 ;
        RECT 765.170 2.390 765.710 4.280 ;
        RECT 766.550 2.390 767.090 4.280 ;
        RECT 767.930 2.390 768.470 4.280 ;
        RECT 769.310 2.390 769.850 4.280 ;
        RECT 770.690 2.390 771.230 4.280 ;
        RECT 772.070 2.390 773.070 4.280 ;
        RECT 773.910 2.390 774.450 4.280 ;
        RECT 775.290 2.390 775.830 4.280 ;
        RECT 776.670 2.390 777.210 4.280 ;
        RECT 778.050 2.390 778.590 4.280 ;
        RECT 779.430 2.390 779.970 4.280 ;
        RECT 780.810 2.390 781.810 4.280 ;
        RECT 782.650 2.390 783.190 4.280 ;
        RECT 784.030 2.390 784.570 4.280 ;
        RECT 785.410 2.390 785.950 4.280 ;
        RECT 786.790 2.390 787.330 4.280 ;
        RECT 788.170 2.390 788.710 4.280 ;
        RECT 789.550 2.390 790.550 4.280 ;
        RECT 791.390 2.390 791.930 4.280 ;
        RECT 792.770 2.390 793.310 4.280 ;
        RECT 794.150 2.390 794.690 4.280 ;
        RECT 795.530 2.390 796.070 4.280 ;
        RECT 796.910 2.390 797.450 4.280 ;
        RECT 798.290 2.390 799.290 4.280 ;
        RECT 800.130 2.390 800.670 4.280 ;
        RECT 801.510 2.390 802.050 4.280 ;
        RECT 802.890 2.390 803.430 4.280 ;
        RECT 804.270 2.390 804.810 4.280 ;
        RECT 805.650 2.390 806.190 4.280 ;
        RECT 807.030 2.390 808.030 4.280 ;
        RECT 808.870 2.390 809.410 4.280 ;
        RECT 810.250 2.390 810.790 4.280 ;
        RECT 811.630 2.390 812.170 4.280 ;
        RECT 813.010 2.390 813.550 4.280 ;
        RECT 814.390 2.390 814.930 4.280 ;
        RECT 815.770 2.390 816.770 4.280 ;
        RECT 817.610 2.390 818.150 4.280 ;
        RECT 818.990 2.390 819.530 4.280 ;
        RECT 820.370 2.390 820.910 4.280 ;
        RECT 821.750 2.390 822.290 4.280 ;
        RECT 823.130 2.390 823.770 4.280 ;
      LAYER met3 ;
        RECT 4.000 827.240 819.500 827.385 ;
        RECT 4.400 826.520 819.500 827.240 ;
        RECT 4.400 825.840 823.795 826.520 ;
        RECT 4.000 814.320 823.795 825.840 ;
        RECT 4.000 812.920 819.500 814.320 ;
        RECT 4.000 812.280 823.795 812.920 ;
        RECT 4.400 810.880 823.795 812.280 ;
        RECT 4.000 800.720 823.795 810.880 ;
        RECT 4.000 799.320 819.500 800.720 ;
        RECT 4.000 797.320 823.795 799.320 ;
        RECT 4.400 795.920 823.795 797.320 ;
        RECT 4.000 787.120 823.795 795.920 ;
        RECT 4.000 785.720 819.500 787.120 ;
        RECT 4.000 782.360 823.795 785.720 ;
        RECT 4.400 780.960 823.795 782.360 ;
        RECT 4.000 773.520 823.795 780.960 ;
        RECT 4.000 772.120 819.500 773.520 ;
        RECT 4.000 767.400 823.795 772.120 ;
        RECT 4.400 766.000 823.795 767.400 ;
        RECT 4.000 759.920 823.795 766.000 ;
        RECT 4.000 758.520 819.500 759.920 ;
        RECT 4.000 752.440 823.795 758.520 ;
        RECT 4.400 751.040 823.795 752.440 ;
        RECT 4.000 746.320 823.795 751.040 ;
        RECT 4.000 744.920 819.500 746.320 ;
        RECT 4.000 737.480 823.795 744.920 ;
        RECT 4.400 736.080 823.795 737.480 ;
        RECT 4.000 732.720 823.795 736.080 ;
        RECT 4.000 731.320 819.500 732.720 ;
        RECT 4.000 722.520 823.795 731.320 ;
        RECT 4.400 721.120 823.795 722.520 ;
        RECT 4.000 718.440 823.795 721.120 ;
        RECT 4.000 717.040 819.500 718.440 ;
        RECT 4.000 707.560 823.795 717.040 ;
        RECT 4.400 706.160 823.795 707.560 ;
        RECT 4.000 704.840 823.795 706.160 ;
        RECT 4.000 703.440 819.500 704.840 ;
        RECT 4.000 692.600 823.795 703.440 ;
        RECT 4.400 691.240 823.795 692.600 ;
        RECT 4.400 691.200 819.500 691.240 ;
        RECT 4.000 689.840 819.500 691.200 ;
        RECT 4.000 677.640 823.795 689.840 ;
        RECT 4.400 676.240 819.500 677.640 ;
        RECT 4.000 664.040 823.795 676.240 ;
        RECT 4.000 663.360 819.500 664.040 ;
        RECT 4.400 662.640 819.500 663.360 ;
        RECT 4.400 661.960 823.795 662.640 ;
        RECT 4.000 650.440 823.795 661.960 ;
        RECT 4.000 649.040 819.500 650.440 ;
        RECT 4.000 648.400 823.795 649.040 ;
        RECT 4.400 647.000 823.795 648.400 ;
        RECT 4.000 636.840 823.795 647.000 ;
        RECT 4.000 635.440 819.500 636.840 ;
        RECT 4.000 633.440 823.795 635.440 ;
        RECT 4.400 632.040 823.795 633.440 ;
        RECT 4.000 623.240 823.795 632.040 ;
        RECT 4.000 621.840 819.500 623.240 ;
        RECT 4.000 618.480 823.795 621.840 ;
        RECT 4.400 617.080 823.795 618.480 ;
        RECT 4.000 609.640 823.795 617.080 ;
        RECT 4.000 608.240 819.500 609.640 ;
        RECT 4.000 603.520 823.795 608.240 ;
        RECT 4.400 602.120 823.795 603.520 ;
        RECT 4.000 595.360 823.795 602.120 ;
        RECT 4.000 593.960 819.500 595.360 ;
        RECT 4.000 588.560 823.795 593.960 ;
        RECT 4.400 587.160 823.795 588.560 ;
        RECT 4.000 581.760 823.795 587.160 ;
        RECT 4.000 580.360 819.500 581.760 ;
        RECT 4.000 573.600 823.795 580.360 ;
        RECT 4.400 572.200 823.795 573.600 ;
        RECT 4.000 568.160 823.795 572.200 ;
        RECT 4.000 566.760 819.500 568.160 ;
        RECT 4.000 558.640 823.795 566.760 ;
        RECT 4.400 557.240 823.795 558.640 ;
        RECT 4.000 554.560 823.795 557.240 ;
        RECT 4.000 553.160 819.500 554.560 ;
        RECT 4.000 543.680 823.795 553.160 ;
        RECT 4.400 542.280 823.795 543.680 ;
        RECT 4.000 540.960 823.795 542.280 ;
        RECT 4.000 539.560 819.500 540.960 ;
        RECT 4.000 528.720 823.795 539.560 ;
        RECT 4.400 527.360 823.795 528.720 ;
        RECT 4.400 527.320 819.500 527.360 ;
        RECT 4.000 525.960 819.500 527.320 ;
        RECT 4.000 513.760 823.795 525.960 ;
        RECT 4.400 512.360 819.500 513.760 ;
        RECT 4.000 500.160 823.795 512.360 ;
        RECT 4.000 499.480 819.500 500.160 ;
        RECT 4.400 498.760 819.500 499.480 ;
        RECT 4.400 498.080 823.795 498.760 ;
        RECT 4.000 486.560 823.795 498.080 ;
        RECT 4.000 485.160 819.500 486.560 ;
        RECT 4.000 484.520 823.795 485.160 ;
        RECT 4.400 483.120 823.795 484.520 ;
        RECT 4.000 472.280 823.795 483.120 ;
        RECT 4.000 470.880 819.500 472.280 ;
        RECT 4.000 469.560 823.795 470.880 ;
        RECT 4.400 468.160 823.795 469.560 ;
        RECT 4.000 458.680 823.795 468.160 ;
        RECT 4.000 457.280 819.500 458.680 ;
        RECT 4.000 454.600 823.795 457.280 ;
        RECT 4.400 453.200 823.795 454.600 ;
        RECT 4.000 445.080 823.795 453.200 ;
        RECT 4.000 443.680 819.500 445.080 ;
        RECT 4.000 439.640 823.795 443.680 ;
        RECT 4.400 438.240 823.795 439.640 ;
        RECT 4.000 431.480 823.795 438.240 ;
        RECT 4.000 430.080 819.500 431.480 ;
        RECT 4.000 424.680 823.795 430.080 ;
        RECT 4.400 423.280 823.795 424.680 ;
        RECT 4.000 417.880 823.795 423.280 ;
        RECT 4.000 416.480 819.500 417.880 ;
        RECT 4.000 409.720 823.795 416.480 ;
        RECT 4.400 408.320 823.795 409.720 ;
        RECT 4.000 404.280 823.795 408.320 ;
        RECT 4.000 402.880 819.500 404.280 ;
        RECT 4.000 394.760 823.795 402.880 ;
        RECT 4.400 393.360 823.795 394.760 ;
        RECT 4.000 390.680 823.795 393.360 ;
        RECT 4.000 389.280 819.500 390.680 ;
        RECT 4.000 379.800 823.795 389.280 ;
        RECT 4.400 378.400 823.795 379.800 ;
        RECT 4.000 377.080 823.795 378.400 ;
        RECT 4.000 375.680 819.500 377.080 ;
        RECT 4.000 364.840 823.795 375.680 ;
        RECT 4.400 363.440 823.795 364.840 ;
        RECT 4.000 362.800 823.795 363.440 ;
        RECT 4.000 361.400 819.500 362.800 ;
        RECT 4.000 349.880 823.795 361.400 ;
        RECT 4.400 349.200 823.795 349.880 ;
        RECT 4.400 348.480 819.500 349.200 ;
        RECT 4.000 347.800 819.500 348.480 ;
        RECT 4.000 335.600 823.795 347.800 ;
        RECT 4.400 334.200 819.500 335.600 ;
        RECT 4.000 322.000 823.795 334.200 ;
        RECT 4.000 320.640 819.500 322.000 ;
        RECT 4.400 320.600 819.500 320.640 ;
        RECT 4.400 319.240 823.795 320.600 ;
        RECT 4.000 308.400 823.795 319.240 ;
        RECT 4.000 307.000 819.500 308.400 ;
        RECT 4.000 305.680 823.795 307.000 ;
        RECT 4.400 304.280 823.795 305.680 ;
        RECT 4.000 294.800 823.795 304.280 ;
        RECT 4.000 293.400 819.500 294.800 ;
        RECT 4.000 290.720 823.795 293.400 ;
        RECT 4.400 289.320 823.795 290.720 ;
        RECT 4.000 281.200 823.795 289.320 ;
        RECT 4.000 279.800 819.500 281.200 ;
        RECT 4.000 275.760 823.795 279.800 ;
        RECT 4.400 274.360 823.795 275.760 ;
        RECT 4.000 267.600 823.795 274.360 ;
        RECT 4.000 266.200 819.500 267.600 ;
        RECT 4.000 260.800 823.795 266.200 ;
        RECT 4.400 259.400 823.795 260.800 ;
        RECT 4.000 254.000 823.795 259.400 ;
        RECT 4.000 252.600 819.500 254.000 ;
        RECT 4.000 245.840 823.795 252.600 ;
        RECT 4.400 244.440 823.795 245.840 ;
        RECT 4.000 239.720 823.795 244.440 ;
        RECT 4.000 238.320 819.500 239.720 ;
        RECT 4.000 230.880 823.795 238.320 ;
        RECT 4.400 229.480 823.795 230.880 ;
        RECT 4.000 226.120 823.795 229.480 ;
        RECT 4.000 224.720 819.500 226.120 ;
        RECT 4.000 215.920 823.795 224.720 ;
        RECT 4.400 214.520 823.795 215.920 ;
        RECT 4.000 212.520 823.795 214.520 ;
        RECT 4.000 211.120 819.500 212.520 ;
        RECT 4.000 200.960 823.795 211.120 ;
        RECT 4.400 199.560 823.795 200.960 ;
        RECT 4.000 198.920 823.795 199.560 ;
        RECT 4.000 197.520 819.500 198.920 ;
        RECT 4.000 186.000 823.795 197.520 ;
        RECT 4.400 185.320 823.795 186.000 ;
        RECT 4.400 184.600 819.500 185.320 ;
        RECT 4.000 183.920 819.500 184.600 ;
        RECT 4.000 171.720 823.795 183.920 ;
        RECT 4.400 170.320 819.500 171.720 ;
        RECT 4.000 158.120 823.795 170.320 ;
        RECT 4.000 156.760 819.500 158.120 ;
        RECT 4.400 156.720 819.500 156.760 ;
        RECT 4.400 155.360 823.795 156.720 ;
        RECT 4.000 144.520 823.795 155.360 ;
        RECT 4.000 143.120 819.500 144.520 ;
        RECT 4.000 141.800 823.795 143.120 ;
        RECT 4.400 140.400 823.795 141.800 ;
        RECT 4.000 130.920 823.795 140.400 ;
        RECT 4.000 129.520 819.500 130.920 ;
        RECT 4.000 126.840 823.795 129.520 ;
        RECT 4.400 125.440 823.795 126.840 ;
        RECT 4.000 116.640 823.795 125.440 ;
        RECT 4.000 115.240 819.500 116.640 ;
        RECT 4.000 111.880 823.795 115.240 ;
        RECT 4.400 110.480 823.795 111.880 ;
        RECT 4.000 103.040 823.795 110.480 ;
        RECT 4.000 101.640 819.500 103.040 ;
        RECT 4.000 96.920 823.795 101.640 ;
        RECT 4.400 95.520 823.795 96.920 ;
        RECT 4.000 89.440 823.795 95.520 ;
        RECT 4.000 88.040 819.500 89.440 ;
        RECT 4.000 81.960 823.795 88.040 ;
        RECT 4.400 80.560 823.795 81.960 ;
        RECT 4.000 75.840 823.795 80.560 ;
        RECT 4.000 74.440 819.500 75.840 ;
        RECT 4.000 67.000 823.795 74.440 ;
        RECT 4.400 65.600 823.795 67.000 ;
        RECT 4.000 62.240 823.795 65.600 ;
        RECT 4.000 60.840 819.500 62.240 ;
        RECT 4.000 52.040 823.795 60.840 ;
        RECT 4.400 50.640 823.795 52.040 ;
        RECT 4.000 48.640 823.795 50.640 ;
        RECT 4.000 47.240 819.500 48.640 ;
        RECT 4.000 37.080 823.795 47.240 ;
        RECT 4.400 35.680 823.795 37.080 ;
        RECT 4.000 35.040 823.795 35.680 ;
        RECT 4.000 33.640 819.500 35.040 ;
        RECT 4.000 22.120 823.795 33.640 ;
        RECT 4.400 21.440 823.795 22.120 ;
        RECT 4.400 20.720 819.500 21.440 ;
        RECT 4.000 20.040 819.500 20.720 ;
        RECT 4.000 7.840 823.795 20.040 ;
        RECT 4.400 6.440 819.500 7.840 ;
        RECT 4.000 2.220 823.795 6.440 ;
      LAYER met4 ;
        RECT 15.935 10.240 20.640 820.585 ;
        RECT 23.040 10.240 97.440 820.585 ;
        RECT 99.840 10.240 174.240 820.585 ;
        RECT 176.640 10.240 251.040 820.585 ;
        RECT 253.440 10.240 327.840 820.585 ;
        RECT 330.240 10.240 404.640 820.585 ;
        RECT 407.040 10.240 481.440 820.585 ;
        RECT 483.840 10.240 558.240 820.585 ;
        RECT 560.640 10.240 635.040 820.585 ;
        RECT 637.440 10.240 711.840 820.585 ;
        RECT 714.240 10.240 788.640 820.585 ;
        RECT 791.040 10.240 815.745 820.585 ;
        RECT 15.935 2.215 815.745 10.240 ;
  END
END user_proj
END LIBRARY

