magic
tech sky130A
magscale 1 2
timestamp 1639392407
<< locali >>
rect 26157 697595 26191 699329
rect 36001 697663 36035 699329
rect 50905 697731 50939 699329
rect 95157 698343 95191 699329
rect 109877 698411 109911 699329
rect 124597 698547 124631 699329
rect 129473 698683 129507 699329
rect 139317 698615 139351 699329
rect 158821 698819 158855 699329
rect 168849 698887 168883 699329
rect 173725 698955 173759 699329
rect 178601 699023 178635 699329
rect 188445 699091 188479 699329
rect 213837 699295 213871 699397
rect 379529 699159 379563 699465
rect 438317 698751 438351 699465
rect 453037 698479 453071 699465
rect 521853 697799 521887 699465
rect 7481 527 7515 697
rect 240517 595 240551 697
rect 196817 391 196851 561
rect 212089 459 212123 561
rect 252385 595 252419 697
rect 307677 663 307711 765
rect 214481 459 214515 561
rect 270049 255 270083 561
rect 279525 255 279559 629
rect 280721 187 280755 561
rect 283113 323 283147 561
rect 310345 51 310379 561
rect 319729 51 319763 629
rect 321017 323 321051 629
rect 328469 255 328503 561
rect 335737 255 335771 629
rect 337393 629 337577 663
rect 337393 595 337427 629
rect 341809 595 341843 697
rect 342361 663 342395 765
rect 338681 119 338715 561
rect 338773 255 338807 357
rect 342177 255 342211 561
rect 347605 459 347639 561
rect 351285 391 351319 765
rect 359289 595 359323 833
rect 372905 663 372939 765
rect 355793 187 355827 357
rect 356345 323 356379 561
rect 358277 323 358311 493
rect 367753 187 367787 425
rect 368213 255 368247 629
rect 373181 595 373215 765
rect 379897 425 380081 459
rect 379897 391 379931 425
rect 380633 255 380667 901
rect 386521 663 386555 901
rect 388269 595 388303 833
rect 389925 595 389959 833
rect 389465 391 389499 561
rect 393237 391 393271 765
rect 395537 391 395571 697
rect 396273 527 396307 969
rect 397745 595 397779 901
rect 405657 663 405691 901
rect 408325 663 408359 969
rect 406853 629 407037 663
rect 414949 663 414983 969
rect 415225 663 415259 901
rect 397837 323 397871 425
rect 396457 187 396491 289
rect 400137 255 400171 629
rect 403081 187 403115 425
rect 406853 391 406887 629
rect 417249 119 417283 629
rect 417341 187 417375 561
rect 422401 527 422435 1037
rect 424977 765 425069 799
rect 423723 561 423873 595
rect 422493 51 422527 493
rect 424517 323 424551 493
rect 424977 255 425011 765
rect 427277 595 427311 969
rect 428013 595 428047 901
rect 428473 663 428507 833
rect 430589 527 430623 833
rect 431877 663 431911 969
rect 435557 663 435591 1037
rect 432061 119 432095 561
rect 432705 51 432739 289
rect 433383 221 433533 255
rect 438409 51 438443 765
rect 441537 595 441571 901
rect 443285 595 443319 697
rect 445033 595 445067 969
rect 446229 595 446263 765
rect 446689 595 446723 1037
rect 442641 323 442675 561
rect 447425 119 447459 561
rect 448253 527 448287 833
rect 448897 187 448931 833
rect 451289 663 451323 901
rect 454233 663 454267 1105
rect 449541 527 449575 629
rect 454509 595 454543 833
rect 455061 595 455095 1037
rect 452301 323 452335 561
rect 455705 391 455739 629
rect 457177 459 457211 765
rect 461317 595 461351 697
rect 463157 663 463191 901
rect 464905 663 464939 833
rect 464997 527 465031 629
rect 467205 527 467239 901
rect 468401 663 468435 1105
rect 468493 595 468527 697
rect 468677 697 468769 731
rect 468677 595 468711 697
rect 469229 663 469263 1105
rect 468493 561 468711 595
rect 469689 527 469723 833
rect 449081 289 449265 323
rect 449081 255 449115 289
rect 470885 51 470919 697
rect 474013 663 474047 1173
rect 476773 663 476807 901
rect 476957 119 476991 629
rect 479625 595 479659 765
rect 483121 595 483155 833
rect 483765 595 483799 1037
rect 479533 391 479567 493
rect 483949 459 483983 697
rect 484041 595 484075 1105
rect 486617 663 486651 901
rect 484961 255 484995 493
rect 489009 459 489043 1173
rect 491217 901 491401 935
rect 491125 459 491159 697
rect 491217 663 491251 901
rect 492137 663 492171 969
rect 493333 663 493367 1173
rect 497841 663 497875 1105
rect 498117 799 498151 1377
rect 499405 595 499439 1037
rect 499497 663 499531 1037
rect 502993 595 503027 1377
rect 504649 663 504683 1241
rect 485053 119 485087 425
rect 503453 187 503487 493
rect 501153 51 501187 153
rect 505201 51 505235 357
rect 507317 323 507351 969
rect 507961 663 507995 969
rect 508605 663 508639 1173
rect 509893 663 509927 1173
rect 513573 663 513607 1105
rect 512561 119 512595 561
rect 513941 187 513975 697
rect 514677 663 514711 901
rect 514769 663 514803 1037
rect 518265 663 518299 1105
rect 520749 663 520783 1241
rect 518357 527 518391 629
rect 522865 663 522899 1037
rect 523049 663 523083 833
rect 523969 663 524003 833
rect 524245 663 524279 969
rect 519461 391 519495 629
rect 526453 527 526487 1173
rect 530133 595 530167 765
rect 530225 663 530259 969
rect 531329 595 531363 901
rect 531881 663 531915 901
rect 534549 595 534583 1105
rect 538781 663 538815 1105
rect 539793 459 539827 1037
rect 540805 595 540839 833
rect 542001 595 542035 969
rect 542185 459 542219 765
rect 554605 663 554639 969
rect 555893 663 555927 1105
rect 556077 799 556111 1037
rect 542277 255 542311 561
rect 550557 323 550591 493
rect 555985 323 556019 697
rect 556077 391 556111 629
rect 558009 323 558043 969
rect 561137 799 561171 1173
rect 561229 595 561263 765
rect 561413 595 561447 1105
<< viali >>
rect 379529 699465 379563 699499
rect 213837 699397 213871 699431
rect 26157 699329 26191 699363
rect 36001 699329 36035 699363
rect 50905 699329 50939 699363
rect 95157 699329 95191 699363
rect 109877 699329 109911 699363
rect 124597 699329 124631 699363
rect 129473 699329 129507 699363
rect 129473 698649 129507 698683
rect 139317 699329 139351 699363
rect 158821 699329 158855 699363
rect 168849 699329 168883 699363
rect 173725 699329 173759 699363
rect 178601 699329 178635 699363
rect 188445 699329 188479 699363
rect 213837 699261 213871 699295
rect 379529 699125 379563 699159
rect 438317 699465 438351 699499
rect 188445 699057 188479 699091
rect 178601 698989 178635 699023
rect 173725 698921 173759 698955
rect 168849 698853 168883 698887
rect 158821 698785 158855 698819
rect 438317 698717 438351 698751
rect 453037 699465 453071 699499
rect 139317 698581 139351 698615
rect 124597 698513 124631 698547
rect 453037 698445 453071 698479
rect 521853 699465 521887 699499
rect 109877 698377 109911 698411
rect 95157 698309 95191 698343
rect 521853 697765 521887 697799
rect 50905 697697 50939 697731
rect 36001 697629 36035 697663
rect 26157 697561 26191 697595
rect 498117 1377 498151 1411
rect 474013 1173 474047 1207
rect 454233 1105 454267 1139
rect 422401 1037 422435 1071
rect 396273 969 396307 1003
rect 380633 901 380667 935
rect 359289 833 359323 867
rect 307677 765 307711 799
rect 7481 697 7515 731
rect 240517 697 240551 731
rect 7481 493 7515 527
rect 196817 561 196851 595
rect 212089 561 212123 595
rect 212089 425 212123 459
rect 214481 561 214515 595
rect 240517 561 240551 595
rect 252385 697 252419 731
rect 342361 765 342395 799
rect 341809 697 341843 731
rect 279525 629 279559 663
rect 307677 629 307711 663
rect 319729 629 319763 663
rect 252385 561 252419 595
rect 270049 561 270083 595
rect 214481 425 214515 459
rect 196817 357 196851 391
rect 270049 221 270083 255
rect 279525 221 279559 255
rect 280721 561 280755 595
rect 283113 561 283147 595
rect 283113 289 283147 323
rect 310345 561 310379 595
rect 280721 153 280755 187
rect 310345 17 310379 51
rect 321017 629 321051 663
rect 335737 629 335771 663
rect 321017 289 321051 323
rect 328469 561 328503 595
rect 328469 221 328503 255
rect 337577 629 337611 663
rect 342361 629 342395 663
rect 351285 765 351319 799
rect 337393 561 337427 595
rect 338681 561 338715 595
rect 341809 561 341843 595
rect 342177 561 342211 595
rect 335737 221 335771 255
rect 338773 357 338807 391
rect 338773 221 338807 255
rect 347605 561 347639 595
rect 347605 425 347639 459
rect 372905 765 372939 799
rect 356345 561 356379 595
rect 359289 561 359323 595
rect 368213 629 368247 663
rect 372905 629 372939 663
rect 373181 765 373215 799
rect 351285 357 351319 391
rect 355793 357 355827 391
rect 342177 221 342211 255
rect 356345 289 356379 323
rect 358277 493 358311 527
rect 358277 289 358311 323
rect 367753 425 367787 459
rect 355793 153 355827 187
rect 373181 561 373215 595
rect 380081 425 380115 459
rect 379897 357 379931 391
rect 368213 221 368247 255
rect 386521 901 386555 935
rect 386521 629 386555 663
rect 388269 833 388303 867
rect 389925 833 389959 867
rect 388269 561 388303 595
rect 389465 561 389499 595
rect 389925 561 389959 595
rect 393237 765 393271 799
rect 389465 357 389499 391
rect 393237 357 393271 391
rect 395537 697 395571 731
rect 408325 969 408359 1003
rect 397745 901 397779 935
rect 405657 901 405691 935
rect 397745 561 397779 595
rect 400137 629 400171 663
rect 405657 629 405691 663
rect 407037 629 407071 663
rect 408325 629 408359 663
rect 414949 969 414983 1003
rect 414949 629 414983 663
rect 415225 901 415259 935
rect 415225 629 415259 663
rect 417249 629 417283 663
rect 396273 493 396307 527
rect 395537 357 395571 391
rect 397837 425 397871 459
rect 380633 221 380667 255
rect 396457 289 396491 323
rect 397837 289 397871 323
rect 367753 153 367787 187
rect 400137 221 400171 255
rect 403081 425 403115 459
rect 396457 153 396491 187
rect 406853 357 406887 391
rect 403081 153 403115 187
rect 338681 85 338715 119
rect 417341 561 417375 595
rect 435557 1037 435591 1071
rect 427277 969 427311 1003
rect 425069 765 425103 799
rect 423689 561 423723 595
rect 423873 561 423907 595
rect 422401 493 422435 527
rect 422493 493 422527 527
rect 417341 153 417375 187
rect 417249 85 417283 119
rect 319729 17 319763 51
rect 424517 493 424551 527
rect 424517 289 424551 323
rect 431877 969 431911 1003
rect 427277 561 427311 595
rect 428013 901 428047 935
rect 428473 833 428507 867
rect 428473 629 428507 663
rect 430589 833 430623 867
rect 428013 561 428047 595
rect 431877 629 431911 663
rect 446689 1037 446723 1071
rect 445033 969 445067 1003
rect 441537 901 441571 935
rect 435557 629 435591 663
rect 438409 765 438443 799
rect 430589 493 430623 527
rect 432061 561 432095 595
rect 424977 221 425011 255
rect 432061 85 432095 119
rect 432705 289 432739 323
rect 422493 17 422527 51
rect 433349 221 433383 255
rect 433533 221 433567 255
rect 432705 17 432739 51
rect 443285 697 443319 731
rect 441537 561 441571 595
rect 442641 561 442675 595
rect 443285 561 443319 595
rect 445033 561 445067 595
rect 446229 765 446263 799
rect 446229 561 446263 595
rect 451289 901 451323 935
rect 448253 833 448287 867
rect 446689 561 446723 595
rect 447425 561 447459 595
rect 442641 289 442675 323
rect 448253 493 448287 527
rect 448897 833 448931 867
rect 449541 629 449575 663
rect 451289 629 451323 663
rect 468401 1105 468435 1139
rect 455061 1037 455095 1071
rect 454233 629 454267 663
rect 454509 833 454543 867
rect 449541 493 449575 527
rect 452301 561 452335 595
rect 454509 561 454543 595
rect 463157 901 463191 935
rect 457177 765 457211 799
rect 455061 561 455095 595
rect 455705 629 455739 663
rect 461317 697 461351 731
rect 467205 901 467239 935
rect 463157 629 463191 663
rect 464905 833 464939 867
rect 464905 629 464939 663
rect 464997 629 465031 663
rect 461317 561 461351 595
rect 464997 493 465031 527
rect 469229 1105 469263 1139
rect 468401 629 468435 663
rect 468493 697 468527 731
rect 468769 697 468803 731
rect 469229 629 469263 663
rect 469689 833 469723 867
rect 467205 493 467239 527
rect 469689 493 469723 527
rect 470885 697 470919 731
rect 457177 425 457211 459
rect 455705 357 455739 391
rect 449265 289 449299 323
rect 452301 289 452335 323
rect 449081 221 449115 255
rect 448897 153 448931 187
rect 447425 85 447459 119
rect 438409 17 438443 51
rect 489009 1173 489043 1207
rect 484041 1105 484075 1139
rect 483765 1037 483799 1071
rect 474013 629 474047 663
rect 476773 901 476807 935
rect 483121 833 483155 867
rect 479625 765 479659 799
rect 476773 629 476807 663
rect 476957 629 476991 663
rect 479625 561 479659 595
rect 483121 561 483155 595
rect 483765 561 483799 595
rect 483949 697 483983 731
rect 479533 493 479567 527
rect 486617 901 486651 935
rect 486617 629 486651 663
rect 484041 561 484075 595
rect 483949 425 483983 459
rect 484961 493 484995 527
rect 479533 357 479567 391
rect 493333 1173 493367 1207
rect 492137 969 492171 1003
rect 491401 901 491435 935
rect 484961 221 484995 255
rect 485053 425 485087 459
rect 489009 425 489043 459
rect 491125 697 491159 731
rect 491217 629 491251 663
rect 492137 629 492171 663
rect 493333 629 493367 663
rect 497841 1105 497875 1139
rect 502993 1377 503027 1411
rect 498117 765 498151 799
rect 499405 1037 499439 1071
rect 497841 629 497875 663
rect 499497 1037 499531 1071
rect 499497 629 499531 663
rect 499405 561 499439 595
rect 504649 1241 504683 1275
rect 520749 1241 520783 1275
rect 508605 1173 508639 1207
rect 504649 629 504683 663
rect 507317 969 507351 1003
rect 502993 561 503027 595
rect 491125 425 491159 459
rect 503453 493 503487 527
rect 476957 85 476991 119
rect 485053 85 485087 119
rect 501153 153 501187 187
rect 503453 153 503487 187
rect 505201 357 505235 391
rect 470885 17 470919 51
rect 501153 17 501187 51
rect 507961 969 507995 1003
rect 507961 629 507995 663
rect 508605 629 508639 663
rect 509893 1173 509927 1207
rect 509893 629 509927 663
rect 513573 1105 513607 1139
rect 518265 1105 518299 1139
rect 514769 1037 514803 1071
rect 514677 901 514711 935
rect 513573 629 513607 663
rect 513941 697 513975 731
rect 507317 289 507351 323
rect 512561 561 512595 595
rect 514677 629 514711 663
rect 514769 629 514803 663
rect 526453 1173 526487 1207
rect 518265 629 518299 663
rect 518357 629 518391 663
rect 518357 493 518391 527
rect 519461 629 519495 663
rect 520749 629 520783 663
rect 522865 1037 522899 1071
rect 524245 969 524279 1003
rect 522865 629 522899 663
rect 523049 833 523083 867
rect 523049 629 523083 663
rect 523969 833 524003 867
rect 523969 629 524003 663
rect 524245 629 524279 663
rect 561137 1173 561171 1207
rect 534549 1105 534583 1139
rect 530225 969 530259 1003
rect 530133 765 530167 799
rect 530225 629 530259 663
rect 531329 901 531363 935
rect 530133 561 530167 595
rect 531881 901 531915 935
rect 531881 629 531915 663
rect 531329 561 531363 595
rect 538781 1105 538815 1139
rect 555893 1105 555927 1139
rect 538781 629 538815 663
rect 539793 1037 539827 1071
rect 534549 561 534583 595
rect 526453 493 526487 527
rect 542001 969 542035 1003
rect 540805 833 540839 867
rect 540805 561 540839 595
rect 554605 969 554639 1003
rect 542001 561 542035 595
rect 542185 765 542219 799
rect 539793 425 539827 459
rect 554605 629 554639 663
rect 556077 1037 556111 1071
rect 556077 765 556111 799
rect 558009 969 558043 1003
rect 555893 629 555927 663
rect 555985 697 556019 731
rect 542185 425 542219 459
rect 542277 561 542311 595
rect 519461 357 519495 391
rect 550557 493 550591 527
rect 550557 289 550591 323
rect 556077 629 556111 663
rect 556077 357 556111 391
rect 555985 289 556019 323
rect 561413 1105 561447 1139
rect 561137 765 561171 799
rect 561229 765 561263 799
rect 561229 561 561263 595
rect 561413 561 561447 595
rect 558009 289 558043 323
rect 542277 221 542311 255
rect 513941 153 513975 187
rect 512561 85 512595 119
rect 505201 17 505235 51
<< metal1 >>
rect 271782 703808 271788 703860
rect 271840 703848 271846 703860
rect 364702 703848 364708 703860
rect 271840 703820 364708 703848
rect 271840 703808 271846 703820
rect 364702 703808 364708 703820
rect 364760 703808 364766 703860
rect 235442 703740 235448 703792
rect 235500 703780 235506 703792
rect 300854 703780 300860 703792
rect 235500 703752 300860 703780
rect 235500 703740 235506 703752
rect 300854 703740 300860 703752
rect 300912 703740 300918 703792
rect 257246 703672 257252 703724
rect 257304 703712 257310 703724
rect 394694 703712 394700 703724
rect 257304 703684 394700 703712
rect 257304 703672 257310 703684
rect 394694 703672 394700 703684
rect 394752 703672 394758 703724
rect 242434 703604 242440 703656
rect 242492 703644 242498 703656
rect 400858 703644 400864 703656
rect 242492 703616 400864 703644
rect 242492 703604 242498 703616
rect 400858 703604 400864 703616
rect 400916 703604 400922 703656
rect 170490 703536 170496 703588
rect 170548 703576 170554 703588
rect 315482 703576 315488 703588
rect 170548 703548 315488 703576
rect 170548 703536 170554 703548
rect 315482 703536 315488 703548
rect 315540 703536 315546 703588
rect 227622 703468 227628 703520
rect 227680 703508 227686 703520
rect 468478 703508 468484 703520
rect 227680 703480 468484 703508
rect 227680 703468 227686 703480
rect 468478 703468 468484 703480
rect 468536 703468 468542 703520
rect 105446 703400 105452 703452
rect 105504 703440 105510 703452
rect 330294 703440 330300 703452
rect 105504 703412 330300 703440
rect 105504 703400 105510 703412
rect 330294 703400 330300 703412
rect 330352 703400 330358 703452
rect 1486 703332 1492 703384
rect 1544 703372 1550 703384
rect 359734 703372 359740 703384
rect 1544 703344 359740 703372
rect 1544 703332 1550 703344
rect 359734 703332 359740 703344
rect 359792 703332 359798 703384
rect 212994 703264 213000 703316
rect 213052 703304 213058 703316
rect 576302 703304 576308 703316
rect 213052 703276 576308 703304
rect 213052 703264 213058 703276
rect 576302 703264 576308 703276
rect 576360 703264 576366 703316
rect 1578 703196 1584 703248
rect 1636 703236 1642 703248
rect 374454 703236 374460 703248
rect 1636 703208 374460 703236
rect 1636 703196 1642 703208
rect 374454 703196 374460 703208
rect 374512 703196 374518 703248
rect 198274 703128 198280 703180
rect 198332 703168 198338 703180
rect 575014 703168 575020 703180
rect 198332 703140 575020 703168
rect 198332 703128 198338 703140
rect 575014 703128 575020 703140
rect 575072 703128 575078 703180
rect 1670 703060 1676 703112
rect 1728 703100 1734 703112
rect 389174 703100 389180 703112
rect 1728 703072 389180 703100
rect 1728 703060 1734 703072
rect 389174 703060 389180 703072
rect 389232 703060 389238 703112
rect 183370 702992 183376 703044
rect 183428 703032 183434 703044
rect 573634 703032 573640 703044
rect 183428 703004 573640 703032
rect 183428 702992 183434 703004
rect 573634 702992 573640 703004
rect 573692 702992 573698 703044
rect 750 702924 756 702976
rect 808 702964 814 702976
rect 394142 702964 394148 702976
rect 808 702936 394148 702964
rect 808 702924 814 702936
rect 394142 702924 394148 702936
rect 394200 702924 394206 702976
rect 1854 702856 1860 702908
rect 1912 702896 1918 702908
rect 403894 702896 403900 702908
rect 1912 702868 403900 702896
rect 1912 702856 1918 702868
rect 403894 702856 403900 702868
rect 403952 702856 403958 702908
rect 2498 702788 2504 702840
rect 2556 702828 2562 702840
rect 462866 702828 462872 702840
rect 2556 702800 462872 702828
rect 2556 702788 2562 702800
rect 462866 702788 462872 702800
rect 462924 702788 462930 702840
rect 382 702720 388 702772
rect 440 702760 446 702772
rect 492674 702760 492680 702772
rect 440 702732 492680 702760
rect 440 702720 446 702732
rect 492674 702720 492680 702732
rect 492732 702720 492738 702772
rect 198 702652 204 702704
rect 256 702692 262 702704
rect 507118 702692 507124 702704
rect 256 702664 507124 702692
rect 256 702652 262 702664
rect 507118 702652 507124 702664
rect 507176 702652 507182 702704
rect 41046 702584 41052 702636
rect 41104 702624 41110 702636
rect 578878 702624 578884 702636
rect 41104 702596 578884 702624
rect 41104 702584 41110 702596
rect 578878 702584 578884 702596
rect 578936 702584 578942 702636
rect 2038 702516 2044 702568
rect 2096 702556 2102 702568
rect 551278 702556 551284 702568
rect 2096 702528 551284 702556
rect 2096 702516 2102 702528
rect 551278 702516 551284 702528
rect 551336 702516 551342 702568
rect 21450 702448 21456 702500
rect 21508 702488 21514 702500
rect 576118 702488 576124 702500
rect 21508 702460 576124 702488
rect 21508 702448 21514 702460
rect 576118 702448 576124 702460
rect 576176 702448 576182 702500
rect 70118 702380 70124 702432
rect 70176 702420 70182 702432
rect 573450 702420 573456 702432
rect 70176 702392 573456 702420
rect 70176 702380 70182 702392
rect 573450 702380 573456 702392
rect 573508 702380 573514 702432
rect 237098 702312 237104 702364
rect 237156 702352 237162 702364
rect 291838 702352 291844 702364
rect 237156 702324 291844 702352
rect 237156 702312 237162 702324
rect 291838 702312 291844 702324
rect 291896 702312 291902 702364
rect 134426 702244 134432 702296
rect 134484 702284 134490 702296
rect 266354 702284 266360 702296
rect 134484 702256 266360 702284
rect 134484 702244 134490 702256
rect 266354 702244 266360 702256
rect 266412 702244 266418 702296
rect 277394 702244 277400 702296
rect 277452 702284 277458 702296
rect 428458 702284 428464 702296
rect 277452 702256 428464 702284
rect 277452 702244 277458 702256
rect 428458 702244 428464 702256
rect 428516 702244 428522 702296
rect 144270 702176 144276 702228
rect 144328 702216 144334 702228
rect 324314 702216 324320 702228
rect 144328 702188 324320 702216
rect 144328 702176 144334 702188
rect 324314 702176 324320 702188
rect 324372 702176 324378 702228
rect 100018 702108 100024 702160
rect 100076 702148 100082 702160
rect 311986 702148 311992 702160
rect 100076 702120 311992 702148
rect 100076 702108 100082 702120
rect 311986 702108 311992 702120
rect 312044 702108 312050 702160
rect 119706 702040 119712 702092
rect 119764 702080 119770 702092
rect 340138 702080 340144 702092
rect 119764 702052 340144 702080
rect 119764 702040 119770 702052
rect 340138 702040 340144 702052
rect 340196 702040 340202 702092
rect 55766 701972 55772 702024
rect 55824 702012 55830 702024
rect 304994 702012 305000 702024
rect 55824 701984 305000 702012
rect 55824 701972 55830 701984
rect 304994 701972 305000 701984
rect 305052 701972 305058 702024
rect 338022 701972 338028 702024
rect 338080 702012 338086 702024
rect 482554 702012 482560 702024
rect 338080 701984 482560 702012
rect 338080 701972 338086 701984
rect 482554 701972 482560 701984
rect 482612 701972 482618 702024
rect 6638 701904 6644 701956
rect 6696 701944 6702 701956
rect 259362 701944 259368 701956
rect 6696 701916 259368 701944
rect 6696 701904 6702 701916
rect 259362 701904 259368 701916
rect 259420 701904 259426 701956
rect 280890 701904 280896 701956
rect 280948 701944 280954 701956
rect 467834 701944 467840 701956
rect 280948 701916 467840 701944
rect 280948 701904 280954 701916
rect 467834 701904 467840 701916
rect 467892 701904 467898 701956
rect 154022 701836 154028 701888
rect 154080 701876 154086 701888
rect 565354 701876 565360 701888
rect 154080 701848 565360 701876
rect 154080 701836 154086 701848
rect 565354 701836 565360 701848
rect 565412 701836 565418 701888
rect 163866 701768 163872 701820
rect 163924 701808 163930 701820
rect 577590 701808 577596 701820
rect 163924 701780 577596 701808
rect 163924 701768 163930 701780
rect 577590 701768 577596 701780
rect 577648 701768 577654 701820
rect 148962 701700 148968 701752
rect 149020 701740 149026 701752
rect 574922 701740 574928 701752
rect 149020 701712 574928 701740
rect 149020 701700 149026 701712
rect 574922 701700 574928 701712
rect 574980 701700 574986 701752
rect 566 701632 572 701684
rect 624 701672 630 701684
rect 443270 701672 443276 701684
rect 624 701644 443276 701672
rect 624 701632 630 701644
rect 443270 701632 443276 701644
rect 443328 701632 443334 701684
rect 114278 701564 114284 701616
rect 114336 701604 114342 701616
rect 574830 701604 574836 701616
rect 114336 701576 574836 701604
rect 114336 701564 114342 701576
rect 574830 701564 574836 701576
rect 574888 701564 574894 701616
rect 4430 701496 4436 701548
rect 4488 701536 4494 701548
rect 472710 701536 472716 701548
rect 4488 701508 472716 701536
rect 4488 701496 4494 701508
rect 472710 701496 472716 701508
rect 472768 701496 472774 701548
rect 90174 701428 90180 701480
rect 90232 701468 90238 701480
rect 566550 701468 566556 701480
rect 90232 701440 566556 701468
rect 90232 701428 90238 701440
rect 566550 701428 566556 701440
rect 566608 701428 566614 701480
rect 2222 701360 2228 701412
rect 2280 701400 2286 701412
rect 487430 701400 487436 701412
rect 2280 701372 487436 701400
rect 2280 701360 2286 701372
rect 487430 701360 487436 701372
rect 487488 701360 487494 701412
rect 85298 701292 85304 701344
rect 85356 701332 85362 701344
rect 570690 701332 570696 701344
rect 85356 701304 570696 701332
rect 85356 701292 85362 701304
rect 570690 701292 570696 701304
rect 570748 701292 570754 701344
rect 75454 701224 75460 701276
rect 75512 701264 75518 701276
rect 570598 701264 570604 701276
rect 75512 701236 570604 701264
rect 75512 701224 75518 701236
rect 570598 701224 570604 701236
rect 570656 701224 570662 701276
rect 290 701156 296 701208
rect 348 701196 354 701208
rect 497274 701196 497280 701208
rect 348 701168 497280 701196
rect 348 701156 354 701168
rect 497274 701156 497280 701168
rect 497332 701156 497338 701208
rect 1302 701088 1308 701140
rect 1360 701128 1366 701140
rect 502334 701128 502340 701140
rect 1360 701100 502340 701128
rect 1360 701088 1366 701100
rect 502334 701088 502340 701100
rect 502392 701088 502398 701140
rect 556890 701088 556896 701140
rect 556948 701128 556954 701140
rect 564434 701128 564440 701140
rect 556948 701100 564440 701128
rect 556948 701088 556954 701100
rect 564434 701088 564440 701100
rect 564492 701088 564498 701140
rect 266998 701020 267004 701072
rect 267056 701060 267062 701072
rect 278590 701060 278596 701072
rect 267056 701032 278596 701060
rect 267056 701020 267062 701032
rect 278590 701020 278596 701032
rect 278648 701020 278654 701072
rect 292482 701020 292488 701072
rect 292540 701060 292546 701072
rect 295886 701060 295892 701072
rect 292540 701032 295892 701060
rect 292540 701020 292546 701032
rect 295886 701020 295892 701032
rect 295944 701020 295950 701072
rect 311894 701020 311900 701072
rect 311952 701060 311958 701072
rect 364610 701060 364616 701072
rect 311952 701032 364616 701060
rect 311952 701020 311958 701032
rect 364610 701020 364616 701032
rect 364668 701020 364674 701072
rect 468570 701020 468576 701072
rect 468628 701060 468634 701072
rect 511994 701060 512000 701072
rect 468628 701032 512000 701060
rect 468628 701020 468634 701032
rect 511994 701020 512000 701032
rect 512052 701020 512058 701072
rect 267642 700952 267648 701004
rect 267700 700992 267706 701004
rect 291378 700992 291384 701004
rect 267700 700964 291384 700992
rect 267700 700952 267706 700964
rect 291378 700952 291384 700964
rect 291436 700952 291442 701004
rect 291838 700952 291844 701004
rect 291896 700992 291902 701004
rect 543458 700992 543464 701004
rect 291896 700964 543464 700992
rect 291896 700952 291902 700964
rect 543458 700952 543464 700964
rect 543516 700952 543522 701004
rect 252278 700884 252284 700936
rect 252336 700924 252342 700936
rect 478506 700924 478512 700936
rect 252336 700896 478512 700924
rect 252336 700884 252342 700896
rect 478506 700884 478512 700896
rect 478564 700884 478570 700936
rect 89162 700816 89168 700868
rect 89220 700856 89226 700868
rect 340046 700856 340052 700868
rect 89220 700828 340052 700856
rect 89220 700816 89226 700828
rect 340046 700816 340052 700828
rect 340104 700816 340110 700868
rect 340138 700816 340144 700868
rect 340196 700856 340202 700868
rect 580626 700856 580632 700868
rect 340196 700828 580632 700856
rect 340196 700816 340202 700828
rect 580626 700816 580632 700828
rect 580684 700816 580690 700868
rect 3418 700748 3424 700800
rect 3476 700788 3482 700800
rect 262858 700788 262864 700800
rect 3476 700760 262864 700788
rect 3476 700748 3482 700760
rect 262858 700748 262864 700760
rect 262916 700748 262922 700800
rect 281350 700748 281356 700800
rect 281408 700788 281414 700800
rect 348786 700788 348792 700800
rect 281408 700760 348792 700788
rect 281408 700748 281414 700760
rect 348786 700748 348792 700760
rect 348844 700748 348850 700800
rect 468478 700748 468484 700800
rect 468536 700788 468542 700800
rect 559650 700788 559656 700800
rect 468536 700760 559656 700788
rect 468536 700748 468542 700760
rect 559650 700748 559656 700760
rect 559708 700748 559714 700800
rect 72970 700680 72976 700732
rect 73028 700720 73034 700732
rect 335354 700720 335360 700732
rect 73028 700692 335360 700720
rect 73028 700680 73034 700692
rect 335354 700680 335360 700692
rect 335412 700680 335418 700732
rect 336642 700680 336648 700732
rect 336700 700720 336706 700732
rect 580350 700720 580356 700732
rect 336700 700692 580356 700720
rect 336700 700680 336706 700692
rect 580350 700680 580356 700692
rect 580408 700680 580414 700732
rect 276842 700612 276848 700664
rect 276900 700652 276906 700664
rect 332502 700652 332508 700664
rect 276900 700624 332508 700652
rect 276900 700612 276906 700624
rect 332502 700612 332508 700624
rect 332560 700612 332566 700664
rect 3970 700544 3976 700596
rect 4028 700584 4034 700596
rect 280890 700584 280896 700596
rect 4028 700556 280896 700584
rect 4028 700544 4034 700556
rect 280890 700544 280896 700556
rect 280948 700544 280954 700596
rect 283834 700544 283840 700596
rect 283892 700584 283898 700596
rect 292482 700584 292488 700596
rect 283892 700556 292488 700584
rect 283892 700544 283898 700556
rect 292482 700544 292488 700556
rect 292540 700544 292546 700596
rect 298094 700544 298100 700596
rect 298152 700584 298158 700596
rect 300118 700584 300124 700596
rect 298152 700556 300124 700584
rect 298152 700544 298158 700556
rect 300118 700544 300124 700556
rect 300176 700544 300182 700596
rect 304994 700544 305000 700596
rect 305052 700584 305058 700596
rect 580442 700584 580448 700596
rect 305052 700556 580448 700584
rect 305052 700544 305058 700556
rect 580442 700544 580448 700556
rect 580500 700544 580506 700596
rect 232682 700476 232688 700528
rect 232740 700516 232746 700528
rect 527174 700516 527180 700528
rect 232740 700488 527180 700516
rect 232740 700476 232746 700488
rect 527174 700476 527180 700488
rect 527232 700476 527238 700528
rect 40494 700408 40500 700460
rect 40552 700448 40558 700460
rect 345198 700448 345204 700460
rect 40552 700420 345204 700448
rect 40552 700408 40558 700420
rect 345198 700408 345204 700420
rect 345256 700408 345262 700460
rect 400858 700408 400864 700460
rect 400916 700448 400922 700460
rect 494790 700448 494796 700460
rect 400916 700420 494796 700448
rect 400916 700408 400922 700420
rect 494790 700408 494796 700420
rect 494848 700408 494854 700460
rect 24302 700340 24308 700392
rect 24360 700380 24366 700392
rect 354950 700380 354956 700392
rect 24360 700352 354956 700380
rect 24360 700340 24366 700352
rect 354950 700340 354956 700352
rect 355008 700340 355014 700392
rect 394694 700340 394700 700392
rect 394752 700380 394758 700392
rect 429838 700380 429844 700392
rect 394752 700352 429844 700380
rect 394752 700340 394758 700352
rect 429838 700340 429844 700352
rect 429896 700340 429902 700392
rect 8110 700272 8116 700324
rect 8168 700312 8174 700324
rect 349890 700312 349896 700324
rect 8168 700284 349896 700312
rect 8168 700272 8174 700284
rect 349890 700272 349896 700284
rect 349948 700272 349954 700324
rect 247402 700204 247408 700256
rect 247460 700244 247466 700256
rect 462314 700244 462320 700256
rect 247460 700216 462320 700244
rect 247460 700204 247466 700216
rect 462314 700204 462320 700216
rect 462372 700204 462378 700256
rect 137830 700136 137836 700188
rect 137888 700176 137894 700188
rect 320772 700176 320778 700188
rect 137888 700148 320778 700176
rect 137888 700136 137894 700148
rect 320772 700136 320778 700148
rect 320830 700136 320836 700188
rect 324314 700136 324320 700188
rect 324372 700176 324378 700188
rect 580810 700176 580816 700188
rect 324372 700148 580816 700176
rect 324372 700136 324378 700148
rect 580810 700136 580816 700148
rect 580868 700136 580874 700188
rect 154114 700068 154120 700120
rect 154172 700108 154178 700120
rect 325648 700108 325654 700120
rect 154172 700080 325654 700108
rect 154172 700068 154178 700080
rect 325648 700068 325654 700080
rect 325706 700068 325712 700120
rect 262122 700000 262128 700052
rect 262180 700040 262186 700052
rect 397454 700040 397460 700052
rect 262180 700012 397460 700040
rect 262180 700000 262186 700012
rect 397454 700000 397460 700012
rect 397512 700000 397518 700052
rect 3326 699932 3332 699984
rect 3384 699972 3390 699984
rect 277302 699972 277308 699984
rect 3384 699944 277308 699972
rect 3384 699932 3390 699944
rect 277302 699932 277308 699944
rect 277360 699932 277366 699984
rect 278590 699932 278596 699984
rect 278648 699972 278654 699984
rect 413646 699972 413652 699984
rect 278648 699944 413652 699972
rect 278648 699932 278654 699944
rect 413646 699932 413652 699944
rect 413704 699932 413710 699984
rect 202690 699864 202696 699916
rect 202748 699904 202754 699916
rect 305730 699904 305736 699916
rect 202748 699876 305736 699904
rect 202748 699864 202754 699876
rect 305730 699864 305736 699876
rect 305788 699864 305794 699916
rect 311986 699864 311992 699916
rect 312044 699904 312050 699916
rect 580534 699904 580540 699916
rect 312044 699876 580540 699904
rect 312044 699864 312050 699876
rect 580534 699864 580540 699876
rect 580592 699864 580598 699916
rect 218974 699796 218980 699848
rect 219032 699836 219038 699848
rect 310606 699836 310612 699848
rect 219032 699808 310612 699836
rect 219032 699796 219038 699808
rect 310606 699796 310612 699808
rect 310664 699796 310670 699848
rect 4246 699728 4252 699780
rect 4304 699768 4310 699780
rect 369762 699768 369768 699780
rect 4304 699740 369768 699768
rect 4304 699728 4310 699740
rect 369762 699728 369768 699740
rect 369820 699728 369826 699780
rect 3786 699660 3792 699712
rect 3844 699700 3850 699712
rect 384298 699700 384304 699712
rect 3844 699672 384304 699700
rect 3844 699660 3850 699672
rect 384298 699660 384304 699672
rect 384356 699660 384362 699712
rect 3142 699592 3148 699644
rect 3200 699632 3206 699644
rect 311894 699632 311900 699644
rect 3200 699604 311900 699632
rect 3200 699592 3206 699604
rect 311894 699592 311900 699604
rect 311952 699592 311958 699644
rect 266354 699524 266360 699576
rect 266412 699564 266418 699576
rect 580718 699564 580724 699576
rect 266412 699536 580724 699564
rect 266412 699524 266418 699536
rect 580718 699524 580724 699536
rect 580776 699524 580782 699576
rect 3878 699456 3884 699508
rect 3936 699496 3942 699508
rect 338022 699496 338028 699508
rect 3936 699468 338028 699496
rect 3936 699456 3942 699468
rect 338022 699456 338028 699468
rect 338080 699456 338086 699508
rect 379514 699496 379520 699508
rect 379475 699468 379520 699496
rect 379514 699456 379520 699468
rect 379572 699456 379578 699508
rect 438302 699496 438308 699508
rect 438263 699468 438308 699496
rect 438302 699456 438308 699468
rect 438360 699456 438366 699508
rect 453022 699496 453028 699508
rect 452983 699468 453028 699496
rect 453022 699456 453028 699468
rect 453080 699456 453086 699508
rect 521838 699496 521844 699508
rect 521799 699468 521844 699496
rect 521838 699456 521844 699468
rect 521896 699456 521902 699508
rect 208118 699388 208124 699440
rect 208176 699428 208182 699440
rect 213825 699431 213883 699437
rect 213825 699428 213837 699431
rect 208176 699400 213837 699428
rect 208176 699388 208182 699400
rect 213825 699397 213837 699400
rect 213871 699397 213883 699431
rect 213825 699391 213883 699397
rect 222838 699388 222844 699440
rect 222896 699428 222902 699440
rect 572162 699428 572168 699440
rect 222896 699400 572168 699428
rect 222896 699388 222902 699400
rect 572162 699388 572168 699400
rect 572220 699388 572226 699440
rect 26142 699360 26148 699372
rect 26103 699332 26148 699360
rect 26142 699320 26148 699332
rect 26200 699320 26206 699372
rect 35986 699360 35992 699372
rect 35947 699332 35992 699360
rect 35986 699320 35992 699332
rect 36044 699320 36050 699372
rect 50890 699360 50896 699372
rect 50851 699332 50896 699360
rect 50890 699320 50896 699332
rect 50948 699320 50954 699372
rect 95142 699360 95148 699372
rect 95103 699332 95148 699360
rect 95142 699320 95148 699332
rect 95200 699320 95206 699372
rect 109862 699360 109868 699372
rect 109823 699332 109868 699360
rect 109862 699320 109868 699332
rect 109920 699320 109926 699372
rect 124582 699360 124588 699372
rect 124543 699332 124588 699360
rect 124582 699320 124588 699332
rect 124640 699320 124646 699372
rect 129458 699360 129464 699372
rect 129419 699332 129464 699360
rect 129458 699320 129464 699332
rect 129516 699320 129522 699372
rect 139302 699360 139308 699372
rect 139263 699332 139308 699360
rect 139302 699320 139308 699332
rect 139360 699320 139366 699372
rect 158806 699360 158812 699372
rect 158767 699332 158812 699360
rect 158806 699320 158812 699332
rect 158864 699320 158870 699372
rect 168834 699360 168840 699372
rect 168795 699332 168840 699360
rect 168834 699320 168840 699332
rect 168892 699320 168898 699372
rect 173710 699360 173716 699372
rect 173671 699332 173716 699360
rect 173710 699320 173716 699332
rect 173768 699320 173774 699372
rect 178586 699360 178592 699372
rect 178547 699332 178592 699360
rect 178586 699320 178592 699332
rect 178644 699320 178650 699372
rect 188430 699360 188436 699372
rect 188391 699332 188436 699360
rect 188430 699320 188436 699332
rect 188488 699320 188494 699372
rect 193214 699320 193220 699372
rect 193272 699360 193278 699372
rect 193272 699332 200114 699360
rect 193272 699320 193278 699332
rect 200086 699224 200114 699332
rect 202966 699320 202972 699372
rect 203024 699360 203030 699372
rect 563698 699360 563704 699372
rect 203024 699332 563704 699360
rect 203024 699320 203030 699332
rect 563698 699320 563704 699332
rect 563756 699320 563762 699372
rect 213825 699295 213883 699301
rect 213825 699261 213837 699295
rect 213871 699292 213883 699295
rect 570874 699292 570880 699304
rect 213871 699264 570880 699292
rect 213871 699261 213883 699264
rect 213825 699255 213883 699261
rect 570874 699252 570880 699264
rect 570932 699252 570938 699304
rect 567838 699224 567844 699236
rect 200086 699196 567844 699224
rect 567838 699184 567844 699196
rect 567896 699184 567902 699236
rect 842 699116 848 699168
rect 900 699156 906 699168
rect 379517 699159 379575 699165
rect 379517 699156 379529 699159
rect 900 699128 379529 699156
rect 900 699116 906 699128
rect 379517 699125 379529 699128
rect 379563 699125 379575 699159
rect 379517 699119 379575 699125
rect 188433 699091 188491 699097
rect 188433 699057 188445 699091
rect 188479 699088 188491 699091
rect 576210 699088 576216 699100
rect 188479 699060 576216 699088
rect 188479 699057 188491 699060
rect 188433 699051 188491 699057
rect 576210 699048 576216 699060
rect 576268 699048 576274 699100
rect 178589 699023 178647 699029
rect 178589 698989 178601 699023
rect 178635 699020 178647 699023
rect 569586 699020 569592 699032
rect 178635 698992 569592 699020
rect 178635 698989 178647 698992
rect 178589 698983 178647 698989
rect 569586 698980 569592 698992
rect 569644 698980 569650 699032
rect 173713 698955 173771 698961
rect 173713 698921 173725 698955
rect 173759 698952 173771 698955
rect 573542 698952 573548 698964
rect 173759 698924 573548 698952
rect 173759 698921 173771 698924
rect 173713 698915 173771 698921
rect 573542 698912 573548 698924
rect 573600 698912 573606 698964
rect 168837 698887 168895 698893
rect 168837 698853 168849 698887
rect 168883 698884 168895 698887
rect 569494 698884 569500 698896
rect 168883 698856 569500 698884
rect 168883 698853 168895 698856
rect 168837 698847 168895 698853
rect 569494 698844 569500 698856
rect 569552 698844 569558 698896
rect 158809 698819 158867 698825
rect 158809 698785 158821 698819
rect 158855 698816 158867 698819
rect 572070 698816 572076 698828
rect 158855 698788 572076 698816
rect 158855 698785 158867 698788
rect 158809 698779 158867 698785
rect 572070 698776 572076 698788
rect 572128 698776 572134 698828
rect 474 698708 480 698760
rect 532 698748 538 698760
rect 438305 698751 438363 698757
rect 438305 698748 438317 698751
rect 532 698720 438317 698748
rect 532 698708 538 698720
rect 438305 698717 438317 698720
rect 438351 698717 438363 698751
rect 438305 698711 438363 698717
rect 129461 698683 129519 698689
rect 129461 698649 129473 698683
rect 129507 698680 129519 698683
rect 566734 698680 566740 698692
rect 129507 698652 566740 698680
rect 129507 698649 129519 698652
rect 129461 698643 129519 698649
rect 566734 698640 566740 698652
rect 566792 698640 566798 698692
rect 139305 698615 139363 698621
rect 139305 698581 139317 698615
rect 139351 698612 139363 698615
rect 578970 698612 578976 698624
rect 139351 698584 578976 698612
rect 139351 698581 139363 698584
rect 139305 698575 139363 698581
rect 578970 698572 578976 698584
rect 579028 698572 579034 698624
rect 124585 698547 124643 698553
rect 124585 698513 124597 698547
rect 124631 698544 124643 698547
rect 570782 698544 570788 698556
rect 124631 698516 570788 698544
rect 124631 698513 124643 698516
rect 124585 698507 124643 698513
rect 570782 698504 570788 698516
rect 570840 698504 570846 698556
rect 2590 698436 2596 698488
rect 2648 698476 2654 698488
rect 453025 698479 453083 698485
rect 453025 698476 453037 698479
rect 2648 698448 453037 698476
rect 2648 698436 2654 698448
rect 453025 698445 453037 698448
rect 453071 698445 453083 698479
rect 453025 698439 453083 698445
rect 109865 698411 109923 698417
rect 109865 698377 109877 698411
rect 109911 698408 109923 698411
rect 569402 698408 569408 698420
rect 109911 698380 569408 698408
rect 109911 698377 109923 698380
rect 109865 698371 109923 698377
rect 569402 698368 569408 698380
rect 569460 698368 569466 698420
rect 95145 698343 95203 698349
rect 95145 698309 95157 698343
rect 95191 698340 95203 698343
rect 565170 698340 565176 698352
rect 95191 698312 565176 698340
rect 95191 698309 95203 698312
rect 95145 698303 95203 698309
rect 565170 698300 565176 698312
rect 565228 698300 565234 698352
rect 106 697756 112 697808
rect 164 697796 170 697808
rect 521841 697799 521899 697805
rect 521841 697796 521853 697799
rect 164 697768 521853 697796
rect 164 697756 170 697768
rect 521841 697765 521853 697768
rect 521887 697765 521899 697799
rect 521841 697759 521899 697765
rect 50893 697731 50951 697737
rect 50893 697697 50905 697731
rect 50939 697728 50951 697731
rect 573358 697728 573364 697740
rect 50939 697700 573364 697728
rect 50939 697697 50951 697700
rect 50893 697691 50951 697697
rect 573358 697688 573364 697700
rect 573416 697688 573422 697740
rect 35989 697663 36047 697669
rect 35989 697629 36001 697663
rect 36035 697660 36047 697663
rect 574738 697660 574744 697672
rect 36035 697632 574744 697660
rect 36035 697629 36047 697632
rect 35989 697623 36047 697629
rect 574738 697620 574744 697632
rect 574796 697620 574802 697672
rect 26145 697595 26203 697601
rect 26145 697561 26157 697595
rect 26191 697592 26203 697595
rect 569218 697592 569224 697604
rect 26191 697564 569224 697592
rect 26191 697561 26203 697564
rect 26145 697555 26203 697561
rect 569218 697552 569224 697564
rect 569276 697552 569282 697604
rect 572162 684428 572168 684480
rect 572220 684468 572226 684480
rect 580166 684468 580172 684480
rect 572220 684440 580172 684468
rect 572220 684428 572226 684440
rect 580166 684428 580172 684440
rect 580224 684428 580230 684480
rect 576302 671984 576308 672036
rect 576360 672024 576366 672036
rect 580166 672024 580172 672036
rect 576360 671996 580172 672024
rect 576360 671984 576366 671996
rect 580166 671984 580172 671996
rect 580224 671984 580230 672036
rect 563698 644376 563704 644428
rect 563756 644416 563762 644428
rect 580166 644416 580172 644428
rect 563756 644388 580172 644416
rect 563756 644376 563762 644388
rect 580166 644376 580172 644388
rect 580224 644376 580230 644428
rect 570874 632000 570880 632052
rect 570932 632040 570938 632052
rect 580166 632040 580172 632052
rect 570932 632012 580172 632040
rect 570932 632000 570938 632012
rect 580166 632000 580172 632012
rect 580224 632000 580230 632052
rect 575014 618196 575020 618248
rect 575072 618236 575078 618248
rect 580166 618236 580172 618248
rect 575072 618208 580172 618236
rect 575072 618196 575078 618208
rect 580166 618196 580172 618208
rect 580224 618196 580230 618248
rect 576210 591948 576216 592000
rect 576268 591988 576274 592000
rect 579982 591988 579988 592000
rect 576268 591960 579988 591988
rect 576268 591948 576274 591960
rect 579982 591948 579988 591960
rect 580040 591948 580046 592000
rect 567838 578144 567844 578196
rect 567896 578184 567902 578196
rect 579798 578184 579804 578196
rect 567896 578156 579804 578184
rect 567896 578144 567902 578156
rect 579798 578144 579804 578156
rect 579856 578144 579862 578196
rect 3786 565836 3792 565888
rect 3844 565876 3850 565888
rect 4338 565876 4344 565888
rect 3844 565848 4344 565876
rect 3844 565836 3850 565848
rect 4338 565836 4344 565848
rect 4396 565836 4402 565888
rect 573634 564340 573640 564392
rect 573692 564380 573698 564392
rect 580166 564380 580172 564392
rect 573692 564352 580172 564380
rect 573692 564340 573698 564352
rect 580166 564340 580172 564352
rect 580224 564340 580230 564392
rect 573542 538160 573548 538212
rect 573600 538200 573606 538212
rect 580166 538200 580172 538212
rect 573600 538172 580172 538200
rect 573600 538160 573606 538172
rect 580166 538160 580172 538172
rect 580224 538160 580230 538212
rect 569586 525716 569592 525768
rect 569644 525756 569650 525768
rect 580166 525756 580172 525768
rect 569644 525728 580172 525756
rect 569644 525716 569650 525728
rect 580166 525716 580172 525728
rect 580224 525716 580230 525768
rect 569494 511912 569500 511964
rect 569552 511952 569558 511964
rect 580166 511952 580172 511964
rect 569552 511924 580172 511952
rect 569552 511912 569558 511924
rect 580166 511912 580172 511924
rect 580224 511912 580230 511964
rect 3142 502256 3148 502308
rect 3200 502296 3206 502308
rect 4430 502296 4436 502308
rect 3200 502268 4436 502296
rect 3200 502256 3206 502268
rect 4430 502256 4436 502268
rect 4488 502256 4494 502308
rect 572070 485732 572076 485784
rect 572128 485772 572134 485784
rect 580166 485772 580172 485784
rect 572128 485744 580172 485772
rect 572128 485732 572134 485744
rect 580166 485732 580172 485744
rect 580224 485732 580230 485784
rect 577590 471928 577596 471980
rect 577648 471968 577654 471980
rect 580902 471968 580908 471980
rect 577648 471940 580908 471968
rect 577648 471928 577654 471940
rect 580902 471928 580908 471940
rect 580960 471928 580966 471980
rect 565354 458124 565360 458176
rect 565412 458164 565418 458176
rect 580166 458164 580172 458176
rect 565412 458136 580172 458164
rect 565412 458124 565418 458136
rect 580166 458124 580172 458136
rect 580224 458124 580230 458176
rect 574922 419432 574928 419484
rect 574980 419472 574986 419484
rect 580166 419472 580172 419484
rect 574980 419444 580172 419472
rect 574980 419432 574986 419444
rect 580166 419432 580172 419444
rect 580224 419432 580230 419484
rect 566734 379448 566740 379500
rect 566792 379488 566798 379500
rect 580166 379488 580172 379500
rect 566792 379460 580172 379488
rect 566792 379448 566798 379460
rect 580166 379448 580172 379460
rect 580224 379448 580230 379500
rect 570782 353200 570788 353252
rect 570840 353240 570846 353252
rect 580166 353240 580172 353252
rect 570840 353212 580172 353240
rect 570840 353200 570846 353212
rect 580166 353200 580172 353212
rect 580224 353200 580230 353252
rect 574830 325592 574836 325644
rect 574888 325632 574894 325644
rect 579982 325632 579988 325644
rect 574888 325604 579988 325632
rect 574888 325592 574894 325604
rect 579982 325592 579988 325604
rect 580040 325592 580046 325644
rect 569402 299412 569408 299464
rect 569460 299452 569466 299464
rect 580166 299452 580172 299464
rect 569460 299424 580172 299452
rect 569460 299412 569466 299424
rect 580166 299412 580172 299424
rect 580224 299412 580230 299464
rect 571978 259360 571984 259412
rect 572036 259400 572042 259412
rect 580166 259400 580172 259412
rect 572036 259372 580172 259400
rect 572036 259360 572042 259372
rect 580166 259360 580172 259372
rect 580224 259360 580230 259412
rect 1302 249704 1308 249756
rect 1360 249744 1366 249756
rect 2774 249744 2780 249756
rect 1360 249716 2780 249744
rect 1360 249704 1366 249716
rect 2774 249704 2780 249716
rect 2832 249704 2838 249756
rect 565170 245556 565176 245608
rect 565228 245596 565234 245608
rect 580166 245596 580172 245608
rect 565228 245568 580172 245596
rect 565228 245556 565234 245568
rect 580166 245556 580172 245568
rect 580224 245556 580230 245608
rect 570690 233180 570696 233232
rect 570748 233220 570754 233232
rect 579614 233220 579620 233232
rect 570748 233192 579620 233220
rect 570748 233180 570754 233192
rect 579614 233180 579620 233192
rect 579672 233180 579678 233232
rect 566550 219376 566556 219428
rect 566608 219416 566614 219428
rect 580166 219416 580172 219428
rect 566608 219388 580172 219416
rect 566608 219376 566614 219388
rect 580166 219376 580172 219388
rect 580224 219376 580230 219428
rect 566642 206932 566648 206984
rect 566700 206972 566706 206984
rect 580166 206972 580172 206984
rect 566700 206944 580172 206972
rect 566700 206932 566706 206944
rect 580166 206932 580172 206944
rect 580224 206932 580230 206984
rect 573450 193128 573456 193180
rect 573508 193168 573514 193180
rect 580166 193168 580172 193180
rect 573508 193140 580172 193168
rect 573508 193128 573514 193140
rect 580166 193128 580172 193140
rect 580224 193128 580230 193180
rect 570598 179324 570604 179376
rect 570656 179364 570662 179376
rect 580166 179364 580172 179376
rect 570656 179336 580172 179364
rect 570656 179324 570662 179336
rect 580166 179324 580172 179336
rect 580224 179324 580230 179376
rect 565262 166948 565268 167000
rect 565320 166988 565326 167000
rect 580166 166988 580172 167000
rect 565320 166960 580172 166988
rect 565320 166948 565326 166960
rect 580166 166948 580172 166960
rect 580224 166948 580230 167000
rect 569310 139340 569316 139392
rect 569368 139380 569374 139392
rect 580166 139380 580172 139392
rect 569368 139352 580172 139380
rect 569368 139340 569374 139352
rect 580166 139340 580172 139352
rect 580224 139340 580230 139392
rect 573358 126896 573364 126948
rect 573416 126936 573422 126948
rect 580166 126936 580172 126948
rect 573416 126908 580172 126936
rect 573416 126896 573422 126908
rect 580166 126896 580172 126908
rect 580224 126896 580230 126948
rect 577498 100648 577504 100700
rect 577556 100688 577562 100700
rect 579798 100688 579804 100700
rect 577556 100660 579804 100688
rect 577556 100648 577562 100660
rect 579798 100648 579804 100660
rect 579856 100648 579862 100700
rect 574738 86912 574744 86964
rect 574796 86952 574802 86964
rect 579614 86952 579620 86964
rect 574796 86924 579620 86952
rect 574796 86912 574802 86924
rect 579614 86912 579620 86924
rect 579672 86912 579678 86964
rect 569218 73108 569224 73160
rect 569276 73148 569282 73160
rect 580166 73148 580172 73160
rect 569276 73120 580172 73148
rect 569276 73108 569282 73120
rect 580166 73108 580172 73120
rect 580224 73108 580230 73160
rect 576118 46860 576124 46912
rect 576176 46900 576182 46912
rect 580166 46900 580172 46912
rect 576176 46872 580172 46900
rect 576176 46860 576182 46872
rect 580166 46860 580172 46872
rect 580224 46860 580230 46912
rect 566458 33056 566464 33108
rect 566516 33096 566522 33108
rect 580166 33096 580172 33108
rect 566516 33068 580172 33096
rect 566516 33056 566522 33068
rect 580166 33056 580172 33068
rect 580224 33056 580230 33108
rect 565078 20612 565084 20664
rect 565136 20652 565142 20664
rect 580166 20652 580172 20664
rect 565136 20624 580172 20652
rect 565136 20612 565142 20624
rect 580166 20612 580172 20624
rect 580224 20612 580230 20664
rect 563606 3136 563612 3188
rect 563664 3176 563670 3188
rect 569126 3176 569132 3188
rect 563664 3148 569132 3176
rect 563664 3136 563670 3148
rect 569126 3136 569132 3148
rect 569184 3136 569190 3188
rect 565906 3068 565912 3120
rect 565964 3108 565970 3120
rect 571518 3108 571524 3120
rect 565964 3080 571524 3108
rect 565964 3068 565970 3080
rect 571518 3068 571524 3080
rect 571576 3068 571582 3120
rect 563698 3000 563704 3052
rect 563756 3040 563762 3052
rect 583386 3040 583392 3052
rect 563756 3012 583392 3040
rect 563756 3000 563762 3012
rect 583386 3000 583392 3012
rect 583444 3000 583450 3052
rect 563514 2864 563520 2916
rect 563572 2904 563578 2916
rect 572714 2904 572720 2916
rect 563572 2876 572720 2904
rect 563572 2864 563578 2876
rect 572714 2864 572720 2876
rect 572772 2864 572778 2916
rect 569862 2796 569868 2848
rect 569920 2836 569926 2848
rect 576302 2836 576308 2848
rect 569920 2808 576308 2836
rect 569920 2796 569926 2808
rect 576302 2796 576308 2808
rect 576360 2796 576366 2848
rect 498105 1411 498163 1417
rect 498105 1377 498117 1411
rect 498151 1408 498163 1411
rect 502981 1411 503039 1417
rect 502981 1408 502993 1411
rect 498151 1380 502993 1408
rect 498151 1377 498163 1380
rect 498105 1371 498163 1377
rect 502981 1377 502993 1380
rect 503027 1377 503039 1411
rect 502981 1371 503039 1377
rect 3050 1300 3056 1352
rect 3108 1340 3114 1352
rect 564434 1340 564440 1352
rect 3108 1312 564440 1340
rect 3108 1300 3114 1312
rect 564434 1300 564440 1312
rect 564492 1300 564498 1352
rect 504637 1275 504695 1281
rect 504637 1241 504649 1275
rect 504683 1272 504695 1275
rect 520737 1275 520795 1281
rect 520737 1272 520749 1275
rect 504683 1244 520749 1272
rect 504683 1241 504695 1244
rect 504637 1235 504695 1241
rect 520737 1241 520749 1244
rect 520783 1241 520795 1275
rect 520737 1235 520795 1241
rect 474001 1207 474059 1213
rect 474001 1173 474013 1207
rect 474047 1204 474059 1207
rect 488997 1207 489055 1213
rect 488997 1204 489009 1207
rect 474047 1176 489009 1204
rect 474047 1173 474059 1176
rect 474001 1167 474059 1173
rect 488997 1173 489009 1176
rect 489043 1173 489055 1207
rect 488997 1167 489055 1173
rect 493321 1207 493379 1213
rect 493321 1173 493333 1207
rect 493367 1204 493379 1207
rect 508593 1207 508651 1213
rect 508593 1204 508605 1207
rect 493367 1176 508605 1204
rect 493367 1173 493379 1176
rect 493321 1167 493379 1173
rect 508593 1173 508605 1176
rect 508639 1173 508651 1207
rect 508593 1167 508651 1173
rect 509881 1207 509939 1213
rect 509881 1173 509893 1207
rect 509927 1204 509939 1207
rect 526441 1207 526499 1213
rect 526441 1204 526453 1207
rect 509927 1176 526453 1204
rect 509927 1173 509939 1176
rect 509881 1167 509939 1173
rect 526441 1173 526453 1176
rect 526487 1173 526499 1207
rect 526441 1167 526499 1173
rect 561125 1207 561183 1213
rect 561125 1173 561137 1207
rect 561171 1204 561183 1207
rect 566826 1204 566832 1216
rect 561171 1176 566832 1204
rect 561171 1173 561183 1176
rect 561125 1167 561183 1173
rect 566826 1164 566832 1176
rect 566884 1164 566890 1216
rect 454221 1139 454279 1145
rect 454221 1105 454233 1139
rect 454267 1136 454279 1139
rect 468389 1139 468447 1145
rect 468389 1136 468401 1139
rect 454267 1108 468401 1136
rect 454267 1105 454279 1108
rect 454221 1099 454279 1105
rect 468389 1105 468401 1108
rect 468435 1105 468447 1139
rect 468389 1099 468447 1105
rect 469217 1139 469275 1145
rect 469217 1105 469229 1139
rect 469263 1136 469275 1139
rect 484029 1139 484087 1145
rect 484029 1136 484041 1139
rect 469263 1108 484041 1136
rect 469263 1105 469275 1108
rect 469217 1099 469275 1105
rect 484029 1105 484041 1108
rect 484075 1105 484087 1139
rect 484029 1099 484087 1105
rect 497829 1139 497887 1145
rect 497829 1105 497841 1139
rect 497875 1136 497887 1139
rect 513561 1139 513619 1145
rect 513561 1136 513573 1139
rect 497875 1108 513573 1136
rect 497875 1105 497887 1108
rect 497829 1099 497887 1105
rect 513561 1105 513573 1108
rect 513607 1105 513619 1139
rect 513561 1099 513619 1105
rect 518253 1139 518311 1145
rect 518253 1105 518265 1139
rect 518299 1136 518311 1139
rect 534537 1139 534595 1145
rect 534537 1136 534549 1139
rect 518299 1108 534549 1136
rect 518299 1105 518311 1108
rect 518253 1099 518311 1105
rect 534537 1105 534549 1108
rect 534583 1105 534595 1139
rect 534537 1099 534595 1105
rect 538769 1139 538827 1145
rect 538769 1105 538781 1139
rect 538815 1136 538827 1139
rect 555881 1139 555939 1145
rect 555881 1136 555893 1139
rect 538815 1108 555893 1136
rect 538815 1105 538827 1108
rect 538769 1099 538827 1105
rect 555881 1105 555893 1108
rect 555927 1105 555939 1139
rect 555881 1099 555939 1105
rect 561401 1139 561459 1145
rect 561401 1105 561413 1139
rect 561447 1136 561459 1139
rect 580994 1136 581000 1148
rect 561447 1108 581000 1136
rect 561447 1105 561459 1108
rect 561401 1099 561459 1105
rect 580994 1096 581000 1108
rect 581052 1096 581058 1148
rect 422389 1071 422447 1077
rect 422389 1037 422401 1071
rect 422435 1068 422447 1071
rect 435545 1071 435603 1077
rect 435545 1068 435557 1071
rect 422435 1040 435557 1068
rect 422435 1037 422447 1040
rect 422389 1031 422447 1037
rect 435545 1037 435557 1040
rect 435591 1037 435603 1071
rect 435545 1031 435603 1037
rect 446677 1071 446735 1077
rect 446677 1037 446689 1071
rect 446723 1068 446735 1071
rect 455049 1071 455107 1077
rect 455049 1068 455061 1071
rect 446723 1040 455061 1068
rect 446723 1037 446735 1040
rect 446677 1031 446735 1037
rect 455049 1037 455061 1040
rect 455095 1037 455107 1071
rect 455049 1031 455107 1037
rect 483753 1071 483811 1077
rect 483753 1037 483765 1071
rect 483799 1068 483811 1071
rect 499393 1071 499451 1077
rect 499393 1068 499405 1071
rect 483799 1040 499405 1068
rect 483799 1037 483811 1040
rect 483753 1031 483811 1037
rect 499393 1037 499405 1040
rect 499439 1037 499451 1071
rect 499393 1031 499451 1037
rect 499485 1071 499543 1077
rect 499485 1037 499497 1071
rect 499531 1068 499543 1071
rect 514757 1071 514815 1077
rect 514757 1068 514769 1071
rect 499531 1040 514769 1068
rect 499531 1037 499543 1040
rect 499485 1031 499543 1037
rect 514757 1037 514769 1040
rect 514803 1037 514815 1071
rect 514757 1031 514815 1037
rect 522853 1071 522911 1077
rect 522853 1037 522865 1071
rect 522899 1068 522911 1071
rect 539781 1071 539839 1077
rect 539781 1068 539793 1071
rect 522899 1040 539793 1068
rect 522899 1037 522911 1040
rect 522853 1031 522911 1037
rect 539781 1037 539793 1040
rect 539827 1037 539839 1071
rect 556065 1071 556123 1077
rect 556065 1068 556077 1071
rect 539781 1031 539839 1037
rect 553366 1040 556077 1068
rect 396261 1003 396319 1009
rect 396261 969 396273 1003
rect 396307 1000 396319 1003
rect 408313 1003 408371 1009
rect 408313 1000 408325 1003
rect 396307 972 408325 1000
rect 396307 969 396319 972
rect 396261 963 396319 969
rect 408313 969 408325 972
rect 408359 969 408371 1003
rect 408313 963 408371 969
rect 414937 1003 414995 1009
rect 414937 969 414949 1003
rect 414983 1000 414995 1003
rect 427265 1003 427323 1009
rect 427265 1000 427277 1003
rect 414983 972 427277 1000
rect 414983 969 414995 972
rect 414937 963 414995 969
rect 427265 969 427277 972
rect 427311 969 427323 1003
rect 427265 963 427323 969
rect 431865 1003 431923 1009
rect 431865 969 431877 1003
rect 431911 1000 431923 1003
rect 445021 1003 445079 1009
rect 445021 1000 445033 1003
rect 431911 972 445033 1000
rect 431911 969 431923 972
rect 431865 963 431923 969
rect 445021 969 445033 972
rect 445067 969 445079 1003
rect 445021 963 445079 969
rect 492125 1003 492183 1009
rect 492125 969 492137 1003
rect 492171 1000 492183 1003
rect 507305 1003 507363 1009
rect 507305 1000 507317 1003
rect 492171 972 507317 1000
rect 492171 969 492183 972
rect 492125 963 492183 969
rect 507305 969 507317 972
rect 507351 969 507363 1003
rect 507305 963 507363 969
rect 507949 1003 508007 1009
rect 507949 969 507961 1003
rect 507995 1000 508007 1003
rect 524233 1003 524291 1009
rect 524233 1000 524245 1003
rect 507995 972 524245 1000
rect 507995 969 508007 972
rect 507949 963 508007 969
rect 524233 969 524245 972
rect 524279 969 524291 1003
rect 524233 963 524291 969
rect 530213 1003 530271 1009
rect 530213 969 530225 1003
rect 530259 1000 530271 1003
rect 541989 1003 542047 1009
rect 541989 1000 542001 1003
rect 530259 972 542001 1000
rect 530259 969 530271 972
rect 530213 963 530271 969
rect 541989 969 542001 972
rect 542035 969 542047 1003
rect 553366 1000 553394 1040
rect 556065 1037 556077 1040
rect 556111 1037 556123 1071
rect 563514 1068 563520 1080
rect 556065 1031 556123 1037
rect 557506 1040 563520 1068
rect 541989 963 542047 969
rect 551020 972 553394 1000
rect 554593 1003 554651 1009
rect 380621 935 380679 941
rect 380621 901 380633 935
rect 380667 932 380679 935
rect 386509 935 386567 941
rect 380667 904 382274 932
rect 380667 901 380679 904
rect 380621 895 380679 901
rect 359277 867 359335 873
rect 359277 833 359289 867
rect 359323 864 359335 867
rect 382246 864 382274 904
rect 386509 901 386521 935
rect 386555 932 386567 935
rect 397733 935 397791 941
rect 397733 932 397745 935
rect 386555 904 397745 932
rect 386555 901 386567 904
rect 386509 895 386567 901
rect 397733 901 397745 904
rect 397779 901 397791 935
rect 397733 895 397791 901
rect 405645 935 405703 941
rect 405645 901 405657 935
rect 405691 932 405703 935
rect 415213 935 415271 941
rect 415213 932 415225 935
rect 405691 904 415225 932
rect 405691 901 405703 904
rect 405645 895 405703 901
rect 415213 901 415225 904
rect 415259 901 415271 935
rect 415213 895 415271 901
rect 428001 935 428059 941
rect 428001 901 428013 935
rect 428047 932 428059 935
rect 441525 935 441583 941
rect 441525 932 441537 935
rect 428047 904 441537 932
rect 428047 901 428059 904
rect 428001 895 428059 901
rect 441525 901 441537 904
rect 441571 901 441583 935
rect 441525 895 441583 901
rect 451277 935 451335 941
rect 451277 901 451289 935
rect 451323 932 451335 935
rect 463145 935 463203 941
rect 463145 932 463157 935
rect 451323 904 463157 932
rect 451323 901 451335 904
rect 451277 895 451335 901
rect 463145 901 463157 904
rect 463191 901 463203 935
rect 463145 895 463203 901
rect 467193 935 467251 941
rect 467193 901 467205 935
rect 467239 932 467251 935
rect 476761 935 476819 941
rect 476761 932 476773 935
rect 467239 904 476773 932
rect 467239 901 467251 904
rect 467193 895 467251 901
rect 476761 901 476773 904
rect 476807 901 476819 935
rect 486605 935 486663 941
rect 486605 932 486617 935
rect 476761 895 476819 901
rect 478846 904 486617 932
rect 388257 867 388315 873
rect 388257 864 388269 867
rect 359323 836 369440 864
rect 382246 836 388269 864
rect 359323 833 359335 836
rect 359277 827 359335 833
rect 307665 799 307723 805
rect 307665 765 307677 799
rect 307711 796 307723 799
rect 342349 799 342407 805
rect 342349 796 342361 799
rect 307711 768 314654 796
rect 307711 765 307723 768
rect 307665 759 307723 765
rect 7469 731 7527 737
rect 7469 697 7481 731
rect 7515 728 7527 731
rect 240505 731 240563 737
rect 240505 728 240517 731
rect 7515 700 11560 728
rect 7515 697 7527 700
rect 7469 691 7527 697
rect 11532 672 11560 700
rect 237346 700 240517 728
rect 1670 620 1676 672
rect 1728 660 1734 672
rect 5350 660 5356 672
rect 1728 632 5356 660
rect 1728 620 1734 632
rect 5350 620 5356 632
rect 5408 620 5414 672
rect 6454 620 6460 672
rect 6512 660 6518 672
rect 10042 660 10048 672
rect 6512 632 10048 660
rect 6512 620 6518 632
rect 10042 620 10048 632
rect 10100 620 10106 672
rect 10152 632 11468 660
rect 566 552 572 604
rect 624 592 630 604
rect 4338 592 4344 604
rect 624 564 4344 592
rect 624 552 630 564
rect 4338 552 4344 564
rect 4396 552 4402 604
rect 5258 552 5264 604
rect 5316 592 5322 604
rect 8846 592 8852 604
rect 5316 564 8852 592
rect 5316 552 5322 564
rect 8846 552 8852 564
rect 8904 552 8910 604
rect 7466 524 7472 536
rect 7427 496 7472 524
rect 7466 484 7472 496
rect 7524 484 7530 536
rect 8570 484 8576 536
rect 8628 524 8634 536
rect 10152 524 10180 632
rect 11146 552 11152 604
rect 11204 552 11210 604
rect 11440 592 11468 632
rect 11514 620 11520 672
rect 11572 620 11578 672
rect 19426 620 19432 672
rect 19484 660 19490 672
rect 22370 660 22376 672
rect 19484 632 22376 660
rect 19484 620 19490 632
rect 22370 620 22376 632
rect 22428 620 22434 672
rect 24854 660 24860 672
rect 22480 632 24860 660
rect 11440 564 11836 592
rect 8628 496 10180 524
rect 11164 524 11192 552
rect 11808 524 11836 564
rect 12342 552 12348 604
rect 12400 592 12406 604
rect 15562 592 15568 604
rect 12400 564 15568 592
rect 12400 552 12406 564
rect 15562 552 15568 564
rect 15620 552 15626 604
rect 21818 552 21824 604
rect 21876 592 21882 604
rect 22480 592 22508 632
rect 24854 620 24860 632
rect 24912 620 24918 672
rect 25314 620 25320 672
rect 25372 660 25378 672
rect 28074 660 28080 672
rect 25372 632 28080 660
rect 25372 620 25378 632
rect 28074 620 28080 632
rect 28132 620 28138 672
rect 28718 620 28724 672
rect 28776 660 28782 672
rect 29178 660 29184 672
rect 28776 632 29184 660
rect 28776 620 28782 632
rect 29178 620 29184 632
rect 29236 620 29242 672
rect 31294 620 31300 672
rect 31352 660 31358 672
rect 33778 660 33784 672
rect 31352 632 33784 660
rect 31352 620 31358 632
rect 33778 620 33784 632
rect 33836 620 33842 672
rect 34790 620 34796 672
rect 34848 660 34854 672
rect 37274 660 37280 672
rect 34848 632 37280 660
rect 34848 620 34854 632
rect 37274 620 37280 632
rect 37332 620 37338 672
rect 38378 620 38384 672
rect 38436 660 38442 672
rect 38436 632 38654 660
rect 38436 620 38442 632
rect 21876 564 22508 592
rect 21876 552 21882 564
rect 23014 552 23020 604
rect 23072 592 23078 604
rect 25774 592 25780 604
rect 23072 564 25780 592
rect 23072 552 23078 564
rect 25774 552 25780 564
rect 25832 552 25838 604
rect 28810 552 28816 604
rect 28868 592 28874 604
rect 28868 564 29040 592
rect 28868 552 28874 564
rect 12618 524 12624 536
rect 11164 496 11284 524
rect 11808 496 12624 524
rect 8628 484 8634 496
rect 3234 416 3240 468
rect 3292 456 3298 468
rect 6638 456 6644 468
rect 3292 428 6644 456
rect 3292 416 3298 428
rect 6638 416 6644 428
rect 6696 416 6702 468
rect 11256 456 11284 496
rect 12618 484 12624 496
rect 12676 484 12682 536
rect 13354 484 13360 536
rect 13412 524 13418 536
rect 16666 524 16672 536
rect 13412 496 16672 524
rect 13412 484 13418 496
rect 16666 484 16672 496
rect 16724 484 16730 536
rect 17402 484 17408 536
rect 17460 524 17466 536
rect 20070 524 20076 536
rect 17460 496 20076 524
rect 17460 484 17466 496
rect 20070 484 20076 496
rect 20128 484 20134 536
rect 29012 524 29040 564
rect 30098 552 30104 604
rect 30156 592 30162 604
rect 32582 592 32588 604
rect 30156 564 32588 592
rect 30156 552 30162 564
rect 32582 552 32588 564
rect 32640 552 32646 604
rect 33594 552 33600 604
rect 33652 592 33658 604
rect 36078 592 36084 604
rect 33652 564 36084 592
rect 33652 552 33658 564
rect 36078 552 36084 564
rect 36136 552 36142 604
rect 37182 552 37188 604
rect 37240 552 37246 604
rect 38626 592 38654 632
rect 40678 620 40684 672
rect 40736 660 40742 672
rect 42794 660 42800 672
rect 40736 632 42800 660
rect 40736 620 40742 632
rect 42794 620 42800 632
rect 42852 620 42858 672
rect 46658 620 46664 672
rect 46716 660 46722 672
rect 48498 660 48504 672
rect 46716 632 48504 660
rect 46716 620 46722 632
rect 48498 620 48504 632
rect 48556 620 48562 672
rect 48958 620 48964 672
rect 49016 660 49022 672
rect 50798 660 50804 672
rect 49016 632 50804 660
rect 49016 620 49022 632
rect 50798 620 50804 632
rect 50856 620 50862 672
rect 53742 620 53748 672
rect 53800 660 53806 672
rect 55398 660 55404 672
rect 53800 632 55404 660
rect 53800 620 53806 632
rect 55398 620 55404 632
rect 55456 620 55462 672
rect 64322 620 64328 672
rect 64380 660 64386 672
rect 65610 660 65616 672
rect 64380 632 65616 660
rect 64380 620 64386 632
rect 65610 620 65616 632
rect 65668 620 65674 672
rect 66714 620 66720 672
rect 66772 660 66778 672
rect 68002 660 68008 672
rect 66772 632 68008 660
rect 66772 620 66778 632
rect 68002 620 68008 632
rect 68060 620 68066 672
rect 69106 620 69112 672
rect 69164 660 69170 672
rect 70578 660 70584 672
rect 69164 632 70584 660
rect 69164 620 69170 632
rect 70578 620 70584 632
rect 70636 620 70642 672
rect 133230 620 133236 672
rect 133288 660 133294 672
rect 134150 660 134156 672
rect 133288 632 134156 660
rect 133288 620 133294 632
rect 134150 620 134156 632
rect 134208 620 134214 672
rect 136174 620 136180 672
rect 136232 660 136238 672
rect 137646 660 137652 672
rect 136232 632 137652 660
rect 136232 620 136238 632
rect 137646 620 137652 632
rect 137704 620 137710 672
rect 138750 620 138756 672
rect 138808 660 138814 672
rect 140038 660 140044 672
rect 138808 632 140044 660
rect 138808 620 138814 632
rect 140038 620 140044 632
rect 140096 620 140102 672
rect 151354 620 151360 672
rect 151412 660 151418 672
rect 153010 660 153016 672
rect 151412 632 153016 660
rect 151412 620 151418 632
rect 153010 620 153016 632
rect 153068 620 153074 672
rect 153654 620 153660 672
rect 153712 660 153718 672
rect 155402 660 155408 672
rect 153712 632 155408 660
rect 153712 620 153718 632
rect 155402 620 155408 632
rect 155460 620 155466 672
rect 162762 620 162768 672
rect 162820 660 162826 672
rect 164878 660 164884 672
rect 162820 632 164884 660
rect 162820 620 162826 632
rect 164878 620 164884 632
rect 164936 620 164942 672
rect 166074 660 166080 672
rect 165908 632 166080 660
rect 40770 592 40776 604
rect 38626 564 40776 592
rect 40770 552 40776 564
rect 40828 552 40834 604
rect 41874 552 41880 604
rect 41932 592 41938 604
rect 43990 592 43996 604
rect 41932 564 43996 592
rect 41932 552 41938 564
rect 43990 552 43996 564
rect 44048 552 44054 604
rect 47854 552 47860 604
rect 47912 592 47918 604
rect 49602 592 49608 604
rect 47912 564 49608 592
rect 47912 552 47918 564
rect 49602 552 49608 564
rect 49660 552 49666 604
rect 50154 552 50160 604
rect 50212 552 50218 604
rect 51350 552 51356 604
rect 51408 592 51414 604
rect 53006 592 53012 604
rect 51408 564 53012 592
rect 51408 552 51414 564
rect 53006 552 53012 564
rect 53064 552 53070 604
rect 54938 552 54944 604
rect 54996 592 55002 604
rect 56410 592 56416 604
rect 54996 564 56416 592
rect 54996 552 55002 564
rect 56410 552 56416 564
rect 56468 552 56474 604
rect 60826 552 60832 604
rect 60884 592 60890 604
rect 62114 592 62120 604
rect 60884 564 62120 592
rect 60884 552 60890 564
rect 62114 552 62120 564
rect 62172 552 62178 604
rect 65518 552 65524 604
rect 65576 592 65582 604
rect 66806 592 66812 604
rect 65576 564 66812 592
rect 65576 552 65582 564
rect 66806 552 66812 564
rect 66864 552 66870 604
rect 70302 552 70308 604
rect 70360 592 70366 604
rect 71222 592 71228 604
rect 70360 564 71228 592
rect 70360 552 70366 564
rect 71222 552 71228 564
rect 71280 552 71286 604
rect 76190 552 76196 604
rect 76248 592 76254 604
rect 76926 592 76932 604
rect 76248 564 76932 592
rect 76248 552 76254 564
rect 76926 552 76932 564
rect 76984 552 76990 604
rect 77386 552 77392 604
rect 77444 592 77450 604
rect 78030 592 78036 604
rect 77444 564 78036 592
rect 77444 552 77450 564
rect 78030 552 78036 564
rect 78088 552 78094 604
rect 78582 552 78588 604
rect 78640 592 78646 604
rect 79134 592 79140 604
rect 78640 564 79140 592
rect 78640 552 78646 564
rect 79134 552 79140 564
rect 79192 552 79198 604
rect 79686 552 79692 604
rect 79744 592 79750 604
rect 80330 592 80336 604
rect 79744 564 80336 592
rect 79744 552 79750 564
rect 80330 552 80336 564
rect 80388 552 80394 604
rect 80882 552 80888 604
rect 80940 592 80946 604
rect 81434 592 81440 604
rect 80940 564 81440 592
rect 80940 552 80946 564
rect 81434 552 81440 564
rect 81492 552 81498 604
rect 82078 552 82084 604
rect 82136 592 82142 604
rect 82722 592 82728 604
rect 82136 564 82728 592
rect 82136 552 82142 564
rect 82722 552 82728 564
rect 82780 552 82786 604
rect 121822 552 121828 604
rect 121880 592 121886 604
rect 122282 592 122288 604
rect 121880 564 122288 592
rect 121880 552 121886 564
rect 122282 552 122288 564
rect 122340 552 122346 604
rect 124122 552 124128 604
rect 124180 592 124186 604
rect 124674 592 124680 604
rect 124180 564 124680 592
rect 124180 552 124186 564
rect 124674 552 124680 564
rect 124732 552 124738 604
rect 125226 552 125232 604
rect 125284 592 125290 604
rect 125870 592 125876 604
rect 125284 564 125876 592
rect 125284 552 125290 564
rect 125870 552 125876 564
rect 125928 552 125934 604
rect 126422 552 126428 604
rect 126480 592 126486 604
rect 126974 592 126980 604
rect 126480 564 126980 592
rect 126480 552 126486 564
rect 126974 552 126980 564
rect 127032 552 127038 604
rect 127526 552 127532 604
rect 127584 592 127590 604
rect 128170 592 128176 604
rect 127584 564 128176 592
rect 127584 552 127590 564
rect 128170 552 128176 564
rect 128228 552 128234 604
rect 128630 552 128636 604
rect 128688 592 128694 604
rect 129366 592 129372 604
rect 128688 564 129372 592
rect 128688 552 128694 564
rect 129366 552 129372 564
rect 129424 552 129430 604
rect 133874 552 133880 604
rect 133932 592 133938 604
rect 135254 592 135260 604
rect 133932 564 135260 592
rect 133932 552 133938 564
rect 135254 552 135260 564
rect 135312 552 135318 604
rect 136450 552 136456 604
rect 136508 552 136514 604
rect 137554 552 137560 604
rect 137612 592 137618 604
rect 138842 592 138848 604
rect 137612 564 138848 592
rect 137612 552 137618 564
rect 138842 552 138848 564
rect 138900 552 138906 604
rect 139946 552 139952 604
rect 140004 592 140010 604
rect 141234 592 141240 604
rect 140004 564 141240 592
rect 140004 552 140010 564
rect 141234 552 141240 564
rect 141292 552 141298 604
rect 144546 552 144552 604
rect 144604 592 144610 604
rect 145926 592 145932 604
rect 144604 564 145932 592
rect 144604 552 144610 564
rect 145926 552 145932 564
rect 145984 552 145990 604
rect 146846 552 146852 604
rect 146904 592 146910 604
rect 148318 592 148324 604
rect 146904 564 148324 592
rect 146904 552 146910 564
rect 148318 552 148324 564
rect 148376 552 148382 604
rect 152550 552 152556 604
rect 152608 592 152614 604
rect 154206 592 154212 604
rect 152608 564 154212 592
rect 152608 552 152614 564
rect 154206 552 154212 564
rect 154264 552 154270 604
rect 154758 552 154764 604
rect 154816 592 154822 604
rect 156598 592 156604 604
rect 154816 564 156604 592
rect 154816 552 154822 564
rect 156598 552 156604 564
rect 156656 552 156662 604
rect 157058 552 157064 604
rect 157116 592 157122 604
rect 158898 592 158904 604
rect 157116 564 158904 592
rect 157116 552 157122 564
rect 158898 552 158904 564
rect 158956 552 158962 604
rect 161566 552 161572 604
rect 161624 592 161630 604
rect 163682 592 163688 604
rect 161624 564 163688 592
rect 161624 552 161630 564
rect 163682 552 163688 564
rect 163740 552 163746 604
rect 31662 524 31668 536
rect 29012 496 31668 524
rect 31662 484 31668 496
rect 31720 484 31726 536
rect 33226 484 33232 536
rect 33284 524 33290 536
rect 34974 524 34980 536
rect 33284 496 34980 524
rect 33284 484 33290 496
rect 34974 484 34980 496
rect 35032 484 35038 536
rect 14458 456 14464 468
rect 11256 428 14464 456
rect 14458 416 14464 428
rect 14516 416 14522 468
rect 14550 416 14556 468
rect 14608 456 14614 468
rect 17862 456 17868 468
rect 14608 428 17868 456
rect 14608 416 14614 428
rect 17862 416 17868 428
rect 17920 416 17926 468
rect 24394 416 24400 468
rect 24452 456 24458 468
rect 26878 456 26884 468
rect 24452 428 26884 456
rect 24452 416 24458 428
rect 26878 416 26884 428
rect 26936 416 26942 468
rect 37200 456 37228 552
rect 50172 524 50200 552
rect 51902 524 51908 536
rect 50172 496 51908 524
rect 51902 484 51908 496
rect 51960 484 51966 536
rect 63494 484 63500 536
rect 63552 524 63558 536
rect 64506 524 64512 536
rect 63552 496 64512 524
rect 63552 484 63558 496
rect 64506 484 64512 496
rect 64564 484 64570 536
rect 67726 484 67732 536
rect 67784 524 67790 536
rect 69382 524 69388 536
rect 67784 496 69388 524
rect 67784 484 67790 496
rect 69382 484 69388 496
rect 69440 484 69446 536
rect 134978 484 134984 536
rect 135036 524 135042 536
rect 136468 524 136496 552
rect 135036 496 136496 524
rect 135036 484 135042 496
rect 141050 484 141056 536
rect 141108 524 141114 536
rect 142062 524 142068 536
rect 141108 496 142068 524
rect 141108 484 141114 496
rect 142062 484 142068 496
rect 142120 484 142126 536
rect 158162 484 158168 536
rect 158220 524 158226 536
rect 159726 524 159732 536
rect 158220 496 159732 524
rect 158220 484 158226 496
rect 159726 484 159732 496
rect 159784 484 159790 536
rect 39850 456 39856 468
rect 37200 428 39856 456
rect 39850 416 39856 428
rect 39908 416 39914 468
rect 163406 416 163412 468
rect 163464 456 163470 468
rect 165908 456 165936 632
rect 166074 620 166080 632
rect 166132 620 166138 672
rect 167086 620 167092 672
rect 167144 660 167150 672
rect 169570 660 169576 672
rect 167144 632 169576 660
rect 167144 620 167150 632
rect 169570 620 169576 632
rect 169628 620 169634 672
rect 180886 620 180892 672
rect 180944 660 180950 672
rect 183738 660 183744 672
rect 180944 632 183744 660
rect 180944 620 180950 632
rect 183738 620 183744 632
rect 183796 620 183802 672
rect 186130 660 186136 672
rect 184216 632 186136 660
rect 165982 552 165988 604
rect 166040 592 166046 604
rect 168374 592 168380 604
rect 166040 564 168380 592
rect 166040 552 166046 564
rect 168374 552 168380 564
rect 168432 552 168438 604
rect 170674 552 170680 604
rect 170732 592 170738 604
rect 173158 592 173164 604
rect 170732 564 173164 592
rect 170732 552 170738 564
rect 173158 552 173164 564
rect 173216 552 173222 604
rect 179782 552 179788 604
rect 179840 592 179846 604
rect 182542 592 182548 604
rect 179840 564 182548 592
rect 179840 552 179846 564
rect 182542 552 182548 564
rect 182600 552 182606 604
rect 183186 552 183192 604
rect 183244 592 183250 604
rect 184216 592 184244 632
rect 186130 620 186136 632
rect 186188 620 186194 672
rect 191098 620 191104 672
rect 191156 660 191162 672
rect 194410 660 194416 672
rect 191156 632 194416 660
rect 191156 620 191162 632
rect 194410 620 194416 632
rect 194468 620 194474 672
rect 211614 620 211620 672
rect 211672 660 211678 672
rect 215662 660 215668 672
rect 211672 632 215668 660
rect 211672 620 211678 632
rect 215662 620 215668 632
rect 215720 620 215726 672
rect 220170 620 220176 672
rect 220228 660 220234 672
rect 225322 660 225328 672
rect 220228 632 225328 660
rect 220228 620 220234 632
rect 225322 620 225328 632
rect 225380 620 225386 672
rect 226150 620 226156 672
rect 226208 660 226214 672
rect 231026 660 231032 672
rect 226208 632 231032 660
rect 226208 620 226214 632
rect 231026 620 231032 632
rect 231084 620 231090 672
rect 234614 660 234620 672
rect 231780 632 234620 660
rect 183244 564 184244 592
rect 183244 552 183250 564
rect 189994 552 190000 604
rect 190052 592 190058 604
rect 193214 592 193220 604
rect 190052 564 193220 592
rect 190052 552 190058 564
rect 193214 552 193220 564
rect 193272 552 193278 604
rect 195606 552 195612 604
rect 195664 552 195670 604
rect 196802 592 196808 604
rect 196763 564 196808 592
rect 196802 552 196808 564
rect 196860 552 196866 604
rect 197906 552 197912 604
rect 197964 552 197970 604
rect 205726 552 205732 604
rect 205784 592 205790 604
rect 209774 592 209780 604
rect 205784 564 209780 592
rect 205784 552 205790 564
rect 209774 552 209780 564
rect 209832 552 209838 604
rect 210418 552 210424 604
rect 210476 592 210482 604
rect 212077 595 212135 601
rect 212077 592 212089 595
rect 210476 564 212089 592
rect 210476 552 210482 564
rect 212077 561 212089 564
rect 212123 561 212135 595
rect 212077 555 212135 561
rect 212166 552 212172 604
rect 212224 552 212230 604
rect 214466 592 214472 604
rect 214427 564 214472 592
rect 214466 552 214472 564
rect 214524 552 214530 604
rect 219986 552 219992 604
rect 220044 592 220050 604
rect 220446 592 220452 604
rect 220044 564 220452 592
rect 220044 552 220050 564
rect 220446 552 220452 564
rect 220504 552 220510 604
rect 223942 552 223948 604
rect 224000 552 224006 604
rect 225046 552 225052 604
rect 225104 592 225110 604
rect 229830 592 229836 604
rect 225104 564 227714 592
rect 225104 552 225110 564
rect 186590 484 186596 536
rect 186648 524 186654 536
rect 189902 524 189908 536
rect 186648 496 189908 524
rect 186648 484 186654 496
rect 189902 484 189908 496
rect 189960 484 189966 536
rect 192294 484 192300 536
rect 192352 524 192358 536
rect 195624 524 195652 552
rect 192352 496 195652 524
rect 192352 484 192358 496
rect 163464 428 165936 456
rect 163464 416 163470 428
rect 187694 416 187700 468
rect 187752 456 187758 468
rect 191006 456 191012 468
rect 187752 428 191012 456
rect 187752 416 187758 428
rect 191006 416 191012 428
rect 191064 416 191070 468
rect 194042 416 194048 468
rect 194100 456 194106 468
rect 197924 456 197952 552
rect 208394 484 208400 536
rect 208452 524 208458 536
rect 212184 524 212212 552
rect 208452 496 212212 524
rect 208452 484 208458 496
rect 212718 484 212724 536
rect 212776 524 212782 536
rect 216582 524 216588 536
rect 212776 496 216588 524
rect 212776 484 212782 496
rect 216582 484 216588 496
rect 216640 484 216646 536
rect 219526 484 219532 536
rect 219584 524 219590 536
rect 223960 524 223988 552
rect 219584 496 223988 524
rect 219584 484 219590 496
rect 227346 484 227352 536
rect 227404 484 227410 536
rect 227686 524 227714 564
rect 229066 564 229836 592
rect 229066 524 229094 564
rect 229830 552 229836 564
rect 229888 552 229894 604
rect 227686 496 229094 524
rect 229646 484 229652 536
rect 229704 524 229710 536
rect 231780 524 231808 632
rect 234614 620 234620 632
rect 234672 620 234678 672
rect 235442 620 235448 672
rect 235500 660 235506 672
rect 237346 660 237374 700
rect 240505 697 240517 700
rect 240551 697 240563 731
rect 252373 731 252431 737
rect 252373 728 252385 731
rect 240505 691 240563 697
rect 246776 700 252385 728
rect 246776 672 246804 700
rect 252373 697 252385 700
rect 252419 697 252431 731
rect 314626 728 314654 768
rect 340846 768 342361 796
rect 340846 728 340874 768
rect 342349 765 342361 768
rect 342395 765 342407 799
rect 351273 799 351331 805
rect 351273 796 351285 799
rect 342349 759 342407 765
rect 343606 768 351285 796
rect 252373 691 252431 697
rect 279252 700 285674 728
rect 279252 672 279280 700
rect 235500 632 237374 660
rect 235500 620 235506 632
rect 237742 620 237748 672
rect 237800 660 237806 672
rect 242894 660 242900 672
rect 237800 632 242900 660
rect 237800 620 237806 632
rect 242894 620 242900 632
rect 242952 620 242958 672
rect 246758 620 246764 672
rect 246816 620 246822 672
rect 247954 620 247960 672
rect 248012 660 248018 672
rect 253474 660 253480 672
rect 248012 632 253480 660
rect 248012 620 248018 632
rect 253474 620 253480 632
rect 253532 620 253538 672
rect 257246 620 257252 672
rect 257304 660 257310 672
rect 258258 660 258264 672
rect 257304 632 258264 660
rect 257304 620 257310 632
rect 258258 620 258264 632
rect 258316 620 258322 672
rect 260650 660 260656 672
rect 259288 632 260656 660
rect 231854 552 231860 604
rect 231912 592 231918 604
rect 237006 592 237012 604
rect 231912 564 237012 592
rect 231912 552 231918 564
rect 237006 552 237012 564
rect 237064 552 237070 604
rect 238110 552 238116 604
rect 238168 552 238174 604
rect 239306 592 239312 604
rect 238404 564 239312 592
rect 229704 496 231808 524
rect 229704 484 229710 496
rect 233142 484 233148 536
rect 233200 524 233206 536
rect 238128 524 238156 552
rect 233200 496 238156 524
rect 233200 484 233206 496
rect 194100 428 197952 456
rect 212077 459 212135 465
rect 194100 416 194106 428
rect 212077 425 212089 459
rect 212123 456 212135 459
rect 214469 459 214527 465
rect 214469 456 214481 459
rect 212123 428 214481 456
rect 212123 425 212135 428
rect 212077 419 212135 425
rect 214469 425 214481 428
rect 214515 425 214527 459
rect 214469 419 214527 425
rect 218422 416 218428 468
rect 218480 456 218486 468
rect 222930 456 222936 468
rect 218480 428 222936 456
rect 218480 416 218486 428
rect 222930 416 222936 428
rect 222988 416 222994 468
rect 227364 456 227392 484
rect 224926 428 227392 456
rect 39298 348 39304 400
rect 39356 388 39362 400
rect 42150 388 42156 400
rect 39356 360 42156 388
rect 39356 348 39362 360
rect 42150 348 42156 360
rect 42208 348 42214 400
rect 42886 348 42892 400
rect 42944 388 42950 400
rect 45094 388 45100 400
rect 42944 360 45100 388
rect 42944 348 42950 360
rect 45094 348 45100 360
rect 45152 348 45158 400
rect 71314 348 71320 400
rect 71372 388 71378 400
rect 72326 388 72332 400
rect 71372 360 72332 388
rect 71372 348 71378 360
rect 72326 348 72332 360
rect 72384 348 72390 400
rect 72418 348 72424 400
rect 72476 388 72482 400
rect 73522 388 73528 400
rect 72476 360 73528 388
rect 72476 348 72482 360
rect 73522 348 73528 360
rect 73580 348 73586 400
rect 73614 348 73620 400
rect 73672 388 73678 400
rect 74626 388 74632 400
rect 73672 360 74632 388
rect 73672 348 73678 360
rect 74626 348 74632 360
rect 74684 348 74690 400
rect 130930 348 130936 400
rect 130988 388 130994 400
rect 131942 388 131948 400
rect 130988 360 131948 388
rect 130988 348 130994 360
rect 131942 348 131948 360
rect 132000 348 132006 400
rect 132034 348 132040 400
rect 132092 388 132098 400
rect 133138 388 133144 400
rect 132092 360 133144 388
rect 132092 348 132098 360
rect 133138 348 133144 360
rect 133196 348 133202 400
rect 160462 348 160468 400
rect 160520 388 160526 400
rect 162670 388 162676 400
rect 160520 360 162676 388
rect 160520 348 160526 360
rect 162670 348 162676 360
rect 162728 348 162734 400
rect 192938 348 192944 400
rect 192996 388 193002 400
rect 196805 391 196863 397
rect 196805 388 196817 391
rect 192996 360 196817 388
rect 192996 348 193002 360
rect 196805 357 196817 360
rect 196851 357 196863 391
rect 196805 351 196863 357
rect 217226 348 217232 400
rect 217284 388 217290 400
rect 221734 388 221740 400
rect 217284 360 221740 388
rect 217284 348 217290 360
rect 221734 348 221740 360
rect 221792 348 221798 400
rect 222470 348 222476 400
rect 222528 388 222534 400
rect 224926 388 224954 428
rect 234338 416 234344 468
rect 234396 456 234402 468
rect 238404 456 238432 564
rect 239306 552 239312 564
rect 239364 552 239370 604
rect 240502 592 240508 604
rect 240463 564 240508 592
rect 240502 552 240508 564
rect 240560 552 240566 604
rect 241146 552 241152 604
rect 241204 592 241210 604
rect 246022 592 246028 604
rect 241204 564 246028 592
rect 241204 552 241210 564
rect 246022 552 246028 564
rect 246080 552 246086 604
rect 249978 552 249984 604
rect 250036 552 250042 604
rect 251174 552 251180 604
rect 251232 552 251238 604
rect 252370 592 252376 604
rect 252331 564 252376 592
rect 252370 552 252376 564
rect 252428 552 252434 604
rect 253382 552 253388 604
rect 253440 552 253446 604
rect 254578 552 254584 604
rect 254636 592 254642 604
rect 259288 592 259316 632
rect 260650 620 260656 632
rect 260708 620 260714 672
rect 262674 620 262680 672
rect 262732 660 262738 672
rect 268838 660 268844 672
rect 262732 632 268844 660
rect 262732 620 262738 632
rect 268838 620 268844 632
rect 268896 620 268902 672
rect 269482 620 269488 672
rect 269540 660 269546 672
rect 276198 660 276204 672
rect 269540 632 276204 660
rect 269540 620 269546 632
rect 276198 620 276204 632
rect 276256 620 276262 672
rect 279234 620 279240 672
rect 279292 620 279298 672
rect 279510 660 279516 672
rect 279471 632 279516 660
rect 279510 620 279516 632
rect 279568 620 279574 672
rect 284294 660 284300 672
rect 280126 632 284300 660
rect 259454 592 259460 604
rect 254636 564 259316 592
rect 259380 564 259460 592
rect 254636 552 254642 564
rect 238846 484 238852 536
rect 238904 524 238910 536
rect 243906 524 243912 536
rect 238904 496 243912 524
rect 238904 484 238910 496
rect 243906 484 243912 496
rect 243964 484 243970 536
rect 248966 524 248972 536
rect 244246 496 248972 524
rect 234396 428 238432 456
rect 234396 416 234402 428
rect 243354 416 243360 468
rect 243412 456 243418 468
rect 244246 456 244274 496
rect 248966 484 248972 496
rect 249024 484 249030 536
rect 243412 428 244274 456
rect 243412 416 243418 428
rect 244550 416 244556 468
rect 244608 456 244614 468
rect 249996 456 250024 552
rect 244608 428 250024 456
rect 244608 416 244614 428
rect 222528 360 224954 388
rect 222528 348 222534 360
rect 242250 348 242256 400
rect 242308 388 242314 400
rect 247310 388 247316 400
rect 242308 360 247316 388
rect 242308 348 242314 360
rect 247310 348 247316 360
rect 247368 348 247374 400
rect 245654 280 245660 332
rect 245712 320 245718 332
rect 251192 320 251220 552
rect 253400 524 253428 552
rect 259380 524 259408 564
rect 259454 552 259460 564
rect 259512 552 259518 604
rect 260466 552 260472 604
rect 260524 592 260530 604
rect 266538 592 266544 604
rect 260524 564 266544 592
rect 260524 552 260530 564
rect 266538 552 266544 564
rect 266596 552 266602 604
rect 267734 552 267740 604
rect 267792 552 267798 604
rect 270034 592 270040 604
rect 269995 564 270040 592
rect 270034 552 270040 564
rect 270092 552 270098 604
rect 271782 552 271788 604
rect 271840 592 271846 604
rect 271840 564 276014 592
rect 271840 552 271846 564
rect 253400 496 259408 524
rect 261570 484 261576 536
rect 261628 524 261634 536
rect 267752 524 267780 552
rect 261628 496 267780 524
rect 261628 484 261634 496
rect 268378 484 268384 536
rect 268436 524 268442 536
rect 274542 524 274548 536
rect 268436 496 274548 524
rect 268436 484 268442 496
rect 274542 484 274548 496
rect 274600 484 274606 536
rect 275986 524 276014 564
rect 277486 552 277492 604
rect 277544 592 277550 604
rect 280126 592 280154 632
rect 284294 620 284300 632
rect 284352 620 284358 672
rect 285646 660 285674 700
rect 304966 700 312676 728
rect 314626 700 315896 728
rect 286594 660 286600 672
rect 285646 632 286600 660
rect 286594 620 286600 632
rect 286652 620 286658 672
rect 291102 620 291108 672
rect 291160 660 291166 672
rect 298462 660 298468 672
rect 291160 632 298468 660
rect 291160 620 291166 632
rect 298462 620 298468 632
rect 298520 620 298526 672
rect 304718 620 304724 672
rect 304776 660 304782 672
rect 304966 660 304994 700
rect 312648 672 312676 700
rect 307662 660 307668 672
rect 304776 632 304994 660
rect 307623 632 307668 660
rect 304776 620 304782 632
rect 307662 620 307668 632
rect 307720 620 307726 672
rect 309962 620 309968 672
rect 310020 660 310026 672
rect 310020 632 312354 660
rect 310020 620 310026 632
rect 280706 592 280712 604
rect 277544 564 280154 592
rect 280667 564 280712 592
rect 277544 552 277550 564
rect 280706 552 280712 564
rect 280764 552 280770 604
rect 283098 592 283104 604
rect 283059 564 283104 592
rect 283098 552 283104 564
rect 283156 552 283162 604
rect 285398 552 285404 604
rect 285456 552 285462 604
rect 288802 552 288808 604
rect 288860 592 288866 604
rect 296070 592 296076 604
rect 288860 564 296076 592
rect 288860 552 288866 564
rect 296070 552 296076 564
rect 296128 552 296134 604
rect 297266 592 297272 604
rect 296364 564 297272 592
rect 278498 524 278504 536
rect 275986 496 278504 524
rect 278498 484 278504 496
rect 278556 484 278562 536
rect 278590 484 278596 536
rect 278648 524 278654 536
rect 285416 524 285444 552
rect 278648 496 285444 524
rect 278648 484 278654 496
rect 286410 484 286416 536
rect 286468 524 286474 536
rect 293310 524 293316 536
rect 286468 496 293316 524
rect 286468 484 286474 496
rect 293310 484 293316 496
rect 293368 484 293374 536
rect 256878 456 256884 468
rect 245712 292 251220 320
rect 251836 428 256884 456
rect 245712 280 245718 292
rect 227346 212 227352 264
rect 227404 252 227410 264
rect 232038 252 232044 264
rect 227404 224 232044 252
rect 227404 212 227410 224
rect 232038 212 232044 224
rect 232096 212 232102 264
rect 233234 212 233240 264
rect 233292 212 233298 264
rect 250898 212 250904 264
rect 250956 252 250962 264
rect 251836 252 251864 428
rect 256878 416 256884 428
rect 256936 416 256942 468
rect 257982 416 257988 468
rect 258040 456 258046 468
rect 258040 416 258074 456
rect 259270 416 259276 468
rect 259328 456 259334 468
rect 264974 456 264980 468
rect 259328 428 264980 456
rect 259328 416 259334 428
rect 264974 416 264980 428
rect 265032 416 265038 468
rect 266078 416 266084 468
rect 266136 456 266142 468
rect 272150 456 272156 468
rect 266136 428 272156 456
rect 266136 416 266142 428
rect 272150 416 272156 428
rect 272208 416 272214 468
rect 280430 416 280436 468
rect 280488 456 280494 468
rect 287514 456 287520 468
rect 280488 428 287520 456
rect 280488 416 280494 428
rect 287514 416 287520 428
rect 287572 416 287578 468
rect 289814 416 289820 468
rect 289872 456 289878 468
rect 296364 456 296392 564
rect 297266 552 297272 564
rect 297324 552 297330 604
rect 300210 552 300216 604
rect 300268 592 300274 604
rect 300268 564 304304 592
rect 300268 552 300274 564
rect 296806 484 296812 536
rect 296864 524 296870 536
rect 303982 524 303988 536
rect 296864 496 303988 524
rect 296864 484 296870 496
rect 303982 484 303988 496
rect 304040 484 304046 536
rect 304276 524 304304 564
rect 307938 552 307944 604
rect 307996 552 308002 604
rect 309042 552 309048 604
rect 309100 552 309106 604
rect 310238 552 310244 604
rect 310296 552 310302 604
rect 310333 595 310391 601
rect 310333 561 310345 595
rect 310379 592 310391 595
rect 311434 592 311440 604
rect 310379 564 311440 592
rect 310379 561 310391 564
rect 310333 555 310391 561
rect 311434 552 311440 564
rect 311492 552 311498 604
rect 307956 524 307984 552
rect 304276 496 307984 524
rect 289872 428 296392 456
rect 289872 416 289878 428
rect 301314 416 301320 468
rect 301372 456 301378 468
rect 309060 456 309088 552
rect 301372 428 309088 456
rect 301372 416 301378 428
rect 258046 388 258074 416
rect 263134 388 263140 400
rect 258046 360 263140 388
rect 263134 348 263140 360
rect 263192 348 263198 400
rect 270678 348 270684 400
rect 270736 388 270742 400
rect 276750 388 276756 400
rect 270736 360 276756 388
rect 270736 348 270742 360
rect 276750 348 276756 360
rect 276808 348 276814 400
rect 281534 348 281540 400
rect 281592 388 281598 400
rect 287054 388 287060 400
rect 281592 360 287060 388
rect 281592 348 281598 360
rect 287054 348 287060 360
rect 287112 348 287118 400
rect 287606 348 287612 400
rect 287664 388 287670 400
rect 293862 388 293868 400
rect 287664 360 293868 388
rect 287664 348 287670 360
rect 293862 348 293868 360
rect 293920 348 293926 400
rect 294506 348 294512 400
rect 294564 388 294570 400
rect 301774 388 301780 400
rect 294564 360 301780 388
rect 294564 348 294570 360
rect 301774 348 301780 360
rect 301832 348 301838 400
rect 306926 388 306932 400
rect 302344 360 306932 388
rect 252002 280 252008 332
rect 252060 320 252066 332
rect 257246 320 257252 332
rect 252060 292 257252 320
rect 252060 280 252066 292
rect 257246 280 257252 292
rect 257304 280 257310 332
rect 275830 280 275836 332
rect 275888 320 275894 332
rect 283101 323 283159 329
rect 283101 320 283113 323
rect 275888 292 283113 320
rect 275888 280 275894 292
rect 283101 289 283113 292
rect 283147 289 283159 323
rect 283101 283 283159 289
rect 284110 280 284116 332
rect 284168 320 284174 332
rect 291194 320 291200 332
rect 284168 292 291200 320
rect 284168 280 284174 292
rect 291194 280 291200 292
rect 291252 280 291258 332
rect 299014 280 299020 332
rect 299072 320 299078 332
rect 302344 320 302372 360
rect 306926 348 306932 360
rect 306984 348 306990 400
rect 299072 292 302372 320
rect 299072 280 299078 292
rect 302418 280 302424 332
rect 302476 320 302482 332
rect 310256 320 310284 552
rect 312326 456 312354 632
rect 312630 620 312636 672
rect 312688 620 312694 672
rect 315868 592 315896 700
rect 318720 700 324268 728
rect 315942 620 315948 672
rect 316000 660 316006 672
rect 318720 660 318748 700
rect 319714 660 319720 672
rect 316000 632 318748 660
rect 319675 632 319720 660
rect 316000 620 316006 632
rect 319714 620 319720 632
rect 319772 620 319778 672
rect 320910 660 320916 672
rect 320560 632 320916 660
rect 316218 592 316224 604
rect 315868 564 316224 592
rect 316218 552 316224 564
rect 316276 552 316282 604
rect 320560 592 320588 632
rect 320910 620 320916 632
rect 320968 620 320974 672
rect 321005 663 321063 669
rect 321005 629 321017 663
rect 321051 660 321063 663
rect 323302 660 323308 672
rect 321051 632 323308 660
rect 321051 629 321063 632
rect 321005 623 321063 629
rect 323302 620 323308 632
rect 323360 620 323366 672
rect 324240 660 324268 700
rect 335372 700 340874 728
rect 341797 731 341855 737
rect 335372 672 335400 700
rect 341797 697 341809 731
rect 341843 728 341855 731
rect 343606 728 343634 768
rect 351273 765 351285 768
rect 351319 765 351331 799
rect 351273 759 351331 765
rect 341843 700 343634 728
rect 341843 697 341855 700
rect 341797 691 341855 697
rect 369412 672 369440 836
rect 388257 833 388269 836
rect 388303 833 388315 867
rect 388257 827 388315 833
rect 389913 867 389971 873
rect 389913 833 389925 867
rect 389959 864 389971 867
rect 428461 867 428519 873
rect 428461 864 428473 867
rect 389959 836 401364 864
rect 389959 833 389971 836
rect 389913 827 389971 833
rect 372893 799 372951 805
rect 372893 796 372905 799
rect 369826 768 372905 796
rect 324406 660 324412 672
rect 324240 632 324412 660
rect 324406 620 324412 632
rect 324464 620 324470 672
rect 329190 660 329196 672
rect 325528 632 329196 660
rect 317064 564 320588 592
rect 312446 484 312452 536
rect 312504 524 312510 536
rect 317064 524 317092 564
rect 320634 552 320640 604
rect 320692 592 320698 604
rect 325528 592 325556 632
rect 329190 620 329196 632
rect 329248 620 329254 672
rect 335354 620 335360 672
rect 335412 620 335418 672
rect 335725 663 335783 669
rect 335725 629 335737 663
rect 335771 660 335783 663
rect 337565 663 337623 669
rect 335771 632 337516 660
rect 335771 629 335783 632
rect 335725 623 335783 629
rect 337488 604 337516 632
rect 337565 629 337577 663
rect 337611 660 337623 663
rect 342349 663 342407 669
rect 337611 632 342300 660
rect 337611 629 337623 632
rect 337565 623 337623 629
rect 320692 564 325556 592
rect 320692 552 320698 564
rect 325602 552 325608 604
rect 325660 552 325666 604
rect 327994 552 328000 604
rect 328052 552 328058 604
rect 328457 595 328515 601
rect 328457 561 328469 595
rect 328503 592 328515 595
rect 332686 592 332692 604
rect 328503 564 332692 592
rect 328503 561 328515 564
rect 328457 555 328515 561
rect 332686 552 332692 564
rect 332744 552 332750 604
rect 334250 552 334256 604
rect 334308 592 334314 604
rect 337381 595 337439 601
rect 337381 592 337393 595
rect 334308 564 337393 592
rect 334308 552 334314 564
rect 337381 561 337393 564
rect 337427 561 337439 595
rect 337381 555 337439 561
rect 337470 552 337476 604
rect 337528 552 337534 604
rect 338666 592 338672 604
rect 338627 564 338672 592
rect 338666 552 338672 564
rect 338724 552 338730 604
rect 339862 552 339868 604
rect 339920 552 339926 604
rect 340966 552 340972 604
rect 341024 552 341030 604
rect 341794 592 341800 604
rect 341755 564 341800 592
rect 341794 552 341800 564
rect 341852 552 341858 604
rect 342162 592 342168 604
rect 342123 564 342168 592
rect 342162 552 342168 564
rect 342220 552 342226 604
rect 342272 592 342300 632
rect 342349 629 342361 663
rect 342395 660 342407 663
rect 344554 660 344560 672
rect 342395 632 344560 660
rect 342395 629 342407 632
rect 342349 623 342407 629
rect 344554 620 344560 632
rect 344612 620 344618 672
rect 347682 620 347688 672
rect 347740 660 347746 672
rect 357526 660 357532 672
rect 347740 632 357532 660
rect 347740 620 347746 632
rect 357526 620 357532 632
rect 357584 620 357590 672
rect 367002 660 367008 672
rect 357820 632 367008 660
rect 343358 592 343364 604
rect 342272 564 343364 592
rect 343358 552 343364 564
rect 343416 552 343422 604
rect 343450 552 343456 604
rect 343508 592 343514 604
rect 345750 592 345756 604
rect 343508 564 345756 592
rect 343508 552 343514 564
rect 345750 552 345756 564
rect 345808 552 345814 604
rect 347593 595 347651 601
rect 347593 561 347605 595
rect 347639 592 347651 595
rect 352834 592 352840 604
rect 347639 564 352840 592
rect 347639 561 347651 564
rect 347593 555 347651 561
rect 352834 552 352840 564
rect 352892 552 352898 604
rect 354030 592 354036 604
rect 353220 564 354036 592
rect 312504 496 317092 524
rect 312504 484 312510 496
rect 317138 484 317144 536
rect 317196 524 317202 536
rect 325620 524 325648 552
rect 317196 496 325648 524
rect 317196 484 317202 496
rect 318150 456 318156 468
rect 312326 428 318156 456
rect 318150 416 318156 428
rect 318208 416 318214 468
rect 319530 416 319536 468
rect 319588 456 319594 468
rect 328012 456 328040 552
rect 330846 484 330852 536
rect 330904 524 330910 536
rect 339880 524 339908 552
rect 330904 496 339908 524
rect 330904 484 330910 496
rect 319588 428 328040 456
rect 319588 416 319594 428
rect 331950 416 331956 468
rect 332008 456 332014 468
rect 340984 456 341012 552
rect 347682 484 347688 536
rect 347740 524 347746 536
rect 353220 524 353248 564
rect 354030 552 354036 564
rect 354088 552 354094 604
rect 356330 592 356336 604
rect 356291 564 356336 592
rect 356330 552 356336 564
rect 356388 552 356394 604
rect 356974 552 356980 604
rect 357032 592 357038 604
rect 357820 592 357848 632
rect 367002 620 367008 632
rect 367060 620 367066 672
rect 368198 660 368204 672
rect 368159 632 368204 660
rect 368198 620 368204 632
rect 368256 620 368262 672
rect 369394 620 369400 672
rect 369452 620 369458 672
rect 359274 592 359280 604
rect 357032 564 357848 592
rect 359235 564 359280 592
rect 357032 552 357038 564
rect 359274 552 359280 564
rect 359332 552 359338 604
rect 362678 552 362684 604
rect 362736 592 362742 604
rect 369826 592 369854 768
rect 372893 765 372905 768
rect 372939 765 372951 799
rect 372893 759 372951 765
rect 373169 799 373227 805
rect 373169 765 373181 799
rect 373215 796 373227 799
rect 393225 799 393283 805
rect 393225 796 393237 799
rect 373215 768 382274 796
rect 373215 765 373227 768
rect 373169 759 373227 765
rect 372586 700 375420 728
rect 370406 620 370412 672
rect 370464 660 370470 672
rect 372586 660 372614 700
rect 372890 660 372896 672
rect 370464 632 372614 660
rect 372851 632 372896 660
rect 370464 620 370470 632
rect 372890 620 372896 632
rect 372948 620 372954 672
rect 375392 660 375420 700
rect 379486 700 381216 728
rect 379486 660 379514 700
rect 381188 672 381216 700
rect 375392 632 379514 660
rect 381170 620 381176 672
rect 381228 620 381234 672
rect 382246 660 382274 768
rect 382798 768 393237 796
rect 382366 660 382372 672
rect 382246 632 382372 660
rect 382366 620 382372 632
rect 382424 620 382430 672
rect 362736 564 369854 592
rect 362736 552 362742 564
rect 370682 552 370688 604
rect 370740 552 370746 604
rect 371602 552 371608 604
rect 371660 592 371666 604
rect 373169 595 373227 601
rect 373169 592 373181 595
rect 371660 564 373181 592
rect 371660 552 371666 564
rect 373169 561 373181 564
rect 373215 561 373227 595
rect 373169 555 373227 561
rect 381998 552 382004 604
rect 382056 592 382062 604
rect 382798 592 382826 768
rect 393225 765 393237 768
rect 393271 765 393283 799
rect 393225 759 393283 765
rect 395525 731 395583 737
rect 395525 728 395537 731
rect 384224 700 395537 728
rect 384224 672 384252 700
rect 395525 697 395537 700
rect 395571 697 395583 731
rect 395525 691 395583 697
rect 401336 672 401364 836
rect 405292 836 414336 864
rect 384206 620 384212 672
rect 384264 620 384270 672
rect 386506 660 386512 672
rect 386467 632 386512 660
rect 386506 620 386512 632
rect 386564 620 386570 672
rect 400122 660 400128 672
rect 387766 632 396580 660
rect 400083 632 400128 660
rect 382056 564 382826 592
rect 382056 552 382062 564
rect 383562 552 383568 604
rect 383620 552 383626 604
rect 385402 552 385408 604
rect 385460 592 385466 604
rect 387766 592 387794 632
rect 396552 604 396580 632
rect 400122 620 400128 632
rect 400180 620 400186 672
rect 401318 620 401324 672
rect 401376 620 401382 672
rect 402422 620 402428 672
rect 402480 660 402486 672
rect 405292 660 405320 836
rect 414308 672 414336 836
rect 416746 836 428473 864
rect 405642 660 405648 672
rect 402480 632 405320 660
rect 405603 632 405648 660
rect 402480 620 402486 632
rect 405642 620 405648 632
rect 405700 620 405706 672
rect 407025 663 407083 669
rect 407025 629 407037 663
rect 407071 660 407083 663
rect 407206 660 407212 672
rect 407071 632 407212 660
rect 407071 629 407083 632
rect 407025 623 407083 629
rect 407206 620 407212 632
rect 407264 620 407270 672
rect 408310 660 408316 672
rect 408271 632 408316 660
rect 408310 620 408316 632
rect 408368 620 408374 672
rect 410794 660 410800 672
rect 409064 632 410800 660
rect 388254 592 388260 604
rect 385460 564 387794 592
rect 388215 564 388260 592
rect 385460 552 385466 564
rect 388254 552 388260 564
rect 388312 552 388318 604
rect 389450 592 389456 604
rect 389411 564 389456 592
rect 389450 552 389456 564
rect 389508 552 389514 604
rect 389910 592 389916 604
rect 389871 564 389916 592
rect 389910 552 389916 564
rect 389968 552 389974 604
rect 391014 552 391020 604
rect 391072 592 391078 604
rect 391072 564 395660 592
rect 391072 552 391078 564
rect 347740 496 353248 524
rect 347740 484 347746 496
rect 354674 484 354680 536
rect 354732 524 354738 536
rect 358265 527 358323 533
rect 358265 524 358277 527
rect 354732 496 358277 524
rect 354732 484 354738 496
rect 358265 493 358277 496
rect 358311 493 358323 527
rect 358265 487 358323 493
rect 358538 484 358544 536
rect 358596 484 358602 536
rect 360378 484 360384 536
rect 360436 524 360442 536
rect 370700 524 370728 552
rect 360436 496 370728 524
rect 360436 484 360442 496
rect 372430 484 372436 536
rect 372488 524 372494 536
rect 383580 524 383608 552
rect 394418 524 394424 536
rect 372488 496 383608 524
rect 387352 496 394424 524
rect 372488 484 372494 496
rect 332008 428 341012 456
rect 332008 416 332014 428
rect 343174 416 343180 468
rect 343232 456 343238 468
rect 347593 459 347651 465
rect 347593 456 347605 459
rect 343232 428 347605 456
rect 343232 416 343238 428
rect 347593 425 347605 428
rect 347639 425 347651 459
rect 347593 419 347651 425
rect 349062 416 349068 468
rect 349120 456 349126 468
rect 358556 456 358584 484
rect 349120 428 358584 456
rect 349120 416 349126 428
rect 363782 416 363788 468
rect 363840 456 363846 468
rect 367741 459 367799 465
rect 363840 428 367692 456
rect 363840 416 363846 428
rect 314746 348 314752 400
rect 314804 388 314810 400
rect 314804 360 318288 388
rect 314804 348 314810 360
rect 302476 292 310284 320
rect 302476 280 302482 292
rect 313642 280 313648 332
rect 313700 320 313706 332
rect 318260 320 318288 360
rect 318334 348 318340 400
rect 318392 388 318398 400
rect 326614 388 326620 400
rect 318392 360 326620 388
rect 318392 348 318398 360
rect 326614 348 326620 360
rect 326672 348 326678 400
rect 327442 348 327448 400
rect 327500 388 327506 400
rect 327500 360 331352 388
rect 327500 348 327506 360
rect 321005 323 321063 329
rect 321005 320 321017 323
rect 313700 292 317552 320
rect 318260 292 321017 320
rect 313700 280 313706 292
rect 250956 224 251864 252
rect 250956 212 250962 224
rect 255682 212 255688 264
rect 255740 252 255746 264
rect 261938 252 261944 264
rect 255740 224 261944 252
rect 255740 212 255746 224
rect 261938 212 261944 224
rect 261996 212 262002 264
rect 263686 212 263692 264
rect 263744 252 263750 264
rect 270037 255 270095 261
rect 270037 252 270049 255
rect 263744 224 270049 252
rect 263744 212 263750 224
rect 270037 221 270049 224
rect 270083 221 270095 255
rect 270037 215 270095 221
rect 272886 212 272892 264
rect 272944 252 272950 264
rect 279513 255 279571 261
rect 279513 252 279525 255
rect 272944 224 279525 252
rect 272944 212 272950 224
rect 279513 221 279525 224
rect 279559 221 279571 255
rect 279513 215 279571 221
rect 297910 212 297916 264
rect 297968 252 297974 264
rect 305730 252 305736 264
rect 297968 224 305736 252
rect 297968 212 297974 224
rect 305730 212 305736 224
rect 305788 212 305794 264
rect 308766 212 308772 264
rect 308824 252 308830 264
rect 316402 252 316408 264
rect 308824 224 316408 252
rect 308824 212 308830 224
rect 316402 212 316408 224
rect 316460 212 316466 264
rect 186958 184 186964 196
rect 184906 156 186964 184
rect 16298 76 16304 128
rect 16356 116 16362 128
rect 18966 116 18972 128
rect 16356 88 18972 116
rect 16356 76 16362 88
rect 18966 76 18972 88
rect 19024 76 19030 128
rect 45738 76 45744 128
rect 45796 116 45802 128
rect 47394 116 47400 128
rect 45796 88 47400 116
rect 45796 76 45802 88
rect 47394 76 47400 88
rect 47452 76 47458 128
rect 129826 76 129832 128
rect 129884 116 129890 128
rect 130286 116 130292 128
rect 129884 88 130292 116
rect 129884 76 129890 88
rect 130286 76 130292 88
rect 130344 76 130350 128
rect 155954 76 155960 128
rect 156012 116 156018 128
rect 157518 116 157524 128
rect 156012 88 157524 116
rect 156012 76 156018 88
rect 157518 76 157524 88
rect 157576 76 157582 128
rect 159358 76 159364 128
rect 159416 116 159422 128
rect 161474 116 161480 128
rect 159416 88 161480 116
rect 159416 76 159422 88
rect 161474 76 161480 88
rect 161532 76 161538 128
rect 184290 76 184296 128
rect 184348 116 184354 128
rect 184906 116 184934 156
rect 186958 144 186964 156
rect 187016 144 187022 196
rect 228542 144 228548 196
rect 228600 184 228606 196
rect 233252 184 233280 212
rect 228600 156 233280 184
rect 228600 144 228606 156
rect 236546 144 236552 196
rect 236604 184 236610 196
rect 241422 184 241428 196
rect 236604 156 241428 184
rect 236604 144 236610 156
rect 241422 144 241428 156
rect 241480 144 241486 196
rect 274082 144 274088 196
rect 274140 184 274146 196
rect 280709 187 280767 193
rect 280709 184 280721 187
rect 274140 156 280721 184
rect 274140 144 274146 156
rect 280709 153 280721 156
rect 280755 153 280767 187
rect 280709 147 280767 153
rect 282914 144 282920 196
rect 282972 184 282978 196
rect 289998 184 290004 196
rect 282972 156 290004 184
rect 282972 144 282978 156
rect 289998 144 290004 156
rect 290056 144 290062 196
rect 292206 144 292212 196
rect 292264 184 292270 196
rect 299382 184 299388 196
rect 292264 156 299388 184
rect 292264 144 292270 156
rect 299382 144 299388 156
rect 299440 144 299446 196
rect 317524 184 317552 292
rect 321005 289 321017 292
rect 321051 289 321063 323
rect 321005 283 321063 289
rect 321554 280 321560 332
rect 321612 320 321618 332
rect 330110 320 330116 332
rect 321612 292 330116 320
rect 321612 280 321618 292
rect 330110 280 330116 292
rect 330168 280 330174 332
rect 331324 320 331352 360
rect 333146 348 333152 400
rect 333204 388 333210 400
rect 338761 391 338819 397
rect 338761 388 338773 391
rect 333204 360 338773 388
rect 333204 348 333210 360
rect 338761 357 338773 360
rect 338807 357 338819 391
rect 338761 351 338819 357
rect 340598 348 340604 400
rect 340656 388 340662 400
rect 350166 388 350172 400
rect 340656 360 350172 388
rect 340656 348 340662 360
rect 350166 348 350172 360
rect 350224 348 350230 400
rect 351270 388 351276 400
rect 351231 360 351276 388
rect 351270 348 351276 360
rect 351328 348 351334 400
rect 352466 348 352472 400
rect 352524 388 352530 400
rect 355781 391 355839 397
rect 355781 388 355793 391
rect 352524 360 355793 388
rect 352524 348 352530 360
rect 355781 357 355793 360
rect 355827 357 355839 391
rect 355781 351 355839 357
rect 355870 348 355876 400
rect 355928 388 355934 400
rect 365990 388 365996 400
rect 355928 360 365996 388
rect 355928 348 355934 360
rect 365990 348 365996 360
rect 366048 348 366054 400
rect 336458 320 336464 332
rect 331324 292 336464 320
rect 336458 280 336464 292
rect 336516 280 336522 332
rect 337194 280 337200 332
rect 337252 320 337258 332
rect 346670 320 346676 332
rect 337252 292 346676 320
rect 337252 280 337258 292
rect 346670 280 346676 292
rect 346728 280 346734 332
rect 356333 323 356391 329
rect 356333 320 356345 323
rect 350506 292 356345 320
rect 328457 255 328515 261
rect 328457 252 328469 255
rect 324286 224 328469 252
rect 321830 184 321836 196
rect 317524 156 321836 184
rect 321830 144 321836 156
rect 321888 144 321894 196
rect 324038 144 324044 196
rect 324096 184 324102 196
rect 324286 184 324314 224
rect 328457 221 328469 224
rect 328503 221 328515 255
rect 328457 215 328515 221
rect 328546 212 328552 264
rect 328604 252 328610 264
rect 335725 255 335783 261
rect 335725 252 335737 255
rect 328604 224 335737 252
rect 328604 212 328610 224
rect 335725 221 335737 224
rect 335771 221 335783 255
rect 335725 215 335783 221
rect 338761 255 338819 261
rect 338761 221 338773 255
rect 338807 252 338819 255
rect 342165 255 342223 261
rect 342165 252 342177 255
rect 338807 224 342177 252
rect 338807 221 338819 224
rect 338761 215 338819 221
rect 342165 221 342177 224
rect 342211 221 342223 255
rect 342165 215 342223 221
rect 346762 212 346768 264
rect 346820 252 346826 264
rect 350506 252 350534 292
rect 356333 289 356345 292
rect 356379 289 356391 323
rect 356333 283 356391 289
rect 358265 323 358323 329
rect 358265 289 358277 323
rect 358311 320 358323 323
rect 364794 320 364800 332
rect 358311 292 364800 320
rect 358311 289 358323 292
rect 358265 283 358323 289
rect 364794 280 364800 292
rect 364852 280 364858 332
rect 367664 320 367692 428
rect 367741 425 367753 459
rect 367787 456 367799 459
rect 367787 428 372614 456
rect 367787 425 367799 428
rect 367741 419 367799 425
rect 372586 388 372614 428
rect 375098 416 375104 468
rect 375156 456 375162 468
rect 379698 456 379704 468
rect 375156 428 379704 456
rect 375156 416 375162 428
rect 379698 416 379704 428
rect 379756 416 379762 468
rect 380069 459 380127 465
rect 380069 425 380081 459
rect 380115 456 380127 459
rect 380115 428 380940 456
rect 380115 425 380127 428
rect 380069 419 380127 425
rect 377398 388 377404 400
rect 372586 360 377404 388
rect 377398 348 377404 360
rect 377456 348 377462 400
rect 378594 348 378600 400
rect 378652 388 378658 400
rect 379885 391 379943 397
rect 379885 388 379897 391
rect 378652 360 379897 388
rect 378652 348 378658 360
rect 379885 357 379897 360
rect 379931 357 379943 391
rect 380912 388 380940 428
rect 383102 416 383108 468
rect 383160 456 383166 468
rect 387352 456 387380 496
rect 394418 484 394424 496
rect 394476 484 394482 536
rect 395632 524 395660 564
rect 396092 564 396396 592
rect 396092 524 396120 564
rect 396258 524 396264 536
rect 395632 496 396120 524
rect 396219 496 396264 524
rect 396258 484 396264 496
rect 396316 484 396322 536
rect 396368 524 396396 564
rect 396534 552 396540 604
rect 396592 552 396598 604
rect 397730 592 397736 604
rect 397691 564 397736 592
rect 397730 552 397736 564
rect 397788 552 397794 604
rect 398834 552 398840 604
rect 398892 592 398898 604
rect 409064 592 409092 632
rect 410794 620 410800 632
rect 410852 620 410858 672
rect 414290 620 414296 672
rect 414348 620 414354 672
rect 414934 660 414940 672
rect 414895 632 414940 660
rect 414934 620 414940 632
rect 414992 620 414998 672
rect 415210 660 415216 672
rect 415171 632 415216 660
rect 415210 620 415216 632
rect 415268 620 415274 672
rect 416038 620 416044 672
rect 416096 660 416102 672
rect 416746 660 416774 836
rect 428461 833 428473 836
rect 428507 833 428519 867
rect 428461 827 428519 833
rect 430577 867 430635 873
rect 430577 833 430589 867
rect 430623 864 430635 867
rect 448241 867 448299 873
rect 448241 864 448253 867
rect 430623 836 434760 864
rect 430623 833 430635 836
rect 430577 827 430635 833
rect 425057 799 425115 805
rect 425057 765 425069 799
rect 425103 796 425115 799
rect 425103 768 434392 796
rect 425103 765 425115 768
rect 425057 759 425115 765
rect 430546 700 432644 728
rect 416096 632 416774 660
rect 417237 663 417295 669
rect 416096 620 416102 632
rect 417237 629 417249 663
rect 417283 660 417295 663
rect 424962 660 424968 672
rect 417283 632 424968 660
rect 417283 629 417295 632
rect 417237 623 417295 629
rect 424962 620 424968 632
rect 425020 620 425026 672
rect 426986 620 426992 672
rect 427044 660 427050 672
rect 428458 660 428464 672
rect 427044 632 428136 660
rect 428419 632 428464 660
rect 427044 620 427050 632
rect 416682 592 416688 604
rect 398892 564 409092 592
rect 409156 564 416688 592
rect 398892 552 398898 564
rect 402698 524 402704 536
rect 396368 496 402704 524
rect 402698 484 402704 496
rect 402756 484 402762 536
rect 404538 484 404544 536
rect 404596 524 404602 536
rect 409156 524 409184 564
rect 416682 552 416688 564
rect 416740 552 416746 604
rect 417329 595 417387 601
rect 417329 561 417341 595
rect 417375 592 417387 595
rect 423677 595 423735 601
rect 423677 592 423689 595
rect 417375 564 423689 592
rect 417375 561 417387 564
rect 417329 555 417387 561
rect 423677 561 423689 564
rect 423723 561 423735 595
rect 423677 555 423735 561
rect 423766 552 423772 604
rect 423824 552 423830 604
rect 423861 595 423919 601
rect 423861 561 423873 595
rect 423907 592 423919 595
rect 426158 592 426164 604
rect 423907 564 426164 592
rect 423907 561 423919 564
rect 423861 555 423919 561
rect 426158 552 426164 564
rect 426216 552 426222 604
rect 427262 592 427268 604
rect 427223 564 427268 592
rect 427262 552 427268 564
rect 427320 552 427326 604
rect 427998 592 428004 604
rect 427959 564 428004 592
rect 427998 552 428004 564
rect 428056 552 428062 604
rect 428108 592 428136 632
rect 428458 620 428464 632
rect 428516 620 428522 672
rect 430546 592 430574 700
rect 431862 660 431868 672
rect 431823 632 431868 660
rect 431862 620 431868 632
rect 431920 620 431926 672
rect 432046 592 432052 604
rect 428108 564 430574 592
rect 432007 564 432052 592
rect 432046 552 432052 564
rect 432104 552 432110 604
rect 432616 592 432644 700
rect 434364 660 434392 768
rect 434732 672 434760 836
rect 437446 836 448253 864
rect 437446 728 437474 836
rect 448241 833 448253 836
rect 448287 833 448299 867
rect 448241 827 448299 833
rect 448885 867 448943 873
rect 448885 833 448897 867
rect 448931 864 448943 867
rect 454497 867 454555 873
rect 454497 864 454509 867
rect 448931 836 454509 864
rect 448931 833 448943 836
rect 448885 827 448943 833
rect 454497 833 454509 836
rect 454543 833 454555 867
rect 454497 827 454555 833
rect 464893 867 464951 873
rect 464893 833 464905 867
rect 464939 864 464951 867
rect 469677 867 469735 873
rect 469677 864 469689 867
rect 464939 836 469689 864
rect 464939 833 464951 836
rect 464893 827 464951 833
rect 469677 833 469689 836
rect 469723 833 469735 867
rect 478846 864 478874 904
rect 486605 901 486617 904
rect 486651 901 486663 935
rect 486605 895 486663 901
rect 491389 935 491447 941
rect 491389 901 491401 935
rect 491435 932 491447 935
rect 514665 935 514723 941
rect 491435 904 500954 932
rect 491435 901 491447 904
rect 491389 895 491447 901
rect 469677 827 469735 833
rect 473326 836 478874 864
rect 483109 867 483167 873
rect 438397 799 438455 805
rect 438397 765 438409 799
rect 438443 796 438455 799
rect 446217 799 446275 805
rect 446217 796 446229 799
rect 438443 768 446229 796
rect 438443 765 438455 768
rect 438397 759 438455 765
rect 446217 765 446229 768
rect 446263 765 446275 799
rect 457165 799 457223 805
rect 457165 796 457177 799
rect 446217 759 446275 765
rect 449176 768 457177 796
rect 435376 700 437474 728
rect 443273 731 443331 737
rect 435376 672 435404 700
rect 443273 697 443285 731
rect 443319 728 443331 731
rect 449176 728 449204 768
rect 457165 765 457177 768
rect 457211 765 457223 799
rect 457165 759 457223 765
rect 461412 768 471008 796
rect 461305 731 461363 737
rect 461305 728 461317 731
rect 443319 700 449204 728
rect 449636 700 461317 728
rect 443319 697 443331 700
rect 443273 691 443331 697
rect 449636 672 449664 700
rect 461305 697 461317 700
rect 461351 697 461363 731
rect 461305 691 461363 697
rect 434438 660 434444 672
rect 434364 632 434444 660
rect 434438 620 434444 632
rect 434496 620 434502 672
rect 434714 620 434720 672
rect 434772 620 434778 672
rect 435358 620 435364 672
rect 435416 620 435422 672
rect 435542 660 435548 672
rect 435503 632 435548 660
rect 435542 620 435548 632
rect 435600 620 435606 672
rect 437474 620 437480 672
rect 437532 660 437538 672
rect 449529 663 449587 669
rect 449529 660 449541 663
rect 437532 632 449541 660
rect 437532 620 437538 632
rect 449529 629 449541 632
rect 449575 629 449587 663
rect 449529 623 449587 629
rect 449618 620 449624 672
rect 449676 620 449682 672
rect 451274 660 451280 672
rect 451235 632 451280 660
rect 451274 620 451280 632
rect 451332 620 451338 672
rect 454218 660 454224 672
rect 454179 632 454224 660
rect 454218 620 454224 632
rect 454276 620 454282 672
rect 455690 660 455696 672
rect 455651 632 455696 660
rect 455690 620 455696 632
rect 455748 620 455754 672
rect 456794 620 456800 672
rect 456852 660 456858 672
rect 461412 660 461440 768
rect 468481 731 468539 737
rect 468481 728 468493 731
rect 463620 700 468493 728
rect 463620 672 463648 700
rect 468481 697 468493 700
rect 468527 697 468539 731
rect 468481 691 468539 697
rect 468757 731 468815 737
rect 468757 697 468769 731
rect 468803 728 468815 731
rect 470873 731 470931 737
rect 470873 728 470885 731
rect 468803 700 470885 728
rect 468803 697 468815 700
rect 468757 691 468815 697
rect 470873 697 470885 700
rect 470919 697 470931 731
rect 470873 691 470931 697
rect 461946 660 461952 672
rect 456852 632 461440 660
rect 461504 632 461952 660
rect 456852 620 456858 632
rect 440326 592 440332 604
rect 432616 564 440332 592
rect 440326 552 440332 564
rect 440384 552 440390 604
rect 441522 592 441528 604
rect 441483 564 441528 592
rect 441522 552 441528 564
rect 441580 552 441586 604
rect 442626 592 442632 604
rect 442587 564 442632 592
rect 442626 552 442632 564
rect 442684 552 442690 604
rect 443270 592 443276 604
rect 443231 564 443276 592
rect 443270 552 443276 564
rect 443328 552 443334 604
rect 445018 592 445024 604
rect 444979 564 445024 592
rect 445018 552 445024 564
rect 445076 552 445082 604
rect 446214 592 446220 604
rect 446175 564 446220 592
rect 446214 552 446220 564
rect 446272 552 446278 604
rect 446674 592 446680 604
rect 446635 564 446680 592
rect 446674 552 446680 564
rect 446732 552 446738 604
rect 447410 592 447416 604
rect 447371 564 447416 592
rect 447410 552 447416 564
rect 447468 552 447474 604
rect 452289 595 452347 601
rect 452289 592 452301 595
rect 448072 564 452301 592
rect 404596 496 409184 524
rect 404596 484 404602 496
rect 409230 484 409236 536
rect 409288 524 409294 536
rect 421006 524 421012 536
rect 409288 496 421012 524
rect 409288 484 409294 496
rect 421006 484 421012 496
rect 421064 484 421070 536
rect 422386 524 422392 536
rect 422347 496 422392 524
rect 422386 484 422392 496
rect 422444 484 422450 536
rect 422481 527 422539 533
rect 422481 493 422493 527
rect 422527 524 422539 527
rect 423784 524 423812 552
rect 422527 496 423812 524
rect 424505 527 424563 533
rect 422527 493 422539 496
rect 422481 487 422539 493
rect 424505 493 424517 527
rect 424551 524 424563 527
rect 430577 527 430635 533
rect 430577 524 430589 527
rect 424551 496 430589 524
rect 424551 493 424563 496
rect 424505 487 424563 493
rect 430577 493 430589 496
rect 430623 493 430635 527
rect 430577 487 430635 493
rect 430666 484 430672 536
rect 430724 524 430730 536
rect 430724 496 437474 524
rect 430724 484 430730 496
rect 383160 428 387380 456
rect 383160 416 383166 428
rect 388806 416 388812 468
rect 388864 456 388870 468
rect 388864 428 391934 456
rect 388864 416 388870 428
rect 389453 391 389511 397
rect 389453 388 389465 391
rect 380912 360 389465 388
rect 379885 351 379943 357
rect 389453 357 389465 360
rect 389499 357 389511 391
rect 389453 351 389511 357
rect 367664 292 368336 320
rect 346820 224 350534 252
rect 346820 212 346826 224
rect 351270 212 351276 264
rect 351328 252 351334 264
rect 351328 224 357296 252
rect 351328 212 351334 224
rect 324096 156 324314 184
rect 324096 144 324102 156
rect 325142 144 325148 196
rect 325200 184 325206 196
rect 333606 184 333612 196
rect 325200 156 333612 184
rect 325200 144 325206 156
rect 333606 144 333612 156
rect 333664 144 333670 196
rect 338298 144 338304 196
rect 338356 184 338362 196
rect 338356 156 344508 184
rect 338356 144 338362 156
rect 184348 88 184934 116
rect 184348 76 184354 88
rect 185486 76 185492 128
rect 185544 116 185550 128
rect 188246 116 188252 128
rect 185544 88 188252 116
rect 185544 76 185550 88
rect 188246 76 188252 88
rect 188304 76 188310 128
rect 213822 76 213828 128
rect 213880 116 213886 128
rect 217870 116 217876 128
rect 213880 88 217876 116
rect 213880 76 213886 88
rect 217870 76 217876 88
rect 217928 76 217934 128
rect 329742 76 329748 128
rect 329800 116 329806 128
rect 338669 119 338727 125
rect 338669 116 338681 119
rect 329800 88 338681 116
rect 329800 76 329806 88
rect 338669 85 338681 88
rect 338715 85 338727 119
rect 338669 79 338727 85
rect 339494 76 339500 128
rect 339552 116 339558 128
rect 344480 116 344508 156
rect 345566 144 345572 196
rect 345624 184 345630 196
rect 354950 184 354956 196
rect 345624 156 354956 184
rect 345624 144 345630 156
rect 354950 144 354956 156
rect 355008 144 355014 196
rect 355781 187 355839 193
rect 355781 153 355793 187
rect 355827 184 355839 187
rect 357158 184 357164 196
rect 355827 156 357164 184
rect 355827 153 355839 156
rect 355781 147 355839 153
rect 357158 144 357164 156
rect 357216 144 357222 196
rect 357268 184 357296 224
rect 358078 212 358084 264
rect 358136 252 358142 264
rect 368201 255 368259 261
rect 368201 252 368213 255
rect 358136 224 368213 252
rect 358136 212 358142 224
rect 368201 221 368213 224
rect 368247 221 368259 255
rect 368308 252 368336 292
rect 369026 280 369032 332
rect 369084 320 369090 332
rect 379790 320 379796 332
rect 369084 292 379796 320
rect 369084 280 369090 292
rect 379790 280 379796 292
rect 379848 280 379854 332
rect 380802 280 380808 332
rect 380860 320 380866 332
rect 391566 320 391572 332
rect 380860 292 391572 320
rect 380860 280 380866 292
rect 391566 280 391572 292
rect 391624 280 391630 332
rect 373902 252 373908 264
rect 368308 224 373908 252
rect 368201 215 368259 221
rect 373902 212 373908 224
rect 373960 212 373966 264
rect 377398 212 377404 264
rect 377456 252 377462 264
rect 380621 255 380679 261
rect 380621 252 380633 255
rect 377456 224 380633 252
rect 377456 212 377462 224
rect 380621 221 380633 224
rect 380667 221 380679 255
rect 391906 252 391934 428
rect 395614 416 395620 468
rect 395672 456 395678 468
rect 397825 459 397883 465
rect 395672 428 397454 456
rect 395672 416 395678 428
rect 393222 388 393228 400
rect 393183 360 393228 388
rect 393222 348 393228 360
rect 393280 348 393286 400
rect 395522 388 395528 400
rect 395483 360 395528 388
rect 395522 348 395528 360
rect 395580 348 395586 400
rect 397426 388 397454 428
rect 397825 425 397837 459
rect 397871 456 397883 459
rect 403069 459 403127 465
rect 403069 456 403081 459
rect 397871 428 403081 456
rect 397871 425 397883 428
rect 397825 419 397883 425
rect 403069 425 403081 428
rect 403115 425 403127 459
rect 403069 419 403127 425
rect 403434 416 403440 468
rect 403492 456 403498 468
rect 415302 456 415308 468
rect 403492 428 415308 456
rect 403492 416 403498 428
rect 415302 416 415308 428
rect 415360 416 415366 468
rect 417142 416 417148 468
rect 417200 456 417206 468
rect 429470 456 429476 468
rect 417200 428 429476 456
rect 417200 416 417206 428
rect 429470 416 429476 428
rect 429528 416 429534 468
rect 432966 456 432972 468
rect 430546 428 432972 456
rect 406841 391 406899 397
rect 406841 388 406853 391
rect 397426 360 406853 388
rect 406841 357 406853 360
rect 406887 357 406899 391
rect 406841 351 406899 357
rect 406930 348 406936 400
rect 406988 388 406994 400
rect 418798 388 418804 400
rect 406988 360 418804 388
rect 406988 348 406994 360
rect 418798 348 418804 360
rect 418856 348 418862 400
rect 420546 348 420552 400
rect 420604 388 420610 400
rect 430546 388 430574 428
rect 432966 416 432972 428
rect 433024 416 433030 468
rect 437446 456 437474 496
rect 438762 484 438768 536
rect 438820 524 438826 536
rect 448072 524 448100 564
rect 452289 561 452301 564
rect 452335 561 452347 595
rect 454494 592 454500 604
rect 454455 564 454500 592
rect 452289 555 452347 561
rect 454494 552 454500 564
rect 454552 552 454558 604
rect 455049 595 455107 601
rect 455049 561 455061 595
rect 455095 592 455107 595
rect 460382 592 460388 604
rect 455095 564 460388 592
rect 455095 561 455107 564
rect 455049 555 455107 561
rect 460382 552 460388 564
rect 460440 552 460446 604
rect 461305 595 461363 601
rect 461305 561 461317 595
rect 461351 592 461363 595
rect 461504 592 461532 632
rect 461946 620 461952 632
rect 462004 620 462010 672
rect 463142 660 463148 672
rect 463103 632 463148 660
rect 463142 620 463148 632
rect 463200 620 463206 672
rect 463602 620 463608 672
rect 463660 620 463666 672
rect 464890 660 464896 672
rect 464851 632 464896 660
rect 464890 620 464896 632
rect 464948 620 464954 672
rect 464985 663 465043 669
rect 464985 629 464997 663
rect 465031 660 465043 663
rect 468386 660 468392 672
rect 465031 632 467696 660
rect 468347 632 468392 660
rect 465031 629 465043 632
rect 464985 623 465043 629
rect 461351 564 461532 592
rect 461351 561 461363 564
rect 461305 555 461363 561
rect 461762 552 461768 604
rect 461820 592 461826 604
rect 467466 592 467472 604
rect 461820 564 467472 592
rect 461820 552 461826 564
rect 467466 552 467472 564
rect 467524 552 467530 604
rect 467668 592 467696 632
rect 468386 620 468392 632
rect 468444 620 468450 672
rect 469214 620 469220 672
rect 469272 660 469278 672
rect 470980 660 471008 768
rect 471054 660 471060 672
rect 469272 632 469317 660
rect 470980 632 471060 660
rect 469272 620 469278 632
rect 471054 620 471060 632
rect 471112 620 471118 672
rect 471698 620 471704 672
rect 471756 660 471762 672
rect 473326 660 473354 836
rect 483109 833 483121 867
rect 483155 864 483167 867
rect 483155 836 498240 864
rect 483155 833 483167 836
rect 483109 827 483167 833
rect 479613 799 479671 805
rect 479613 765 479625 799
rect 479659 796 479671 799
rect 498105 799 498163 805
rect 498105 796 498117 799
rect 479659 768 488534 796
rect 479659 765 479671 768
rect 479613 759 479671 765
rect 483937 731 483995 737
rect 483937 697 483949 731
rect 483983 728 483995 731
rect 488506 728 488534 768
rect 491312 768 498117 796
rect 491113 731 491171 737
rect 491113 728 491125 731
rect 483983 700 487844 728
rect 488506 700 491125 728
rect 483983 697 483995 700
rect 483937 691 483995 697
rect 487816 672 487844 700
rect 491113 697 491125 700
rect 491159 697 491171 731
rect 491113 691 491171 697
rect 473998 660 474004 672
rect 471756 632 473354 660
rect 473959 632 474004 660
rect 471756 620 471762 632
rect 473998 620 474004 632
rect 474056 620 474062 672
rect 476758 660 476764 672
rect 476719 632 476764 660
rect 476758 620 476764 632
rect 476816 620 476822 672
rect 476942 660 476948 672
rect 476903 632 476948 660
rect 476942 620 476948 632
rect 477000 620 477006 672
rect 485130 660 485136 672
rect 478846 632 485136 660
rect 473446 592 473452 604
rect 467668 564 473452 592
rect 473446 552 473452 564
rect 473504 552 473510 604
rect 475102 552 475108 604
rect 475160 592 475166 604
rect 478846 592 478874 632
rect 485130 620 485136 632
rect 485188 620 485194 672
rect 486602 660 486608 672
rect 486563 632 486608 660
rect 486602 620 486608 632
rect 486660 620 486666 672
rect 487798 620 487804 672
rect 487856 620 487862 672
rect 488534 620 488540 672
rect 488592 660 488598 672
rect 491205 663 491263 669
rect 491205 660 491217 663
rect 488592 632 491217 660
rect 488592 620 488598 632
rect 491205 629 491217 632
rect 491251 629 491263 663
rect 491205 623 491263 629
rect 479610 592 479616 604
rect 475160 564 478874 592
rect 479571 564 479616 592
rect 475160 552 475166 564
rect 479610 552 479616 564
rect 479668 552 479674 604
rect 483106 592 483112 604
rect 483067 564 483112 592
rect 483106 552 483112 564
rect 483164 552 483170 604
rect 483750 592 483756 604
rect 483711 564 483756 592
rect 483750 552 483756 564
rect 483808 552 483814 604
rect 484026 592 484032 604
rect 483987 564 484032 592
rect 484026 552 484032 564
rect 484084 552 484090 604
rect 485222 552 485228 604
rect 485280 552 485286 604
rect 486326 552 486332 604
rect 486384 592 486390 604
rect 486384 564 487154 592
rect 486384 552 486390 564
rect 448238 524 448244 536
rect 438820 496 448100 524
rect 448199 496 448244 524
rect 438820 484 438826 496
rect 448238 484 448244 496
rect 448296 484 448302 536
rect 449529 527 449587 533
rect 449529 493 449541 527
rect 449575 524 449587 527
rect 450630 524 450636 536
rect 449575 496 450636 524
rect 449575 493 449587 496
rect 449529 487 449587 493
rect 450630 484 450636 496
rect 450688 484 450694 536
rect 458266 524 458272 536
rect 454006 496 458272 524
rect 443638 456 443644 468
rect 437446 428 443644 456
rect 443638 416 443644 428
rect 443696 416 443702 468
rect 444466 416 444472 468
rect 444524 456 444530 468
rect 454006 456 454034 496
rect 458266 484 458272 496
rect 458324 484 458330 536
rect 459002 484 459008 536
rect 459060 524 459066 536
rect 464985 527 465043 533
rect 464985 524 464997 527
rect 459060 496 464997 524
rect 459060 484 459066 496
rect 464985 493 464997 496
rect 465031 493 465043 527
rect 467190 524 467196 536
rect 467151 496 467196 524
rect 464985 487 465043 493
rect 467190 484 467196 496
rect 467248 484 467254 536
rect 468294 484 468300 536
rect 468352 524 468358 536
rect 469490 524 469496 536
rect 468352 496 469496 524
rect 468352 484 468358 496
rect 469490 484 469496 496
rect 469548 484 469554 536
rect 469677 527 469735 533
rect 469677 493 469689 527
rect 469723 524 469735 527
rect 479521 527 479579 533
rect 479521 524 479533 527
rect 469723 496 479533 524
rect 469723 493 469735 496
rect 469677 487 469735 493
rect 479521 493 479533 496
rect 479567 493 479579 527
rect 479521 487 479579 493
rect 480806 484 480812 536
rect 480864 524 480870 536
rect 484949 527 485007 533
rect 484949 524 484961 527
rect 480864 496 484961 524
rect 480864 484 480870 496
rect 484949 493 484961 496
rect 484995 493 485007 527
rect 484949 487 485007 493
rect 457162 456 457168 468
rect 444524 428 454034 456
rect 457123 428 457168 456
rect 444524 416 444530 428
rect 457162 416 457168 428
rect 457220 416 457226 468
rect 457898 416 457904 468
rect 457956 456 457962 468
rect 471974 456 471980 468
rect 457956 428 471980 456
rect 457956 416 457962 428
rect 471974 416 471980 428
rect 472032 416 472038 468
rect 472802 416 472808 468
rect 472860 456 472866 468
rect 483937 459 483995 465
rect 483937 456 483949 459
rect 472860 428 483949 456
rect 472860 416 472866 428
rect 483937 425 483949 428
rect 483983 425 483995 459
rect 485041 459 485099 465
rect 485041 456 485053 459
rect 483937 419 483995 425
rect 484044 428 485053 456
rect 437566 388 437572 400
rect 420604 360 430574 388
rect 432616 360 437572 388
rect 420604 348 420610 360
rect 396445 323 396503 329
rect 396445 289 396457 323
rect 396491 320 396503 323
rect 397825 323 397883 329
rect 397825 320 397837 323
rect 396491 292 397837 320
rect 396491 289 396503 292
rect 396445 283 396503 289
rect 397825 289 397837 292
rect 397871 289 397883 323
rect 409414 320 409420 332
rect 397825 283 397883 289
rect 400416 292 409420 320
rect 400125 255 400183 261
rect 400125 252 400137 255
rect 391906 224 400137 252
rect 380621 215 380679 221
rect 400125 221 400137 224
rect 400171 221 400183 255
rect 400125 215 400183 221
rect 360838 184 360844 196
rect 357268 156 360844 184
rect 360838 144 360844 156
rect 360896 144 360902 196
rect 366726 144 366732 196
rect 366784 184 366790 196
rect 367741 187 367799 193
rect 367741 184 367753 187
rect 366784 156 367753 184
rect 366784 144 366790 156
rect 367741 153 367753 156
rect 367787 153 367799 187
rect 367741 147 367799 153
rect 367830 144 367836 196
rect 367888 184 367894 196
rect 367888 156 373764 184
rect 367888 144 367894 156
rect 347682 116 347688 128
rect 339552 88 344416 116
rect 344480 88 347688 116
rect 339552 76 339558 88
rect 44082 8 44088 60
rect 44140 48 44146 60
rect 46198 48 46204 60
rect 44140 20 46204 48
rect 44140 8 44146 20
rect 46198 8 46204 20
rect 46256 8 46262 60
rect 215018 8 215024 60
rect 215076 48 215082 60
rect 219434 48 219440 60
rect 215076 20 219440 48
rect 215076 8 215082 20
rect 219434 8 219440 20
rect 219492 8 219498 60
rect 256878 8 256884 60
rect 256936 48 256942 60
rect 262766 48 262772 60
rect 256936 20 262772 48
rect 256936 8 256942 20
rect 262766 8 262772 20
rect 262824 8 262830 60
rect 264882 8 264888 60
rect 264940 48 264946 60
rect 271046 48 271052 60
rect 264940 20 271052 48
rect 264940 8 264946 20
rect 271046 8 271052 20
rect 271104 8 271110 60
rect 293402 8 293408 60
rect 293460 48 293466 60
rect 300486 48 300492 60
rect 293460 20 300492 48
rect 293460 8 293466 20
rect 300486 8 300492 20
rect 300544 8 300550 60
rect 303614 8 303620 60
rect 303672 48 303678 60
rect 310333 51 310391 57
rect 310333 48 310345 51
rect 303672 20 310345 48
rect 303672 8 303678 20
rect 310333 17 310345 20
rect 310379 17 310391 51
rect 310333 11 310391 17
rect 311066 8 311072 60
rect 311124 48 311130 60
rect 319717 51 319775 57
rect 319717 48 319729 51
rect 311124 20 319729 48
rect 311124 8 311130 20
rect 319717 17 319729 20
rect 319763 17 319775 51
rect 319717 11 319775 17
rect 322842 8 322848 60
rect 322900 48 322906 60
rect 331214 48 331220 60
rect 322900 20 331220 48
rect 322900 8 322906 20
rect 331214 8 331220 20
rect 331272 8 331278 60
rect 344388 48 344416 88
rect 347682 76 347688 88
rect 347740 76 347746 128
rect 349430 76 349436 128
rect 349488 76 349494 128
rect 353570 76 353576 128
rect 353628 116 353634 128
rect 363690 116 363696 128
rect 353628 88 363696 116
rect 353628 76 353634 88
rect 363690 76 363696 88
rect 363748 76 363754 128
rect 373736 116 373764 156
rect 373810 144 373816 196
rect 373868 184 373874 196
rect 384574 184 384580 196
rect 373868 156 384580 184
rect 373868 144 373874 156
rect 384574 144 384580 156
rect 384632 144 384638 196
rect 393958 144 393964 196
rect 394016 184 394022 196
rect 396445 187 396503 193
rect 396445 184 396457 187
rect 394016 156 396457 184
rect 394016 144 394022 156
rect 396445 153 396457 156
rect 396491 153 396503 187
rect 396445 147 396503 153
rect 397454 144 397460 196
rect 397512 184 397518 196
rect 400416 184 400444 292
rect 409414 280 409420 292
rect 409472 280 409478 332
rect 410334 280 410340 332
rect 410392 320 410398 332
rect 422754 320 422760 332
rect 410392 292 422760 320
rect 410392 280 410398 292
rect 422754 280 422760 292
rect 422812 280 422818 332
rect 423490 280 423496 332
rect 423548 320 423554 332
rect 424505 323 424563 329
rect 424505 320 424517 323
rect 423548 292 424517 320
rect 423548 280 423554 292
rect 424505 289 424517 292
rect 424551 289 424563 323
rect 424505 283 424563 289
rect 424686 280 424692 332
rect 424744 320 424750 332
rect 432616 320 432644 360
rect 437566 348 437572 360
rect 437624 348 437630 400
rect 442166 348 442172 400
rect 442224 388 442230 400
rect 455693 391 455751 397
rect 455693 388 455705 391
rect 442224 360 455705 388
rect 442224 348 442230 360
rect 455693 357 455705 360
rect 455739 357 455751 391
rect 455693 351 455751 357
rect 460198 348 460204 400
rect 460256 388 460262 400
rect 474366 388 474372 400
rect 460256 360 474372 388
rect 460256 348 460262 360
rect 474366 348 474372 360
rect 474424 348 474430 400
rect 479518 388 479524 400
rect 479479 360 479524 388
rect 479518 348 479524 360
rect 479576 348 479582 400
rect 481450 348 481456 400
rect 481508 388 481514 400
rect 484044 388 484072 428
rect 485041 425 485053 428
rect 485087 425 485099 459
rect 485041 419 485099 425
rect 485240 388 485268 552
rect 487126 524 487154 564
rect 487522 552 487528 604
rect 487580 592 487586 604
rect 491312 592 491340 768
rect 498105 765 498117 768
rect 498151 765 498163 799
rect 498105 759 498163 765
rect 498212 672 498240 836
rect 492122 660 492128 672
rect 492083 632 492128 660
rect 492122 620 492128 632
rect 492180 620 492186 672
rect 493318 660 493324 672
rect 493279 632 493324 660
rect 493318 620 493324 632
rect 493376 620 493382 672
rect 497826 660 497832 672
rect 497787 632 497832 660
rect 497826 620 497832 632
rect 497884 620 497890 672
rect 498194 620 498200 672
rect 498252 620 498258 672
rect 498930 620 498936 672
rect 498988 660 498994 672
rect 499485 663 499543 669
rect 499485 660 499497 663
rect 498988 632 499497 660
rect 498988 620 498994 632
rect 499485 629 499497 632
rect 499531 629 499543 663
rect 500926 660 500954 904
rect 514665 901 514677 935
rect 514711 932 514723 935
rect 531317 935 531375 941
rect 531317 932 531329 935
rect 514711 904 531329 932
rect 514711 901 514723 904
rect 514665 895 514723 901
rect 531317 901 531329 904
rect 531363 901 531375 935
rect 531317 895 531375 901
rect 531869 935 531927 941
rect 531869 901 531881 935
rect 531915 932 531927 935
rect 531915 904 546494 932
rect 531915 901 531927 904
rect 531869 895 531927 901
rect 523037 867 523095 873
rect 523037 864 523049 867
rect 507826 836 523049 864
rect 504174 660 504180 672
rect 500926 632 504180 660
rect 499485 623 499543 629
rect 504174 620 504180 632
rect 504232 620 504238 672
rect 504634 660 504640 672
rect 504595 632 504640 660
rect 504634 620 504640 632
rect 504692 620 504698 672
rect 506934 620 506940 672
rect 506992 660 506998 672
rect 507826 660 507854 836
rect 523037 833 523049 836
rect 523083 833 523095 867
rect 523037 827 523095 833
rect 523957 867 524015 873
rect 523957 833 523969 867
rect 524003 864 524015 867
rect 540793 867 540851 873
rect 540793 864 540805 867
rect 524003 836 540805 864
rect 524003 833 524015 836
rect 523957 827 524015 833
rect 540793 833 540805 836
rect 540839 833 540851 867
rect 540793 827 540851 833
rect 530121 799 530179 805
rect 530121 796 530133 799
rect 513300 768 530133 796
rect 513300 672 513328 768
rect 530121 765 530133 768
rect 530167 765 530179 799
rect 542173 799 542231 805
rect 542173 796 542185 799
rect 530121 759 530179 765
rect 538876 768 542185 796
rect 513929 731 513987 737
rect 513929 697 513941 731
rect 513975 728 513987 731
rect 513975 700 519584 728
rect 513975 697 513987 700
rect 513929 691 513987 697
rect 519556 672 519584 700
rect 520108 700 532694 728
rect 520108 672 520136 700
rect 506992 632 507854 660
rect 506992 620 506998 632
rect 507946 620 507952 672
rect 508004 660 508010 672
rect 508590 660 508596 672
rect 508004 632 508049 660
rect 508551 632 508596 660
rect 508004 620 508010 632
rect 508590 620 508596 632
rect 508648 620 508654 672
rect 509878 660 509884 672
rect 509839 632 509884 660
rect 509878 620 509884 632
rect 509936 620 509942 672
rect 511184 632 512500 660
rect 487580 564 491340 592
rect 487580 552 487586 564
rect 492858 552 492864 604
rect 492916 592 492922 604
rect 493502 592 493508 604
rect 492916 564 493508 592
rect 492916 552 492922 564
rect 493502 552 493508 564
rect 493560 552 493566 604
rect 499390 592 499396 604
rect 499351 564 499396 592
rect 499390 552 499396 564
rect 499448 552 499454 604
rect 501782 552 501788 604
rect 501840 552 501846 604
rect 502978 592 502984 604
rect 502939 564 502984 592
rect 502978 552 502984 564
rect 503036 552 503042 604
rect 501800 524 501828 552
rect 487126 496 501828 524
rect 503441 527 503499 533
rect 503441 493 503453 527
rect 503487 524 503499 527
rect 511184 524 511212 632
rect 512472 604 512500 632
rect 513282 620 513288 672
rect 513340 620 513346 672
rect 513558 660 513564 672
rect 513519 632 513564 660
rect 513558 620 513564 632
rect 513616 620 513622 672
rect 514662 660 514668 672
rect 514623 632 514668 660
rect 514662 620 514668 632
rect 514720 620 514726 672
rect 514754 620 514760 672
rect 514812 660 514818 672
rect 518250 660 518256 672
rect 514812 632 514857 660
rect 518211 632 518256 660
rect 514812 620 514818 632
rect 518250 620 518256 632
rect 518308 620 518314 672
rect 518345 663 518403 669
rect 518345 629 518357 663
rect 518391 660 518403 663
rect 519449 663 519507 669
rect 519449 660 519461 663
rect 518391 632 519461 660
rect 518391 629 518403 632
rect 518345 623 518403 629
rect 519449 629 519461 632
rect 519495 629 519507 663
rect 519449 623 519507 629
rect 519538 620 519544 672
rect 519596 620 519602 672
rect 520090 620 520096 672
rect 520148 620 520154 672
rect 520734 660 520740 672
rect 520695 632 520740 660
rect 520734 620 520740 632
rect 520792 620 520798 672
rect 522850 660 522856 672
rect 522811 632 522856 660
rect 522850 620 522856 632
rect 522908 620 522914 672
rect 523034 660 523040 672
rect 522995 632 523040 660
rect 523034 620 523040 632
rect 523092 620 523098 672
rect 523954 660 523960 672
rect 523915 632 523960 660
rect 523954 620 523960 632
rect 524012 620 524018 672
rect 524230 660 524236 672
rect 524191 632 524236 660
rect 524230 620 524236 632
rect 524288 620 524294 672
rect 525058 620 525064 672
rect 525116 660 525122 672
rect 530213 663 530271 669
rect 530213 660 530225 663
rect 525116 632 530225 660
rect 525116 620 525122 632
rect 530213 629 530225 632
rect 530259 629 530271 663
rect 531866 660 531872 672
rect 531827 632 531872 660
rect 530213 623 530271 629
rect 531866 620 531872 632
rect 531924 620 531930 672
rect 532666 660 532694 700
rect 535822 660 535828 672
rect 532666 632 535828 660
rect 535822 620 535828 632
rect 535880 620 535886 672
rect 538766 660 538772 672
rect 538727 632 538772 660
rect 538766 620 538772 632
rect 538824 620 538830 672
rect 511258 552 511264 604
rect 511316 552 511322 604
rect 512454 552 512460 604
rect 512512 552 512518 604
rect 512549 595 512607 601
rect 512549 561 512561 595
rect 512595 592 512607 595
rect 515950 592 515956 604
rect 512595 564 515956 592
rect 512595 561 512607 564
rect 512549 555 512607 561
rect 515950 552 515956 564
rect 516008 552 516014 604
rect 517054 552 517060 604
rect 517112 592 517118 604
rect 529934 592 529940 604
rect 517112 564 529940 592
rect 517112 552 517118 564
rect 529934 552 529940 564
rect 529992 552 529998 604
rect 530118 592 530124 604
rect 530079 564 530124 592
rect 530118 552 530124 564
rect 530176 552 530182 604
rect 531314 592 531320 604
rect 531275 564 531320 592
rect 531314 552 531320 564
rect 531372 552 531378 604
rect 534534 592 534540 604
rect 534495 564 534540 592
rect 534534 552 534540 564
rect 534592 552 534598 604
rect 503487 496 511212 524
rect 503487 493 503499 496
rect 503441 487 503499 493
rect 488994 456 489000 468
rect 488955 428 489000 456
rect 488994 416 489000 428
rect 489052 416 489058 468
rect 491113 459 491171 465
rect 491113 425 491125 459
rect 491159 456 491171 459
rect 491478 456 491484 468
rect 491159 428 491484 456
rect 491159 425 491171 428
rect 491113 419 491171 425
rect 491478 416 491484 428
rect 491536 416 491542 468
rect 495526 416 495532 468
rect 495584 456 495590 468
rect 511276 456 511304 552
rect 518345 527 518403 533
rect 518345 524 518357 527
rect 495584 428 511304 456
rect 512104 496 518357 524
rect 495584 416 495590 428
rect 481508 360 484072 388
rect 484136 360 485268 388
rect 481508 348 481514 360
rect 424744 292 432644 320
rect 432693 323 432751 329
rect 424744 280 424750 292
rect 432693 289 432705 323
rect 432739 320 432751 323
rect 442629 323 442687 329
rect 442629 320 442641 323
rect 432739 292 442641 320
rect 432739 289 432751 292
rect 432693 283 432751 289
rect 442629 289 442641 292
rect 442675 289 442687 323
rect 442629 283 442687 289
rect 445570 280 445576 332
rect 445628 320 445634 332
rect 449253 323 449311 329
rect 445628 292 449204 320
rect 445628 280 445634 292
rect 401134 212 401140 264
rect 401192 252 401198 264
rect 401192 224 404768 252
rect 401192 212 401198 224
rect 397512 156 400444 184
rect 403069 187 403127 193
rect 397512 144 397518 156
rect 403069 153 403081 187
rect 403115 184 403127 187
rect 404740 184 404768 224
rect 408126 212 408132 264
rect 408184 252 408190 264
rect 419902 252 419908 264
rect 408184 224 419908 252
rect 408184 212 408190 224
rect 419902 212 419908 224
rect 419960 212 419966 264
rect 421742 212 421748 264
rect 421800 252 421806 264
rect 424965 255 425023 261
rect 424965 252 424977 255
rect 421800 224 424977 252
rect 421800 212 421806 224
rect 424965 221 424977 224
rect 425011 221 425023 255
rect 424965 215 425023 221
rect 425790 212 425796 264
rect 425848 252 425854 264
rect 433337 255 433395 261
rect 433337 252 433349 255
rect 425848 224 433349 252
rect 425848 212 425854 224
rect 433337 221 433349 224
rect 433383 221 433395 255
rect 433337 215 433395 221
rect 433521 255 433579 261
rect 433521 221 433533 255
rect 433567 252 433579 255
rect 438762 252 438768 264
rect 433567 224 438768 252
rect 433567 221 433579 224
rect 433521 215 433579 221
rect 438762 212 438768 224
rect 438820 212 438826 264
rect 449069 255 449127 261
rect 449069 252 449081 255
rect 440206 224 449081 252
rect 412910 184 412916 196
rect 403115 156 404676 184
rect 404740 156 412916 184
rect 403115 153 403127 156
rect 403069 147 403127 153
rect 378686 116 378692 128
rect 373736 88 378692 116
rect 378686 76 378692 88
rect 378744 76 378750 128
rect 379514 76 379520 128
rect 379572 116 379578 128
rect 390278 116 390284 128
rect 379572 88 390284 116
rect 379572 76 379578 88
rect 390278 76 390284 88
rect 390336 76 390342 128
rect 393314 76 393320 128
rect 393372 116 393378 128
rect 404538 116 404544 128
rect 393372 88 404544 116
rect 393372 76 393378 88
rect 404538 76 404544 88
rect 404596 76 404602 128
rect 404648 116 404676 156
rect 412910 144 412916 156
rect 412968 144 412974 196
rect 413738 144 413744 196
rect 413796 184 413802 196
rect 417329 187 417387 193
rect 417329 184 417341 187
rect 413796 156 417341 184
rect 413796 144 413802 156
rect 417329 153 417341 156
rect 417375 153 417387 187
rect 417329 147 417387 153
rect 436462 144 436468 196
rect 436520 184 436526 196
rect 440206 184 440234 224
rect 449069 221 449081 224
rect 449115 221 449127 255
rect 449176 252 449204 292
rect 449253 289 449265 323
rect 449299 320 449311 323
rect 449986 320 449992 332
rect 449299 292 449992 320
rect 449299 289 449311 292
rect 449253 283 449311 289
rect 449986 280 449992 292
rect 450044 280 450050 332
rect 452286 320 452292 332
rect 452247 292 452292 320
rect 452286 280 452292 292
rect 452344 280 452350 332
rect 452378 280 452384 332
rect 452436 320 452442 332
rect 465902 320 465908 332
rect 452436 292 465908 320
rect 452436 280 452442 292
rect 465902 280 465908 292
rect 465960 280 465966 332
rect 470594 280 470600 332
rect 470652 320 470658 332
rect 484136 320 484164 360
rect 489730 348 489736 400
rect 489788 388 489794 400
rect 505094 388 505100 400
rect 489788 360 505100 388
rect 489788 348 489794 360
rect 505094 348 505100 360
rect 505152 348 505158 400
rect 505189 391 505247 397
rect 505189 357 505201 391
rect 505235 388 505247 391
rect 509786 388 509792 400
rect 505235 360 509792 388
rect 505235 357 505247 360
rect 505189 351 505247 357
rect 509786 348 509792 360
rect 509844 348 509850 400
rect 510982 348 510988 400
rect 511040 388 511046 400
rect 512104 388 512132 496
rect 518345 493 518357 496
rect 518391 493 518403 527
rect 518345 487 518403 493
rect 519354 484 519360 536
rect 519412 524 519418 536
rect 520090 524 520096 536
rect 519412 496 520096 524
rect 519412 484 519418 496
rect 520090 484 520096 496
rect 520148 484 520154 536
rect 526438 524 526444 536
rect 526399 496 526444 524
rect 526438 484 526444 496
rect 526496 484 526502 536
rect 527174 484 527180 536
rect 527232 524 527238 536
rect 538876 524 538904 768
rect 542173 765 542185 768
rect 542219 765 542231 799
rect 546466 796 546494 904
rect 546466 768 548380 796
rect 542173 759 542231 765
rect 527232 496 538904 524
rect 538968 700 546724 728
rect 527232 484 527238 496
rect 512178 416 512184 468
rect 512236 456 512242 468
rect 528830 456 528836 468
rect 512236 428 528836 456
rect 512236 416 512242 428
rect 528830 416 528836 428
rect 528888 416 528894 468
rect 538968 456 538996 700
rect 546696 672 546724 700
rect 548352 672 548380 768
rect 539134 620 539140 672
rect 539192 660 539198 672
rect 543734 660 543740 672
rect 539192 632 543740 660
rect 539192 620 539198 632
rect 543734 620 543740 632
rect 543792 620 543798 672
rect 546678 620 546684 672
rect 546736 620 546742 672
rect 548334 620 548340 672
rect 548392 620 548398 672
rect 548978 620 548984 672
rect 549036 660 549042 672
rect 551020 660 551048 972
rect 554593 969 554605 1003
rect 554639 1000 554651 1003
rect 557506 1000 557534 1040
rect 563514 1028 563520 1040
rect 563572 1028 563578 1080
rect 554639 972 557534 1000
rect 557997 1003 558055 1009
rect 554639 969 554651 972
rect 554593 963 554651 969
rect 557997 969 558009 1003
rect 558043 1000 558055 1003
rect 569862 1000 569868 1012
rect 558043 972 569868 1000
rect 558043 969 558055 972
rect 557997 963 558055 969
rect 569862 960 569868 972
rect 569920 960 569926 1012
rect 563606 932 563612 944
rect 553366 904 563612 932
rect 553366 796 553394 904
rect 563606 892 563612 904
rect 563664 892 563670 944
rect 565906 864 565912 876
rect 552124 768 553394 796
rect 555344 836 565912 864
rect 549036 632 551048 660
rect 549036 620 549042 632
rect 551186 620 551192 672
rect 551244 660 551250 672
rect 552124 660 552152 768
rect 555344 728 555372 836
rect 565906 824 565912 836
rect 565964 824 565970 876
rect 556065 799 556123 805
rect 556065 765 556077 799
rect 556111 796 556123 799
rect 561125 799 561183 805
rect 561125 796 561137 799
rect 556111 768 561137 796
rect 556111 765 556123 768
rect 556065 759 556123 765
rect 561125 765 561137 768
rect 561171 765 561183 799
rect 561125 759 561183 765
rect 561217 799 561275 805
rect 561217 765 561229 799
rect 561263 796 561275 799
rect 565630 796 565636 808
rect 561263 768 565636 796
rect 561263 765 561275 768
rect 561217 759 561275 765
rect 565630 756 565636 768
rect 565688 756 565694 808
rect 565814 756 565820 808
rect 565872 796 565878 808
rect 568022 796 568028 808
rect 565872 768 568028 796
rect 565872 756 565878 768
rect 568022 756 568028 768
rect 568080 756 568086 808
rect 553366 700 555372 728
rect 555973 731 556031 737
rect 553366 672 553394 700
rect 555973 697 555985 731
rect 556019 728 556031 731
rect 570322 728 570328 740
rect 556019 700 570328 728
rect 556019 697 556031 700
rect 555973 691 556031 697
rect 570322 688 570328 700
rect 570380 688 570386 740
rect 551244 632 552152 660
rect 551244 620 551250 632
rect 553302 620 553308 672
rect 553360 632 553394 672
rect 554590 660 554596 672
rect 554551 632 554596 660
rect 553360 620 553366 632
rect 554590 620 554596 632
rect 554648 620 554654 672
rect 555878 660 555884 672
rect 555839 632 555884 660
rect 555878 620 555884 632
rect 555936 620 555942 672
rect 556065 663 556123 669
rect 556065 629 556077 663
rect 556111 660 556123 663
rect 565814 660 565820 672
rect 556111 632 565820 660
rect 556111 629 556123 632
rect 556065 623 556123 629
rect 565814 620 565820 632
rect 565872 620 565878 672
rect 540790 592 540796 604
rect 540751 564 540796 592
rect 540790 552 540796 564
rect 540848 552 540854 604
rect 541986 552 541992 604
rect 542044 592 542050 604
rect 542265 595 542323 601
rect 542044 564 542089 592
rect 542044 552 542050 564
rect 542265 561 542277 595
rect 542311 592 542323 595
rect 550266 592 550272 604
rect 542311 564 550272 592
rect 542311 561 542323 564
rect 542265 555 542323 561
rect 550266 552 550272 564
rect 550324 552 550330 604
rect 561217 595 561275 601
rect 561217 592 561229 595
rect 550468 564 561229 592
rect 544194 484 544200 536
rect 544252 484 544258 536
rect 547690 484 547696 536
rect 547748 524 547754 536
rect 550468 524 550496 564
rect 561217 561 561229 564
rect 561263 561 561275 595
rect 561398 592 561404 604
rect 561359 564 561404 592
rect 561217 555 561275 561
rect 561398 552 561404 564
rect 561456 552 561462 604
rect 562042 552 562048 604
rect 562100 552 562106 604
rect 573910 592 573916 604
rect 567166 564 573916 592
rect 547748 496 550496 524
rect 550545 527 550603 533
rect 547748 484 547754 496
rect 550545 493 550557 527
rect 550591 524 550603 527
rect 562060 524 562088 552
rect 550591 496 562088 524
rect 550591 493 550603 496
rect 550545 487 550603 493
rect 539778 456 539784 468
rect 532666 428 538996 456
rect 539739 428 539784 456
rect 511040 360 512132 388
rect 519449 391 519507 397
rect 511040 348 511046 360
rect 519449 357 519461 391
rect 519495 388 519507 391
rect 527634 388 527640 400
rect 519495 360 527640 388
rect 519495 357 519507 360
rect 519449 351 519507 357
rect 527634 348 527640 360
rect 527692 348 527698 400
rect 529658 348 529664 400
rect 529716 388 529722 400
rect 532666 388 532694 428
rect 539778 416 539784 428
rect 539836 416 539842 468
rect 542173 459 542231 465
rect 542173 425 542185 459
rect 542219 456 542231 459
rect 544212 456 544240 484
rect 542219 428 544240 456
rect 542219 425 542231 428
rect 542173 419 542231 425
rect 550082 416 550088 468
rect 550140 456 550146 468
rect 550140 428 555740 456
rect 550140 416 550146 428
rect 529716 360 532694 388
rect 529716 348 529722 360
rect 536466 348 536472 400
rect 536524 388 536530 400
rect 553578 388 553584 400
rect 536524 360 553584 388
rect 536524 348 536530 360
rect 553578 348 553584 360
rect 553636 348 553642 400
rect 555712 388 555740 428
rect 555786 416 555792 468
rect 555844 456 555850 468
rect 567166 456 567194 564
rect 573910 552 573916 564
rect 573968 552 573974 604
rect 575106 552 575112 604
rect 575164 552 575170 604
rect 555844 428 567194 456
rect 555844 416 555850 428
rect 556065 391 556123 397
rect 556065 388 556077 391
rect 555712 360 556077 388
rect 556065 357 556077 360
rect 556111 357 556123 391
rect 556065 351 556123 357
rect 556890 348 556896 400
rect 556948 388 556954 400
rect 575124 388 575152 552
rect 556948 360 575152 388
rect 556948 348 556954 360
rect 490190 320 490196 332
rect 470652 292 484164 320
rect 484780 292 490196 320
rect 470652 280 470658 292
rect 459370 252 459376 264
rect 449176 224 459376 252
rect 449069 215 449127 221
rect 459370 212 459376 224
rect 459428 212 459434 264
rect 461394 212 461400 264
rect 461452 252 461458 264
rect 475470 252 475476 264
rect 461452 224 475476 252
rect 461452 212 461458 224
rect 475470 212 475476 224
rect 475528 212 475534 264
rect 436520 156 440234 184
rect 436520 144 436526 156
rect 441062 144 441068 196
rect 441120 184 441126 196
rect 448885 187 448943 193
rect 448885 184 448897 187
rect 441120 156 448897 184
rect 441120 144 441126 156
rect 448885 153 448897 156
rect 448931 153 448943 187
rect 448885 147 448943 153
rect 448974 144 448980 196
rect 449032 184 449038 196
rect 462498 184 462504 196
rect 449032 156 462504 184
rect 449032 144 449038 156
rect 462498 144 462504 156
rect 462556 144 462562 196
rect 465994 144 466000 196
rect 466052 184 466058 196
rect 480714 184 480720 196
rect 466052 156 480720 184
rect 466052 144 466058 156
rect 480714 144 480720 156
rect 480772 144 480778 196
rect 405734 116 405740 128
rect 404648 88 405740 116
rect 405734 76 405740 88
rect 405792 76 405798 128
rect 411622 116 411628 128
rect 408466 88 411628 116
rect 349448 48 349476 76
rect 344388 20 349476 48
rect 350166 8 350172 60
rect 350224 48 350230 60
rect 359734 48 359740 60
rect 350224 20 359740 48
rect 350224 8 350230 20
rect 359734 8 359740 20
rect 359792 8 359798 60
rect 361482 8 361488 60
rect 361540 48 361546 60
rect 371878 48 371884 60
rect 361540 20 371884 48
rect 361540 8 361546 20
rect 371878 8 371884 20
rect 371936 8 371942 60
rect 376294 8 376300 60
rect 376352 48 376358 60
rect 386966 48 386972 60
rect 376352 20 386972 48
rect 376352 8 376358 20
rect 386966 8 386972 20
rect 387024 8 387030 60
rect 387610 8 387616 60
rect 387668 48 387674 60
rect 399110 48 399116 60
rect 387668 20 399116 48
rect 387668 8 387674 20
rect 399110 8 399116 20
rect 399168 8 399174 60
rect 399938 8 399944 60
rect 399996 48 400002 60
rect 408466 48 408494 88
rect 411622 76 411628 88
rect 411680 76 411686 128
rect 412634 76 412640 128
rect 412692 116 412698 128
rect 417237 119 417295 125
rect 417237 116 417249 119
rect 412692 88 417249 116
rect 412692 76 412698 88
rect 417237 85 417249 88
rect 417283 85 417295 119
rect 417237 79 417295 85
rect 419442 76 419448 128
rect 419500 116 419506 128
rect 432049 119 432107 125
rect 432049 116 432061 119
rect 419500 88 432061 116
rect 419500 76 419506 88
rect 432049 85 432061 88
rect 432095 85 432107 119
rect 432049 79 432107 85
rect 434254 76 434260 128
rect 434312 116 434318 128
rect 447413 119 447471 125
rect 447413 116 447425 119
rect 434312 88 447425 116
rect 434312 76 434318 88
rect 447413 85 447425 88
rect 447459 85 447471 119
rect 447413 79 447471 85
rect 447870 76 447876 128
rect 447928 116 447934 128
rect 459554 116 459560 128
rect 447928 88 459560 116
rect 447928 76 447934 88
rect 459554 76 459560 88
rect 459612 76 459618 128
rect 462406 76 462412 128
rect 462464 116 462470 128
rect 476945 119 477003 125
rect 476945 116 476957 119
rect 462464 88 476957 116
rect 462464 76 462470 88
rect 476945 85 476957 88
rect 476991 85 477003 119
rect 476945 79 477003 85
rect 477402 76 477408 128
rect 477460 116 477466 128
rect 484780 116 484808 292
rect 490190 280 490196 292
rect 490248 280 490254 332
rect 490926 280 490932 332
rect 490984 320 490990 332
rect 506198 320 506204 332
rect 490984 292 506204 320
rect 490984 280 490990 292
rect 506198 280 506204 292
rect 506256 280 506262 332
rect 507302 320 507308 332
rect 507263 292 507308 320
rect 507302 280 507308 292
rect 507360 280 507366 332
rect 509234 280 509240 332
rect 509292 320 509298 332
rect 525150 320 525156 332
rect 509292 292 525156 320
rect 509292 280 509298 292
rect 525150 280 525156 292
rect 525208 280 525214 332
rect 526254 280 526260 332
rect 526312 320 526318 332
rect 543458 320 543464 332
rect 526312 292 543464 320
rect 526312 280 526318 292
rect 543458 280 543464 292
rect 543516 280 543522 332
rect 544194 280 544200 332
rect 544252 320 544258 332
rect 550545 323 550603 329
rect 550545 320 550557 323
rect 544252 292 550557 320
rect 544252 280 544258 292
rect 550545 289 550557 292
rect 550591 289 550603 323
rect 550545 283 550603 289
rect 552382 280 552388 332
rect 552440 320 552446 332
rect 555973 323 556031 329
rect 555973 320 555985 323
rect 552440 292 555985 320
rect 552440 280 552446 292
rect 555973 289 555985 292
rect 556019 289 556031 323
rect 557994 320 558000 332
rect 557955 292 558000 320
rect 555973 283 556031 289
rect 557994 280 558000 292
rect 558052 280 558058 332
rect 559006 280 559012 332
rect 559064 320 559070 332
rect 576762 320 576768 332
rect 559064 292 576768 320
rect 559064 280 559070 292
rect 576762 280 576768 292
rect 576820 280 576826 332
rect 484949 255 485007 261
rect 484949 221 484961 255
rect 484995 252 485007 255
rect 492674 252 492680 264
rect 484995 224 492680 252
rect 484995 221 485007 224
rect 484949 215 485007 221
rect 492674 212 492680 224
rect 492732 212 492738 264
rect 494422 212 494428 264
rect 494480 252 494486 264
rect 499942 252 499948 264
rect 494480 224 499948 252
rect 494480 212 494486 224
rect 499942 212 499948 224
rect 500000 212 500006 264
rect 502334 212 502340 264
rect 502392 252 502398 264
rect 518618 252 518624 264
rect 502392 224 518624 252
rect 502392 212 502398 224
rect 518618 212 518624 224
rect 518676 212 518682 264
rect 520366 212 520372 264
rect 520424 252 520430 264
rect 536926 252 536932 264
rect 520424 224 536932 252
rect 520424 212 520430 224
rect 536926 212 536932 224
rect 536984 212 536990 264
rect 538858 212 538864 264
rect 538916 252 538922 264
rect 542265 255 542323 261
rect 542265 252 542277 255
rect 538916 224 542277 252
rect 538916 212 538922 224
rect 542265 221 542277 224
rect 542311 221 542323 255
rect 542265 215 542323 221
rect 542814 212 542820 264
rect 542872 252 542878 264
rect 560662 252 560668 264
rect 542872 224 560668 252
rect 542872 212 542878 224
rect 560662 212 560668 224
rect 560720 212 560726 264
rect 562594 212 562600 264
rect 562652 252 562658 264
rect 581822 252 581828 264
rect 562652 224 581828 252
rect 562652 212 562658 224
rect 581822 212 581828 224
rect 581880 212 581886 264
rect 484854 144 484860 196
rect 484912 184 484918 196
rect 500310 184 500316 196
rect 484912 156 500316 184
rect 484912 144 484918 156
rect 500310 144 500316 156
rect 500368 144 500374 196
rect 501141 187 501199 193
rect 501141 153 501153 187
rect 501187 184 501199 187
rect 503441 187 503499 193
rect 503441 184 503453 187
rect 501187 156 503453 184
rect 501187 153 501199 156
rect 501141 147 501199 153
rect 503441 153 503453 156
rect 503487 153 503499 187
rect 503441 147 503499 153
rect 503530 144 503536 196
rect 503588 184 503594 196
rect 513929 187 513987 193
rect 513929 184 513941 187
rect 503588 156 513941 184
rect 503588 144 503594 156
rect 513929 153 513941 156
rect 513975 153 513987 187
rect 513929 147 513987 153
rect 521562 144 521568 196
rect 521620 184 521626 196
rect 538030 184 538036 196
rect 521620 156 538036 184
rect 521620 144 521626 156
rect 538030 144 538036 156
rect 538088 144 538094 196
rect 539870 144 539876 196
rect 539928 184 539934 196
rect 557166 184 557172 196
rect 539928 156 557172 184
rect 539928 144 539934 156
rect 557166 144 557172 156
rect 557224 144 557230 196
rect 560202 144 560208 196
rect 560260 184 560266 196
rect 578326 184 578332 196
rect 560260 156 578332 184
rect 560260 144 560266 156
rect 578326 144 578332 156
rect 578384 144 578390 196
rect 477460 88 484808 116
rect 485041 119 485099 125
rect 477460 76 477466 88
rect 485041 85 485053 119
rect 485087 116 485099 119
rect 496814 116 496820 128
rect 485087 88 496820 116
rect 485087 85 485099 88
rect 485041 79 485099 85
rect 496814 76 496820 88
rect 496872 76 496878 128
rect 500126 76 500132 128
rect 500184 116 500190 128
rect 512549 119 512607 125
rect 512549 116 512561 119
rect 500184 88 512561 116
rect 500184 76 500190 88
rect 512549 85 512561 88
rect 512595 85 512607 119
rect 512549 79 512607 85
rect 515582 76 515588 128
rect 515640 116 515646 128
rect 532326 116 532332 128
rect 515640 88 532332 116
rect 515640 76 515646 88
rect 532326 76 532332 88
rect 532384 76 532390 128
rect 545666 116 545672 128
rect 532666 88 545672 116
rect 399996 20 408494 48
rect 399996 8 400002 20
rect 411530 8 411536 60
rect 411588 48 411594 60
rect 422481 51 422539 57
rect 422481 48 422493 51
rect 411588 20 422493 48
rect 411588 8 411594 20
rect 422481 17 422493 20
rect 422527 17 422539 51
rect 422481 11 422539 17
rect 429470 8 429476 60
rect 429528 48 429534 60
rect 432693 51 432751 57
rect 432693 48 432705 51
rect 429528 20 432705 48
rect 429528 8 429534 20
rect 432693 17 432705 20
rect 432739 17 432751 51
rect 432693 11 432751 17
rect 433058 8 433064 60
rect 433116 48 433122 60
rect 438397 51 438455 57
rect 438397 48 438409 51
rect 433116 20 438409 48
rect 433116 8 433122 20
rect 438397 17 438409 20
rect 438443 17 438455 51
rect 438397 11 438455 17
rect 439866 8 439872 60
rect 439924 48 439930 60
rect 453482 48 453488 60
rect 439924 20 453488 48
rect 439924 8 439930 20
rect 453482 8 453488 20
rect 453540 8 453546 60
rect 455322 8 455328 60
rect 455380 48 455386 60
rect 469582 48 469588 60
rect 455380 20 469588 48
rect 455380 8 455386 20
rect 469582 8 469588 20
rect 469640 8 469646 60
rect 470873 51 470931 57
rect 470873 17 470885 51
rect 470919 48 470931 51
rect 477862 48 477868 60
rect 470919 20 477868 48
rect 470919 17 470931 20
rect 470873 11 470931 17
rect 477862 8 477868 20
rect 477920 8 477926 60
rect 478506 8 478512 60
rect 478564 48 478570 60
rect 490282 48 490288 60
rect 478564 20 490288 48
rect 478564 8 478570 20
rect 490282 8 490288 20
rect 490340 8 490346 60
rect 496722 8 496728 60
rect 496780 48 496786 60
rect 501141 51 501199 57
rect 501141 48 501153 51
rect 496780 20 501153 48
rect 496780 8 496786 20
rect 501141 17 501153 20
rect 501187 17 501199 51
rect 501141 11 501199 17
rect 501230 8 501236 60
rect 501288 48 501294 60
rect 505189 51 505247 57
rect 505189 48 505201 51
rect 501288 20 505201 48
rect 501288 8 501294 20
rect 505189 17 505201 20
rect 505235 17 505247 51
rect 505189 11 505247 17
rect 505738 8 505744 60
rect 505796 48 505802 60
rect 521654 48 521660 60
rect 505796 20 521660 48
rect 505796 8 505802 20
rect 521654 8 521660 20
rect 521712 8 521718 60
rect 528462 8 528468 60
rect 528520 48 528526 60
rect 532666 48 532694 88
rect 545666 76 545672 88
rect 545724 76 545730 128
rect 546494 76 546500 128
rect 546552 116 546558 128
rect 564618 116 564624 128
rect 546552 88 564624 116
rect 546552 76 546558 88
rect 564618 76 564624 88
rect 564676 76 564682 128
rect 528520 20 532694 48
rect 528520 8 528526 20
rect 545114 8 545120 60
rect 545172 48 545178 60
rect 563054 48 563060 60
rect 545172 20 563060 48
rect 545172 8 545178 20
rect 563054 8 563060 20
rect 563112 8 563118 60
<< via1 >>
rect 271788 703808 271840 703860
rect 364708 703808 364760 703860
rect 235448 703740 235500 703792
rect 300860 703740 300912 703792
rect 257252 703672 257304 703724
rect 394700 703672 394752 703724
rect 242440 703604 242492 703656
rect 400864 703604 400916 703656
rect 170496 703536 170548 703588
rect 315488 703536 315540 703588
rect 227628 703468 227680 703520
rect 468484 703468 468536 703520
rect 105452 703400 105504 703452
rect 330300 703400 330352 703452
rect 1492 703332 1544 703384
rect 359740 703332 359792 703384
rect 213000 703264 213052 703316
rect 576308 703264 576360 703316
rect 1584 703196 1636 703248
rect 374460 703196 374512 703248
rect 198280 703128 198332 703180
rect 575020 703128 575072 703180
rect 1676 703060 1728 703112
rect 389180 703060 389232 703112
rect 183376 702992 183428 703044
rect 573640 702992 573692 703044
rect 756 702924 808 702976
rect 394148 702924 394200 702976
rect 1860 702856 1912 702908
rect 403900 702856 403952 702908
rect 2504 702788 2556 702840
rect 462872 702788 462924 702840
rect 388 702720 440 702772
rect 492680 702720 492732 702772
rect 204 702652 256 702704
rect 507124 702652 507176 702704
rect 41052 702584 41104 702636
rect 578884 702584 578936 702636
rect 2044 702516 2096 702568
rect 551284 702516 551336 702568
rect 21456 702448 21508 702500
rect 576124 702448 576176 702500
rect 70124 702380 70176 702432
rect 573456 702380 573508 702432
rect 237104 702312 237156 702364
rect 291844 702312 291896 702364
rect 134432 702244 134484 702296
rect 266360 702244 266412 702296
rect 277400 702244 277452 702296
rect 428464 702244 428516 702296
rect 144276 702176 144328 702228
rect 324320 702176 324372 702228
rect 100024 702108 100076 702160
rect 311992 702108 312044 702160
rect 119712 702040 119764 702092
rect 340144 702040 340196 702092
rect 55772 701972 55824 702024
rect 305000 701972 305052 702024
rect 338028 701972 338080 702024
rect 482560 701972 482612 702024
rect 6644 701904 6696 701956
rect 259368 701904 259420 701956
rect 280896 701904 280948 701956
rect 467840 701904 467892 701956
rect 154028 701836 154080 701888
rect 565360 701836 565412 701888
rect 163872 701768 163924 701820
rect 577596 701768 577648 701820
rect 148968 701700 149020 701752
rect 574928 701700 574980 701752
rect 572 701632 624 701684
rect 443276 701632 443328 701684
rect 114284 701564 114336 701616
rect 574836 701564 574888 701616
rect 4436 701496 4488 701548
rect 472716 701496 472768 701548
rect 90180 701428 90232 701480
rect 566556 701428 566608 701480
rect 2228 701360 2280 701412
rect 487436 701360 487488 701412
rect 85304 701292 85356 701344
rect 570696 701292 570748 701344
rect 75460 701224 75512 701276
rect 570604 701224 570656 701276
rect 296 701156 348 701208
rect 497280 701156 497332 701208
rect 1308 701088 1360 701140
rect 502340 701088 502392 701140
rect 556896 701088 556948 701140
rect 564440 701088 564492 701140
rect 267004 701020 267056 701072
rect 278596 701020 278648 701072
rect 292488 701020 292540 701072
rect 295892 701020 295944 701072
rect 311900 701020 311952 701072
rect 364616 701020 364668 701072
rect 468576 701020 468628 701072
rect 512000 701020 512052 701072
rect 267648 700952 267700 701004
rect 291384 700952 291436 701004
rect 291844 700952 291896 701004
rect 543464 700952 543516 701004
rect 252284 700884 252336 700936
rect 478512 700884 478564 700936
rect 89168 700816 89220 700868
rect 340052 700816 340104 700868
rect 340144 700816 340196 700868
rect 580632 700816 580684 700868
rect 3424 700748 3476 700800
rect 262864 700748 262916 700800
rect 281356 700748 281408 700800
rect 348792 700748 348844 700800
rect 468484 700748 468536 700800
rect 559656 700748 559708 700800
rect 72976 700680 73028 700732
rect 335360 700680 335412 700732
rect 336648 700680 336700 700732
rect 580356 700680 580408 700732
rect 276848 700612 276900 700664
rect 332508 700612 332560 700664
rect 3976 700544 4028 700596
rect 280896 700544 280948 700596
rect 283840 700544 283892 700596
rect 292488 700544 292540 700596
rect 298100 700544 298152 700596
rect 300124 700544 300176 700596
rect 305000 700544 305052 700596
rect 580448 700544 580500 700596
rect 232688 700476 232740 700528
rect 527180 700476 527232 700528
rect 40500 700408 40552 700460
rect 345204 700408 345256 700460
rect 400864 700408 400916 700460
rect 494796 700408 494848 700460
rect 24308 700340 24360 700392
rect 354956 700340 355008 700392
rect 394700 700340 394752 700392
rect 429844 700340 429896 700392
rect 8116 700272 8168 700324
rect 349896 700272 349948 700324
rect 247408 700204 247460 700256
rect 462320 700204 462372 700256
rect 137836 700136 137888 700188
rect 320778 700136 320830 700188
rect 324320 700136 324372 700188
rect 580816 700136 580868 700188
rect 154120 700068 154172 700120
rect 325654 700068 325706 700120
rect 262128 700000 262180 700052
rect 397460 700000 397512 700052
rect 3332 699932 3384 699984
rect 277308 699932 277360 699984
rect 278596 699932 278648 699984
rect 413652 699932 413704 699984
rect 202696 699864 202748 699916
rect 305736 699864 305788 699916
rect 311992 699864 312044 699916
rect 580540 699864 580592 699916
rect 218980 699796 219032 699848
rect 310612 699796 310664 699848
rect 4252 699728 4304 699780
rect 369768 699728 369820 699780
rect 3792 699660 3844 699712
rect 384304 699660 384356 699712
rect 3148 699592 3200 699644
rect 311900 699592 311952 699644
rect 266360 699524 266412 699576
rect 580724 699524 580776 699576
rect 3884 699456 3936 699508
rect 338028 699456 338080 699508
rect 379520 699499 379572 699508
rect 379520 699465 379529 699499
rect 379529 699465 379563 699499
rect 379563 699465 379572 699499
rect 379520 699456 379572 699465
rect 438308 699499 438360 699508
rect 438308 699465 438317 699499
rect 438317 699465 438351 699499
rect 438351 699465 438360 699499
rect 438308 699456 438360 699465
rect 453028 699499 453080 699508
rect 453028 699465 453037 699499
rect 453037 699465 453071 699499
rect 453071 699465 453080 699499
rect 453028 699456 453080 699465
rect 521844 699499 521896 699508
rect 521844 699465 521853 699499
rect 521853 699465 521887 699499
rect 521887 699465 521896 699499
rect 521844 699456 521896 699465
rect 208124 699388 208176 699440
rect 222844 699388 222896 699440
rect 572168 699388 572220 699440
rect 26148 699363 26200 699372
rect 26148 699329 26157 699363
rect 26157 699329 26191 699363
rect 26191 699329 26200 699363
rect 26148 699320 26200 699329
rect 35992 699363 36044 699372
rect 35992 699329 36001 699363
rect 36001 699329 36035 699363
rect 36035 699329 36044 699363
rect 35992 699320 36044 699329
rect 50896 699363 50948 699372
rect 50896 699329 50905 699363
rect 50905 699329 50939 699363
rect 50939 699329 50948 699363
rect 50896 699320 50948 699329
rect 95148 699363 95200 699372
rect 95148 699329 95157 699363
rect 95157 699329 95191 699363
rect 95191 699329 95200 699363
rect 95148 699320 95200 699329
rect 109868 699363 109920 699372
rect 109868 699329 109877 699363
rect 109877 699329 109911 699363
rect 109911 699329 109920 699363
rect 109868 699320 109920 699329
rect 124588 699363 124640 699372
rect 124588 699329 124597 699363
rect 124597 699329 124631 699363
rect 124631 699329 124640 699363
rect 124588 699320 124640 699329
rect 129464 699363 129516 699372
rect 129464 699329 129473 699363
rect 129473 699329 129507 699363
rect 129507 699329 129516 699363
rect 129464 699320 129516 699329
rect 139308 699363 139360 699372
rect 139308 699329 139317 699363
rect 139317 699329 139351 699363
rect 139351 699329 139360 699363
rect 139308 699320 139360 699329
rect 158812 699363 158864 699372
rect 158812 699329 158821 699363
rect 158821 699329 158855 699363
rect 158855 699329 158864 699363
rect 158812 699320 158864 699329
rect 168840 699363 168892 699372
rect 168840 699329 168849 699363
rect 168849 699329 168883 699363
rect 168883 699329 168892 699363
rect 168840 699320 168892 699329
rect 173716 699363 173768 699372
rect 173716 699329 173725 699363
rect 173725 699329 173759 699363
rect 173759 699329 173768 699363
rect 173716 699320 173768 699329
rect 178592 699363 178644 699372
rect 178592 699329 178601 699363
rect 178601 699329 178635 699363
rect 178635 699329 178644 699363
rect 178592 699320 178644 699329
rect 188436 699363 188488 699372
rect 188436 699329 188445 699363
rect 188445 699329 188479 699363
rect 188479 699329 188488 699363
rect 188436 699320 188488 699329
rect 193220 699320 193272 699372
rect 202972 699320 203024 699372
rect 563704 699320 563756 699372
rect 570880 699252 570932 699304
rect 567844 699184 567896 699236
rect 848 699116 900 699168
rect 576216 699048 576268 699100
rect 569592 698980 569644 699032
rect 573548 698912 573600 698964
rect 569500 698844 569552 698896
rect 572076 698776 572128 698828
rect 480 698708 532 698760
rect 566740 698640 566792 698692
rect 578976 698572 579028 698624
rect 570788 698504 570840 698556
rect 2596 698436 2648 698488
rect 569408 698368 569460 698420
rect 565176 698300 565228 698352
rect 112 697756 164 697808
rect 573364 697688 573416 697740
rect 574744 697620 574796 697672
rect 569224 697552 569276 697604
rect 572168 684428 572220 684480
rect 580172 684428 580224 684480
rect 576308 671984 576360 672036
rect 580172 671984 580224 672036
rect 563704 644376 563756 644428
rect 580172 644376 580224 644428
rect 570880 632000 570932 632052
rect 580172 632000 580224 632052
rect 575020 618196 575072 618248
rect 580172 618196 580224 618248
rect 576216 591948 576268 592000
rect 579988 591948 580040 592000
rect 567844 578144 567896 578196
rect 579804 578144 579856 578196
rect 3792 565836 3844 565888
rect 4344 565836 4396 565888
rect 573640 564340 573692 564392
rect 580172 564340 580224 564392
rect 573548 538160 573600 538212
rect 580172 538160 580224 538212
rect 569592 525716 569644 525768
rect 580172 525716 580224 525768
rect 569500 511912 569552 511964
rect 580172 511912 580224 511964
rect 3148 502256 3200 502308
rect 4436 502256 4488 502308
rect 572076 485732 572128 485784
rect 580172 485732 580224 485784
rect 577596 471928 577648 471980
rect 580908 471928 580960 471980
rect 565360 458124 565412 458176
rect 580172 458124 580224 458176
rect 574928 419432 574980 419484
rect 580172 419432 580224 419484
rect 566740 379448 566792 379500
rect 580172 379448 580224 379500
rect 570788 353200 570840 353252
rect 580172 353200 580224 353252
rect 574836 325592 574888 325644
rect 579988 325592 580040 325644
rect 569408 299412 569460 299464
rect 580172 299412 580224 299464
rect 571984 259360 572036 259412
rect 580172 259360 580224 259412
rect 1308 249704 1360 249756
rect 2780 249704 2832 249756
rect 565176 245556 565228 245608
rect 580172 245556 580224 245608
rect 570696 233180 570748 233232
rect 579620 233180 579672 233232
rect 566556 219376 566608 219428
rect 580172 219376 580224 219428
rect 566648 206932 566700 206984
rect 580172 206932 580224 206984
rect 573456 193128 573508 193180
rect 580172 193128 580224 193180
rect 570604 179324 570656 179376
rect 580172 179324 580224 179376
rect 565268 166948 565320 167000
rect 580172 166948 580224 167000
rect 569316 139340 569368 139392
rect 580172 139340 580224 139392
rect 573364 126896 573416 126948
rect 580172 126896 580224 126948
rect 577504 100648 577556 100700
rect 579804 100648 579856 100700
rect 574744 86912 574796 86964
rect 579620 86912 579672 86964
rect 569224 73108 569276 73160
rect 580172 73108 580224 73160
rect 576124 46860 576176 46912
rect 580172 46860 580224 46912
rect 566464 33056 566516 33108
rect 580172 33056 580224 33108
rect 565084 20612 565136 20664
rect 580172 20612 580224 20664
rect 563612 3136 563664 3188
rect 569132 3136 569184 3188
rect 565912 3068 565964 3120
rect 571524 3068 571576 3120
rect 563704 3000 563756 3052
rect 583392 3000 583444 3052
rect 563520 2864 563572 2916
rect 572720 2864 572772 2916
rect 569868 2796 569920 2848
rect 576308 2796 576360 2848
rect 3056 1300 3108 1352
rect 564440 1300 564492 1352
rect 566832 1164 566884 1216
rect 581000 1096 581052 1148
rect 1676 620 1728 672
rect 5356 620 5408 672
rect 6460 620 6512 672
rect 10048 620 10100 672
rect 572 552 624 604
rect 4344 552 4396 604
rect 5264 552 5316 604
rect 8852 552 8904 604
rect 7472 527 7524 536
rect 7472 493 7481 527
rect 7481 493 7515 527
rect 7515 493 7524 527
rect 7472 484 7524 493
rect 8576 484 8628 536
rect 11152 552 11204 604
rect 11520 620 11572 672
rect 19432 620 19484 672
rect 22376 620 22428 672
rect 12348 552 12400 604
rect 15568 552 15620 604
rect 21824 552 21876 604
rect 24860 620 24912 672
rect 25320 620 25372 672
rect 28080 620 28132 672
rect 28724 620 28776 672
rect 29184 620 29236 672
rect 31300 620 31352 672
rect 33784 620 33836 672
rect 34796 620 34848 672
rect 37280 620 37332 672
rect 38384 620 38436 672
rect 23020 552 23072 604
rect 25780 552 25832 604
rect 28816 552 28868 604
rect 3240 416 3292 468
rect 6644 416 6696 468
rect 12624 484 12676 536
rect 13360 484 13412 536
rect 16672 484 16724 536
rect 17408 484 17460 536
rect 20076 484 20128 536
rect 30104 552 30156 604
rect 32588 552 32640 604
rect 33600 552 33652 604
rect 36084 552 36136 604
rect 37188 552 37240 604
rect 40684 620 40736 672
rect 42800 620 42852 672
rect 46664 620 46716 672
rect 48504 620 48556 672
rect 48964 620 49016 672
rect 50804 620 50856 672
rect 53748 620 53800 672
rect 55404 620 55456 672
rect 64328 620 64380 672
rect 65616 620 65668 672
rect 66720 620 66772 672
rect 68008 620 68060 672
rect 69112 620 69164 672
rect 70584 620 70636 672
rect 133236 620 133288 672
rect 134156 620 134208 672
rect 136180 620 136232 672
rect 137652 620 137704 672
rect 138756 620 138808 672
rect 140044 620 140096 672
rect 151360 620 151412 672
rect 153016 620 153068 672
rect 153660 620 153712 672
rect 155408 620 155460 672
rect 162768 620 162820 672
rect 164884 620 164936 672
rect 40776 552 40828 604
rect 41880 552 41932 604
rect 43996 552 44048 604
rect 47860 552 47912 604
rect 49608 552 49660 604
rect 50160 552 50212 604
rect 51356 552 51408 604
rect 53012 552 53064 604
rect 54944 552 54996 604
rect 56416 552 56468 604
rect 60832 552 60884 604
rect 62120 552 62172 604
rect 65524 552 65576 604
rect 66812 552 66864 604
rect 70308 552 70360 604
rect 71228 552 71280 604
rect 76196 552 76248 604
rect 76932 552 76984 604
rect 77392 552 77444 604
rect 78036 552 78088 604
rect 78588 552 78640 604
rect 79140 552 79192 604
rect 79692 552 79744 604
rect 80336 552 80388 604
rect 80888 552 80940 604
rect 81440 552 81492 604
rect 82084 552 82136 604
rect 82728 552 82780 604
rect 121828 552 121880 604
rect 122288 552 122340 604
rect 124128 552 124180 604
rect 124680 552 124732 604
rect 125232 552 125284 604
rect 125876 552 125928 604
rect 126428 552 126480 604
rect 126980 552 127032 604
rect 127532 552 127584 604
rect 128176 552 128228 604
rect 128636 552 128688 604
rect 129372 552 129424 604
rect 133880 552 133932 604
rect 135260 552 135312 604
rect 136456 552 136508 604
rect 137560 552 137612 604
rect 138848 552 138900 604
rect 139952 552 140004 604
rect 141240 552 141292 604
rect 144552 552 144604 604
rect 145932 552 145984 604
rect 146852 552 146904 604
rect 148324 552 148376 604
rect 152556 552 152608 604
rect 154212 552 154264 604
rect 154764 552 154816 604
rect 156604 552 156656 604
rect 157064 552 157116 604
rect 158904 552 158956 604
rect 161572 552 161624 604
rect 163688 552 163740 604
rect 31668 484 31720 536
rect 33232 484 33284 536
rect 34980 484 35032 536
rect 14464 416 14516 468
rect 14556 416 14608 468
rect 17868 416 17920 468
rect 24400 416 24452 468
rect 26884 416 26936 468
rect 51908 484 51960 536
rect 63500 484 63552 536
rect 64512 484 64564 536
rect 67732 484 67784 536
rect 69388 484 69440 536
rect 134984 484 135036 536
rect 141056 484 141108 536
rect 142068 484 142120 536
rect 158168 484 158220 536
rect 159732 484 159784 536
rect 39856 416 39908 468
rect 163412 416 163464 468
rect 166080 620 166132 672
rect 167092 620 167144 672
rect 169576 620 169628 672
rect 180892 620 180944 672
rect 183744 620 183796 672
rect 165988 552 166040 604
rect 168380 552 168432 604
rect 170680 552 170732 604
rect 173164 552 173216 604
rect 179788 552 179840 604
rect 182548 552 182600 604
rect 183192 552 183244 604
rect 186136 620 186188 672
rect 191104 620 191156 672
rect 194416 620 194468 672
rect 211620 620 211672 672
rect 215668 620 215720 672
rect 220176 620 220228 672
rect 225328 620 225380 672
rect 226156 620 226208 672
rect 231032 620 231084 672
rect 190000 552 190052 604
rect 193220 552 193272 604
rect 195612 552 195664 604
rect 196808 595 196860 604
rect 196808 561 196817 595
rect 196817 561 196851 595
rect 196851 561 196860 595
rect 196808 552 196860 561
rect 197912 552 197964 604
rect 205732 552 205784 604
rect 209780 552 209832 604
rect 210424 552 210476 604
rect 212172 552 212224 604
rect 214472 595 214524 604
rect 214472 561 214481 595
rect 214481 561 214515 595
rect 214515 561 214524 595
rect 214472 552 214524 561
rect 219992 552 220044 604
rect 220452 552 220504 604
rect 223948 552 224000 604
rect 225052 552 225104 604
rect 186596 484 186648 536
rect 189908 484 189960 536
rect 192300 484 192352 536
rect 187700 416 187752 468
rect 191012 416 191064 468
rect 194048 416 194100 468
rect 208400 484 208452 536
rect 212724 484 212776 536
rect 216588 484 216640 536
rect 219532 484 219584 536
rect 227352 484 227404 536
rect 229836 552 229888 604
rect 229652 484 229704 536
rect 234620 620 234672 672
rect 235448 620 235500 672
rect 237748 620 237800 672
rect 242900 620 242952 672
rect 246764 620 246816 672
rect 247960 620 248012 672
rect 253480 620 253532 672
rect 257252 620 257304 672
rect 258264 620 258316 672
rect 231860 552 231912 604
rect 237012 552 237064 604
rect 238116 552 238168 604
rect 233148 484 233200 536
rect 218428 416 218480 468
rect 222936 416 222988 468
rect 39304 348 39356 400
rect 42156 348 42208 400
rect 42892 348 42944 400
rect 45100 348 45152 400
rect 71320 348 71372 400
rect 72332 348 72384 400
rect 72424 348 72476 400
rect 73528 348 73580 400
rect 73620 348 73672 400
rect 74632 348 74684 400
rect 130936 348 130988 400
rect 131948 348 132000 400
rect 132040 348 132092 400
rect 133144 348 133196 400
rect 160468 348 160520 400
rect 162676 348 162728 400
rect 192944 348 192996 400
rect 217232 348 217284 400
rect 221740 348 221792 400
rect 222476 348 222528 400
rect 234344 416 234396 468
rect 239312 552 239364 604
rect 240508 595 240560 604
rect 240508 561 240517 595
rect 240517 561 240551 595
rect 240551 561 240560 595
rect 240508 552 240560 561
rect 241152 552 241204 604
rect 246028 552 246080 604
rect 249984 552 250036 604
rect 251180 552 251232 604
rect 252376 595 252428 604
rect 252376 561 252385 595
rect 252385 561 252419 595
rect 252419 561 252428 595
rect 252376 552 252428 561
rect 253388 552 253440 604
rect 254584 552 254636 604
rect 260656 620 260708 672
rect 262680 620 262732 672
rect 268844 620 268896 672
rect 269488 620 269540 672
rect 276204 620 276256 672
rect 279240 620 279292 672
rect 279516 663 279568 672
rect 279516 629 279525 663
rect 279525 629 279559 663
rect 279559 629 279568 663
rect 279516 620 279568 629
rect 238852 484 238904 536
rect 243912 484 243964 536
rect 243360 416 243412 468
rect 248972 484 249024 536
rect 244556 416 244608 468
rect 242256 348 242308 400
rect 247316 348 247368 400
rect 245660 280 245712 332
rect 259460 552 259512 604
rect 260472 552 260524 604
rect 266544 552 266596 604
rect 267740 552 267792 604
rect 270040 595 270092 604
rect 270040 561 270049 595
rect 270049 561 270083 595
rect 270083 561 270092 595
rect 270040 552 270092 561
rect 271788 552 271840 604
rect 261576 484 261628 536
rect 268384 484 268436 536
rect 274548 484 274600 536
rect 277492 552 277544 604
rect 284300 620 284352 672
rect 286600 620 286652 672
rect 291108 620 291160 672
rect 298468 620 298520 672
rect 304724 620 304776 672
rect 307668 663 307720 672
rect 307668 629 307677 663
rect 307677 629 307711 663
rect 307711 629 307720 663
rect 307668 620 307720 629
rect 309968 620 310020 672
rect 280712 595 280764 604
rect 280712 561 280721 595
rect 280721 561 280755 595
rect 280755 561 280764 595
rect 280712 552 280764 561
rect 283104 595 283156 604
rect 283104 561 283113 595
rect 283113 561 283147 595
rect 283147 561 283156 595
rect 283104 552 283156 561
rect 285404 552 285456 604
rect 288808 552 288860 604
rect 296076 552 296128 604
rect 278504 484 278556 536
rect 278596 484 278648 536
rect 286416 484 286468 536
rect 293316 484 293368 536
rect 227352 212 227404 264
rect 232044 212 232096 264
rect 233240 212 233292 264
rect 250904 212 250956 264
rect 256884 416 256936 468
rect 257988 416 258040 468
rect 259276 416 259328 468
rect 264980 416 265032 468
rect 266084 416 266136 468
rect 272156 416 272208 468
rect 280436 416 280488 468
rect 287520 416 287572 468
rect 289820 416 289872 468
rect 297272 552 297324 604
rect 300216 552 300268 604
rect 296812 484 296864 536
rect 303988 484 304040 536
rect 307944 552 307996 604
rect 309048 552 309100 604
rect 310244 552 310296 604
rect 311440 552 311492 604
rect 301320 416 301372 468
rect 263140 348 263192 400
rect 270684 348 270736 400
rect 276756 348 276808 400
rect 281540 348 281592 400
rect 287060 348 287112 400
rect 287612 348 287664 400
rect 293868 348 293920 400
rect 294512 348 294564 400
rect 301780 348 301832 400
rect 252008 280 252060 332
rect 257252 280 257304 332
rect 275836 280 275888 332
rect 284116 280 284168 332
rect 291200 280 291252 332
rect 299020 280 299072 332
rect 306932 348 306984 400
rect 302424 280 302476 332
rect 312636 620 312688 672
rect 315948 620 316000 672
rect 319720 663 319772 672
rect 319720 629 319729 663
rect 319729 629 319763 663
rect 319763 629 319772 663
rect 319720 620 319772 629
rect 316224 552 316276 604
rect 320916 620 320968 672
rect 323308 620 323360 672
rect 324412 620 324464 672
rect 312452 484 312504 536
rect 320640 552 320692 604
rect 329196 620 329248 672
rect 335360 620 335412 672
rect 325608 552 325660 604
rect 328000 552 328052 604
rect 332692 552 332744 604
rect 334256 552 334308 604
rect 337476 552 337528 604
rect 338672 595 338724 604
rect 338672 561 338681 595
rect 338681 561 338715 595
rect 338715 561 338724 595
rect 338672 552 338724 561
rect 339868 552 339920 604
rect 340972 552 341024 604
rect 341800 595 341852 604
rect 341800 561 341809 595
rect 341809 561 341843 595
rect 341843 561 341852 595
rect 341800 552 341852 561
rect 342168 595 342220 604
rect 342168 561 342177 595
rect 342177 561 342211 595
rect 342211 561 342220 595
rect 342168 552 342220 561
rect 344560 620 344612 672
rect 347688 620 347740 672
rect 357532 620 357584 672
rect 343364 552 343416 604
rect 343456 552 343508 604
rect 345756 552 345808 604
rect 352840 552 352892 604
rect 317144 484 317196 536
rect 318156 416 318208 468
rect 319536 416 319588 468
rect 330852 484 330904 536
rect 331956 416 332008 468
rect 347688 484 347740 536
rect 354036 552 354088 604
rect 356336 595 356388 604
rect 356336 561 356345 595
rect 356345 561 356379 595
rect 356379 561 356388 595
rect 356336 552 356388 561
rect 356980 552 357032 604
rect 367008 620 367060 672
rect 368204 663 368256 672
rect 368204 629 368213 663
rect 368213 629 368247 663
rect 368247 629 368256 663
rect 368204 620 368256 629
rect 369400 620 369452 672
rect 359280 595 359332 604
rect 359280 561 359289 595
rect 359289 561 359323 595
rect 359323 561 359332 595
rect 359280 552 359332 561
rect 362684 552 362736 604
rect 370412 620 370464 672
rect 372896 663 372948 672
rect 372896 629 372905 663
rect 372905 629 372939 663
rect 372939 629 372948 663
rect 372896 620 372948 629
rect 381176 620 381228 672
rect 382372 620 382424 672
rect 370688 552 370740 604
rect 371608 552 371660 604
rect 382004 552 382056 604
rect 384212 620 384264 672
rect 386512 663 386564 672
rect 386512 629 386521 663
rect 386521 629 386555 663
rect 386555 629 386564 663
rect 386512 620 386564 629
rect 400128 663 400180 672
rect 383568 552 383620 604
rect 385408 552 385460 604
rect 400128 629 400137 663
rect 400137 629 400171 663
rect 400171 629 400180 663
rect 400128 620 400180 629
rect 401324 620 401376 672
rect 402428 620 402480 672
rect 405648 663 405700 672
rect 405648 629 405657 663
rect 405657 629 405691 663
rect 405691 629 405700 663
rect 405648 620 405700 629
rect 407212 620 407264 672
rect 408316 663 408368 672
rect 408316 629 408325 663
rect 408325 629 408359 663
rect 408359 629 408368 663
rect 408316 620 408368 629
rect 388260 595 388312 604
rect 388260 561 388269 595
rect 388269 561 388303 595
rect 388303 561 388312 595
rect 388260 552 388312 561
rect 389456 595 389508 604
rect 389456 561 389465 595
rect 389465 561 389499 595
rect 389499 561 389508 595
rect 389456 552 389508 561
rect 389916 595 389968 604
rect 389916 561 389925 595
rect 389925 561 389959 595
rect 389959 561 389968 595
rect 389916 552 389968 561
rect 391020 552 391072 604
rect 354680 484 354732 536
rect 358544 484 358596 536
rect 360384 484 360436 536
rect 372436 484 372488 536
rect 343180 416 343232 468
rect 349068 416 349120 468
rect 363788 416 363840 468
rect 314752 348 314804 400
rect 313648 280 313700 332
rect 318340 348 318392 400
rect 326620 348 326672 400
rect 327448 348 327500 400
rect 255688 212 255740 264
rect 261944 212 261996 264
rect 263692 212 263744 264
rect 272892 212 272944 264
rect 297916 212 297968 264
rect 305736 212 305788 264
rect 308772 212 308824 264
rect 316408 212 316460 264
rect 16304 76 16356 128
rect 18972 76 19024 128
rect 45744 76 45796 128
rect 47400 76 47452 128
rect 129832 76 129884 128
rect 130292 76 130344 128
rect 155960 76 156012 128
rect 157524 76 157576 128
rect 159364 76 159416 128
rect 161480 76 161532 128
rect 184296 76 184348 128
rect 186964 144 187016 196
rect 228548 144 228600 196
rect 236552 144 236604 196
rect 241428 144 241480 196
rect 274088 144 274140 196
rect 282920 144 282972 196
rect 290004 144 290056 196
rect 292212 144 292264 196
rect 299388 144 299440 196
rect 321560 280 321612 332
rect 330116 280 330168 332
rect 333152 348 333204 400
rect 340604 348 340656 400
rect 350172 348 350224 400
rect 351276 391 351328 400
rect 351276 357 351285 391
rect 351285 357 351319 391
rect 351319 357 351328 391
rect 351276 348 351328 357
rect 352472 348 352524 400
rect 355876 348 355928 400
rect 365996 348 366048 400
rect 336464 280 336516 332
rect 337200 280 337252 332
rect 346676 280 346728 332
rect 321836 144 321888 196
rect 324044 144 324096 196
rect 328552 212 328604 264
rect 346768 212 346820 264
rect 364800 280 364852 332
rect 375104 416 375156 468
rect 379704 416 379756 468
rect 377404 348 377456 400
rect 378600 348 378652 400
rect 383108 416 383160 468
rect 394424 484 394476 536
rect 396264 527 396316 536
rect 396264 493 396273 527
rect 396273 493 396307 527
rect 396307 493 396316 527
rect 396264 484 396316 493
rect 396540 552 396592 604
rect 397736 595 397788 604
rect 397736 561 397745 595
rect 397745 561 397779 595
rect 397779 561 397788 595
rect 397736 552 397788 561
rect 398840 552 398892 604
rect 410800 620 410852 672
rect 414296 620 414348 672
rect 414940 663 414992 672
rect 414940 629 414949 663
rect 414949 629 414983 663
rect 414983 629 414992 663
rect 414940 620 414992 629
rect 415216 663 415268 672
rect 415216 629 415225 663
rect 415225 629 415259 663
rect 415259 629 415268 663
rect 415216 620 415268 629
rect 416044 620 416096 672
rect 424968 620 425020 672
rect 426992 620 427044 672
rect 428464 663 428516 672
rect 402704 484 402756 536
rect 404544 484 404596 536
rect 416688 552 416740 604
rect 423772 552 423824 604
rect 426164 552 426216 604
rect 427268 595 427320 604
rect 427268 561 427277 595
rect 427277 561 427311 595
rect 427311 561 427320 595
rect 427268 552 427320 561
rect 428004 595 428056 604
rect 428004 561 428013 595
rect 428013 561 428047 595
rect 428047 561 428056 595
rect 428004 552 428056 561
rect 428464 629 428473 663
rect 428473 629 428507 663
rect 428507 629 428516 663
rect 428464 620 428516 629
rect 431868 663 431920 672
rect 431868 629 431877 663
rect 431877 629 431911 663
rect 431911 629 431920 663
rect 431868 620 431920 629
rect 432052 595 432104 604
rect 432052 561 432061 595
rect 432061 561 432095 595
rect 432095 561 432104 595
rect 432052 552 432104 561
rect 434444 620 434496 672
rect 434720 620 434772 672
rect 435364 620 435416 672
rect 435548 663 435600 672
rect 435548 629 435557 663
rect 435557 629 435591 663
rect 435591 629 435600 663
rect 435548 620 435600 629
rect 437480 620 437532 672
rect 449624 620 449676 672
rect 451280 663 451332 672
rect 451280 629 451289 663
rect 451289 629 451323 663
rect 451323 629 451332 663
rect 451280 620 451332 629
rect 454224 663 454276 672
rect 454224 629 454233 663
rect 454233 629 454267 663
rect 454267 629 454276 663
rect 454224 620 454276 629
rect 455696 663 455748 672
rect 455696 629 455705 663
rect 455705 629 455739 663
rect 455739 629 455748 663
rect 455696 620 455748 629
rect 456800 620 456852 672
rect 440332 552 440384 604
rect 441528 595 441580 604
rect 441528 561 441537 595
rect 441537 561 441571 595
rect 441571 561 441580 595
rect 441528 552 441580 561
rect 442632 595 442684 604
rect 442632 561 442641 595
rect 442641 561 442675 595
rect 442675 561 442684 595
rect 442632 552 442684 561
rect 443276 595 443328 604
rect 443276 561 443285 595
rect 443285 561 443319 595
rect 443319 561 443328 595
rect 443276 552 443328 561
rect 445024 595 445076 604
rect 445024 561 445033 595
rect 445033 561 445067 595
rect 445067 561 445076 595
rect 445024 552 445076 561
rect 446220 595 446272 604
rect 446220 561 446229 595
rect 446229 561 446263 595
rect 446263 561 446272 595
rect 446220 552 446272 561
rect 446680 595 446732 604
rect 446680 561 446689 595
rect 446689 561 446723 595
rect 446723 561 446732 595
rect 446680 552 446732 561
rect 447416 595 447468 604
rect 447416 561 447425 595
rect 447425 561 447459 595
rect 447459 561 447468 595
rect 447416 552 447468 561
rect 409236 484 409288 536
rect 421012 484 421064 536
rect 422392 527 422444 536
rect 422392 493 422401 527
rect 422401 493 422435 527
rect 422435 493 422444 527
rect 422392 484 422444 493
rect 430672 484 430724 536
rect 388812 416 388864 468
rect 351276 212 351328 264
rect 325148 144 325200 196
rect 333612 144 333664 196
rect 338304 144 338356 196
rect 185492 76 185544 128
rect 188252 76 188304 128
rect 213828 76 213880 128
rect 217876 76 217928 128
rect 329748 76 329800 128
rect 339500 76 339552 128
rect 345572 144 345624 196
rect 354956 144 355008 196
rect 357164 144 357216 196
rect 358084 212 358136 264
rect 369032 280 369084 332
rect 379796 280 379848 332
rect 380808 280 380860 332
rect 391572 280 391624 332
rect 373908 212 373960 264
rect 377404 212 377456 264
rect 395620 416 395672 468
rect 393228 391 393280 400
rect 393228 357 393237 391
rect 393237 357 393271 391
rect 393271 357 393280 391
rect 393228 348 393280 357
rect 395528 391 395580 400
rect 395528 357 395537 391
rect 395537 357 395571 391
rect 395571 357 395580 391
rect 395528 348 395580 357
rect 403440 416 403492 468
rect 415308 416 415360 468
rect 417148 416 417200 468
rect 429476 416 429528 468
rect 406936 348 406988 400
rect 418804 348 418856 400
rect 420552 348 420604 400
rect 432972 416 433024 468
rect 438768 484 438820 536
rect 454500 595 454552 604
rect 454500 561 454509 595
rect 454509 561 454543 595
rect 454543 561 454552 595
rect 454500 552 454552 561
rect 460388 552 460440 604
rect 461952 620 462004 672
rect 463148 663 463200 672
rect 463148 629 463157 663
rect 463157 629 463191 663
rect 463191 629 463200 663
rect 463148 620 463200 629
rect 463608 620 463660 672
rect 464896 663 464948 672
rect 464896 629 464905 663
rect 464905 629 464939 663
rect 464939 629 464948 663
rect 464896 620 464948 629
rect 468392 663 468444 672
rect 461768 552 461820 604
rect 467472 552 467524 604
rect 468392 629 468401 663
rect 468401 629 468435 663
rect 468435 629 468444 663
rect 468392 620 468444 629
rect 469220 663 469272 672
rect 469220 629 469229 663
rect 469229 629 469263 663
rect 469263 629 469272 663
rect 469220 620 469272 629
rect 471060 620 471112 672
rect 471704 620 471756 672
rect 474004 663 474056 672
rect 474004 629 474013 663
rect 474013 629 474047 663
rect 474047 629 474056 663
rect 474004 620 474056 629
rect 476764 663 476816 672
rect 476764 629 476773 663
rect 476773 629 476807 663
rect 476807 629 476816 663
rect 476764 620 476816 629
rect 476948 663 477000 672
rect 476948 629 476957 663
rect 476957 629 476991 663
rect 476991 629 477000 663
rect 476948 620 477000 629
rect 473452 552 473504 604
rect 475108 552 475160 604
rect 485136 620 485188 672
rect 486608 663 486660 672
rect 486608 629 486617 663
rect 486617 629 486651 663
rect 486651 629 486660 663
rect 486608 620 486660 629
rect 487804 620 487856 672
rect 488540 620 488592 672
rect 479616 595 479668 604
rect 479616 561 479625 595
rect 479625 561 479659 595
rect 479659 561 479668 595
rect 479616 552 479668 561
rect 483112 595 483164 604
rect 483112 561 483121 595
rect 483121 561 483155 595
rect 483155 561 483164 595
rect 483112 552 483164 561
rect 483756 595 483808 604
rect 483756 561 483765 595
rect 483765 561 483799 595
rect 483799 561 483808 595
rect 483756 552 483808 561
rect 484032 595 484084 604
rect 484032 561 484041 595
rect 484041 561 484075 595
rect 484075 561 484084 595
rect 484032 552 484084 561
rect 485228 552 485280 604
rect 486332 552 486384 604
rect 448244 527 448296 536
rect 448244 493 448253 527
rect 448253 493 448287 527
rect 448287 493 448296 527
rect 448244 484 448296 493
rect 450636 484 450688 536
rect 443644 416 443696 468
rect 444472 416 444524 468
rect 458272 484 458324 536
rect 459008 484 459060 536
rect 467196 527 467248 536
rect 467196 493 467205 527
rect 467205 493 467239 527
rect 467239 493 467248 527
rect 467196 484 467248 493
rect 468300 484 468352 536
rect 469496 484 469548 536
rect 480812 484 480864 536
rect 457168 459 457220 468
rect 457168 425 457177 459
rect 457177 425 457211 459
rect 457211 425 457220 459
rect 457168 416 457220 425
rect 457904 416 457956 468
rect 471980 416 472032 468
rect 472808 416 472860 468
rect 360844 144 360896 196
rect 366732 144 366784 196
rect 367836 144 367888 196
rect 44088 8 44140 60
rect 46204 8 46256 60
rect 215024 8 215076 60
rect 219440 8 219492 60
rect 256884 8 256936 60
rect 262772 8 262824 60
rect 264888 8 264940 60
rect 271052 8 271104 60
rect 293408 8 293460 60
rect 300492 8 300544 60
rect 303620 8 303672 60
rect 311072 8 311124 60
rect 322848 8 322900 60
rect 331220 8 331272 60
rect 347688 76 347740 128
rect 349436 76 349488 128
rect 353576 76 353628 128
rect 363696 76 363748 128
rect 373816 144 373868 196
rect 384580 144 384632 196
rect 393964 144 394016 196
rect 397460 144 397512 196
rect 409420 280 409472 332
rect 410340 280 410392 332
rect 422760 280 422812 332
rect 423496 280 423548 332
rect 424692 280 424744 332
rect 437572 348 437624 400
rect 442172 348 442224 400
rect 460204 348 460256 400
rect 474372 348 474424 400
rect 479524 391 479576 400
rect 479524 357 479533 391
rect 479533 357 479567 391
rect 479567 357 479576 391
rect 479524 348 479576 357
rect 481456 348 481508 400
rect 487528 552 487580 604
rect 492128 663 492180 672
rect 492128 629 492137 663
rect 492137 629 492171 663
rect 492171 629 492180 663
rect 492128 620 492180 629
rect 493324 663 493376 672
rect 493324 629 493333 663
rect 493333 629 493367 663
rect 493367 629 493376 663
rect 493324 620 493376 629
rect 497832 663 497884 672
rect 497832 629 497841 663
rect 497841 629 497875 663
rect 497875 629 497884 663
rect 497832 620 497884 629
rect 498200 620 498252 672
rect 498936 620 498988 672
rect 504180 620 504232 672
rect 504640 663 504692 672
rect 504640 629 504649 663
rect 504649 629 504683 663
rect 504683 629 504692 663
rect 504640 620 504692 629
rect 506940 620 506992 672
rect 507952 663 508004 672
rect 507952 629 507961 663
rect 507961 629 507995 663
rect 507995 629 508004 663
rect 508596 663 508648 672
rect 507952 620 508004 629
rect 508596 629 508605 663
rect 508605 629 508639 663
rect 508639 629 508648 663
rect 508596 620 508648 629
rect 509884 663 509936 672
rect 509884 629 509893 663
rect 509893 629 509927 663
rect 509927 629 509936 663
rect 509884 620 509936 629
rect 492864 552 492916 604
rect 493508 552 493560 604
rect 499396 595 499448 604
rect 499396 561 499405 595
rect 499405 561 499439 595
rect 499439 561 499448 595
rect 499396 552 499448 561
rect 501788 552 501840 604
rect 502984 595 503036 604
rect 502984 561 502993 595
rect 502993 561 503027 595
rect 503027 561 503036 595
rect 502984 552 503036 561
rect 513288 620 513340 672
rect 513564 663 513616 672
rect 513564 629 513573 663
rect 513573 629 513607 663
rect 513607 629 513616 663
rect 513564 620 513616 629
rect 514668 663 514720 672
rect 514668 629 514677 663
rect 514677 629 514711 663
rect 514711 629 514720 663
rect 514668 620 514720 629
rect 514760 663 514812 672
rect 514760 629 514769 663
rect 514769 629 514803 663
rect 514803 629 514812 663
rect 518256 663 518308 672
rect 514760 620 514812 629
rect 518256 629 518265 663
rect 518265 629 518299 663
rect 518299 629 518308 663
rect 518256 620 518308 629
rect 519544 620 519596 672
rect 520096 620 520148 672
rect 520740 663 520792 672
rect 520740 629 520749 663
rect 520749 629 520783 663
rect 520783 629 520792 663
rect 520740 620 520792 629
rect 522856 663 522908 672
rect 522856 629 522865 663
rect 522865 629 522899 663
rect 522899 629 522908 663
rect 522856 620 522908 629
rect 523040 663 523092 672
rect 523040 629 523049 663
rect 523049 629 523083 663
rect 523083 629 523092 663
rect 523040 620 523092 629
rect 523960 663 524012 672
rect 523960 629 523969 663
rect 523969 629 524003 663
rect 524003 629 524012 663
rect 523960 620 524012 629
rect 524236 663 524288 672
rect 524236 629 524245 663
rect 524245 629 524279 663
rect 524279 629 524288 663
rect 524236 620 524288 629
rect 525064 620 525116 672
rect 531872 663 531924 672
rect 531872 629 531881 663
rect 531881 629 531915 663
rect 531915 629 531924 663
rect 531872 620 531924 629
rect 535828 620 535880 672
rect 538772 663 538824 672
rect 538772 629 538781 663
rect 538781 629 538815 663
rect 538815 629 538824 663
rect 538772 620 538824 629
rect 511264 552 511316 604
rect 512460 552 512512 604
rect 515956 552 516008 604
rect 517060 552 517112 604
rect 529940 552 529992 604
rect 530124 595 530176 604
rect 530124 561 530133 595
rect 530133 561 530167 595
rect 530167 561 530176 595
rect 530124 552 530176 561
rect 531320 595 531372 604
rect 531320 561 531329 595
rect 531329 561 531363 595
rect 531363 561 531372 595
rect 531320 552 531372 561
rect 534540 595 534592 604
rect 534540 561 534549 595
rect 534549 561 534583 595
rect 534583 561 534592 595
rect 534540 552 534592 561
rect 489000 459 489052 468
rect 489000 425 489009 459
rect 489009 425 489043 459
rect 489043 425 489052 459
rect 489000 416 489052 425
rect 491484 416 491536 468
rect 495532 416 495584 468
rect 445576 280 445628 332
rect 401140 212 401192 264
rect 408132 212 408184 264
rect 419908 212 419960 264
rect 421748 212 421800 264
rect 425796 212 425848 264
rect 438768 212 438820 264
rect 378692 76 378744 128
rect 379520 76 379572 128
rect 390284 76 390336 128
rect 393320 76 393372 128
rect 404544 76 404596 128
rect 412916 144 412968 196
rect 413744 144 413796 196
rect 436468 144 436520 196
rect 449992 280 450044 332
rect 452292 323 452344 332
rect 452292 289 452301 323
rect 452301 289 452335 323
rect 452335 289 452344 323
rect 452292 280 452344 289
rect 452384 280 452436 332
rect 465908 280 465960 332
rect 470600 280 470652 332
rect 489736 348 489788 400
rect 505100 348 505152 400
rect 509792 348 509844 400
rect 510988 348 511040 400
rect 519360 484 519412 536
rect 520096 484 520148 536
rect 526444 527 526496 536
rect 526444 493 526453 527
rect 526453 493 526487 527
rect 526487 493 526496 527
rect 526444 484 526496 493
rect 527180 484 527232 536
rect 512184 416 512236 468
rect 528836 416 528888 468
rect 539140 620 539192 672
rect 543740 620 543792 672
rect 546684 620 546736 672
rect 548340 620 548392 672
rect 548984 620 549036 672
rect 563520 1028 563572 1080
rect 569868 960 569920 1012
rect 563612 892 563664 944
rect 551192 620 551244 672
rect 565912 824 565964 876
rect 565636 756 565688 808
rect 565820 756 565872 808
rect 568028 756 568080 808
rect 570328 688 570380 740
rect 553308 620 553360 672
rect 554596 663 554648 672
rect 554596 629 554605 663
rect 554605 629 554639 663
rect 554639 629 554648 663
rect 554596 620 554648 629
rect 555884 663 555936 672
rect 555884 629 555893 663
rect 555893 629 555927 663
rect 555927 629 555936 663
rect 555884 620 555936 629
rect 565820 620 565872 672
rect 540796 595 540848 604
rect 540796 561 540805 595
rect 540805 561 540839 595
rect 540839 561 540848 595
rect 540796 552 540848 561
rect 541992 595 542044 604
rect 541992 561 542001 595
rect 542001 561 542035 595
rect 542035 561 542044 595
rect 541992 552 542044 561
rect 550272 552 550324 604
rect 544200 484 544252 536
rect 547696 484 547748 536
rect 561404 595 561456 604
rect 561404 561 561413 595
rect 561413 561 561447 595
rect 561447 561 561456 595
rect 561404 552 561456 561
rect 562048 552 562100 604
rect 539784 459 539836 468
rect 527640 348 527692 400
rect 529664 348 529716 400
rect 539784 425 539793 459
rect 539793 425 539827 459
rect 539827 425 539836 459
rect 539784 416 539836 425
rect 550088 416 550140 468
rect 536472 348 536524 400
rect 553584 348 553636 400
rect 555792 416 555844 468
rect 573916 552 573968 604
rect 575112 552 575164 604
rect 556896 348 556948 400
rect 459376 212 459428 264
rect 461400 212 461452 264
rect 475476 212 475528 264
rect 441068 144 441120 196
rect 448980 144 449032 196
rect 462504 144 462556 196
rect 466000 144 466052 196
rect 480720 144 480772 196
rect 405740 76 405792 128
rect 350172 8 350224 60
rect 359740 8 359792 60
rect 361488 8 361540 60
rect 371884 8 371936 60
rect 376300 8 376352 60
rect 386972 8 387024 60
rect 387616 8 387668 60
rect 399116 8 399168 60
rect 399944 8 399996 60
rect 411628 76 411680 128
rect 412640 76 412692 128
rect 419448 76 419500 128
rect 434260 76 434312 128
rect 447876 76 447928 128
rect 459560 76 459612 128
rect 462412 76 462464 128
rect 477408 76 477460 128
rect 490196 280 490248 332
rect 490932 280 490984 332
rect 506204 280 506256 332
rect 507308 323 507360 332
rect 507308 289 507317 323
rect 507317 289 507351 323
rect 507351 289 507360 323
rect 507308 280 507360 289
rect 509240 280 509292 332
rect 525156 280 525208 332
rect 526260 280 526312 332
rect 543464 280 543516 332
rect 544200 280 544252 332
rect 552388 280 552440 332
rect 558000 323 558052 332
rect 558000 289 558009 323
rect 558009 289 558043 323
rect 558043 289 558052 323
rect 558000 280 558052 289
rect 559012 280 559064 332
rect 576768 280 576820 332
rect 492680 212 492732 264
rect 494428 212 494480 264
rect 499948 212 500000 264
rect 502340 212 502392 264
rect 518624 212 518676 264
rect 520372 212 520424 264
rect 536932 212 536984 264
rect 538864 212 538916 264
rect 542820 212 542872 264
rect 560668 212 560720 264
rect 562600 212 562652 264
rect 581828 212 581880 264
rect 484860 144 484912 196
rect 500316 144 500368 196
rect 503536 144 503588 196
rect 521568 144 521620 196
rect 538036 144 538088 196
rect 539876 144 539928 196
rect 557172 144 557224 196
rect 560208 144 560260 196
rect 578332 144 578384 196
rect 496820 76 496872 128
rect 500132 76 500184 128
rect 515588 76 515640 128
rect 532332 76 532384 128
rect 411536 8 411588 60
rect 429476 8 429528 60
rect 433064 8 433116 60
rect 439872 8 439924 60
rect 453488 8 453540 60
rect 455328 8 455380 60
rect 469588 8 469640 60
rect 477868 8 477920 60
rect 478512 8 478564 60
rect 490288 8 490340 60
rect 496728 8 496780 60
rect 501236 8 501288 60
rect 505744 8 505796 60
rect 521660 8 521712 60
rect 528468 8 528520 60
rect 545672 76 545724 128
rect 546500 76 546552 128
rect 564624 76 564676 128
rect 545120 8 545172 60
rect 563060 8 563112 60
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 170496 703588 170548 703594
rect 170496 703530 170548 703536
rect 1492 703384 1544 703390
rect 1492 703326 1544 703332
rect 756 702976 808 702982
rect 756 702918 808 702924
rect 388 702772 440 702778
rect 388 702714 440 702720
rect 204 702704 256 702710
rect 204 702646 256 702652
rect 18 700768 74 700777
rect 18 700703 74 700712
rect 32 71913 60 700703
rect 112 697808 164 697814
rect 112 697750 164 697756
rect 124 111217 152 697750
rect 216 163441 244 702646
rect 296 701208 348 701214
rect 296 701150 348 701156
rect 308 209774 336 701150
rect 400 229094 428 702714
rect 572 701684 624 701690
rect 572 701626 624 701632
rect 480 698760 532 698766
rect 480 698702 532 698708
rect 492 397474 520 698702
rect 584 410553 612 701626
rect 662 698184 718 698193
rect 662 698119 718 698128
rect 676 449585 704 698119
rect 768 553897 796 702918
rect 1308 701140 1360 701146
rect 1308 701082 1360 701088
rect 848 699168 900 699174
rect 848 699110 900 699116
rect 860 606121 888 699110
rect 846 606112 902 606121
rect 846 606047 902 606056
rect 754 553888 810 553897
rect 754 553823 810 553832
rect 662 449576 718 449585
rect 662 449511 718 449520
rect 570 410544 626 410553
rect 570 410479 626 410488
rect 570 397488 626 397497
rect 492 397446 570 397474
rect 570 397423 626 397432
rect 1320 249762 1348 701082
rect 1504 684321 1532 703326
rect 1584 703248 1636 703254
rect 1584 703190 1636 703196
rect 1490 684312 1546 684321
rect 1490 684247 1546 684256
rect 1596 632097 1624 703190
rect 1676 703112 1728 703118
rect 1676 703054 1728 703060
rect 1582 632088 1638 632097
rect 1582 632023 1638 632032
rect 1688 580009 1716 703054
rect 1860 702908 1912 702914
rect 1860 702850 1912 702856
rect 1766 697776 1822 697785
rect 1766 697711 1822 697720
rect 1674 580000 1730 580009
rect 1674 579935 1730 579944
rect 1780 475697 1808 697711
rect 1872 527921 1900 702850
rect 2504 702840 2556 702846
rect 2504 702782 2556 702788
rect 2044 702568 2096 702574
rect 2044 702510 2096 702516
rect 1950 698048 2006 698057
rect 1950 697983 2006 697992
rect 1858 527912 1914 527921
rect 1858 527847 1914 527856
rect 1766 475688 1822 475697
rect 1766 475623 1822 475632
rect 1964 423609 1992 697983
rect 1950 423600 2006 423609
rect 1950 423535 2006 423544
rect 1308 249756 1360 249762
rect 1308 249698 1360 249704
rect 400 229066 612 229094
rect 584 214985 612 229066
rect 570 214976 626 214985
rect 570 214911 626 214920
rect 308 209746 612 209774
rect 584 188873 612 209746
rect 570 188864 626 188873
rect 570 188799 626 188808
rect 202 163432 258 163441
rect 202 163367 258 163376
rect 110 111208 166 111217
rect 110 111143 166 111152
rect 18 71904 74 71913
rect 18 71839 74 71848
rect 2056 32473 2084 702510
rect 2134 702128 2190 702137
rect 2134 702063 2190 702072
rect 2148 58585 2176 702063
rect 2318 701584 2374 701593
rect 2318 701519 2374 701528
rect 2228 701412 2280 701418
rect 2228 701354 2280 701360
rect 2240 254153 2268 701354
rect 2226 254144 2282 254153
rect 2226 254079 2282 254088
rect 2332 84697 2360 701519
rect 2410 697640 2466 697649
rect 2410 697575 2466 697584
rect 2424 267209 2452 697575
rect 2516 319297 2544 702782
rect 6644 701956 6696 701962
rect 6644 701898 6696 701904
rect 4436 701548 4488 701554
rect 4436 701490 4488 701496
rect 4342 701448 4398 701457
rect 4342 701383 4398 701392
rect 3424 700800 3476 700806
rect 3424 700742 3476 700748
rect 2870 700632 2926 700641
rect 2870 700567 2926 700576
rect 2596 698488 2648 698494
rect 2596 698430 2648 698436
rect 2608 345409 2636 698430
rect 2686 697912 2742 697921
rect 2686 697847 2742 697856
rect 2700 371385 2728 697847
rect 2884 566953 2912 700567
rect 3238 700496 3294 700505
rect 3238 700431 3294 700440
rect 3054 700360 3110 700369
rect 3054 700295 3110 700304
rect 2870 566944 2926 566953
rect 2870 566879 2926 566888
rect 3068 514865 3096 700295
rect 3148 699644 3200 699650
rect 3148 699586 3200 699592
rect 3160 658209 3188 699586
rect 3146 658200 3202 658209
rect 3146 658135 3202 658144
rect 3054 514856 3110 514865
rect 3054 514791 3110 514800
rect 3148 502308 3200 502314
rect 3148 502250 3200 502256
rect 2686 371376 2742 371385
rect 2686 371311 2742 371320
rect 2594 345400 2650 345409
rect 2594 345335 2650 345344
rect 2502 319288 2558 319297
rect 2502 319223 2558 319232
rect 3160 306241 3188 502250
rect 3252 501809 3280 700431
rect 3332 699984 3384 699990
rect 3332 699926 3384 699932
rect 3238 501800 3294 501809
rect 3238 501735 3294 501744
rect 3344 462641 3372 699926
rect 3330 462632 3386 462641
rect 3330 462567 3386 462576
rect 3146 306232 3202 306241
rect 3146 306167 3202 306176
rect 2410 267200 2466 267209
rect 2410 267135 2466 267144
rect 2780 249756 2832 249762
rect 2780 249698 2832 249704
rect 2792 201929 2820 249698
rect 2778 201920 2834 201929
rect 2778 201855 2834 201864
rect 2318 84688 2374 84697
rect 2318 84623 2374 84632
rect 2134 58576 2190 58585
rect 2134 58511 2190 58520
rect 2042 32464 2098 32473
rect 2042 32399 2098 32408
rect 3436 19417 3464 700742
rect 3976 700596 4028 700602
rect 3976 700538 4028 700544
rect 3606 699952 3662 699961
rect 3606 699887 3662 699896
rect 3514 698592 3570 698601
rect 3514 698527 3570 698536
rect 3528 45529 3556 698527
rect 3620 149841 3648 699887
rect 3792 699712 3844 699718
rect 3792 699654 3844 699660
rect 3698 699000 3754 699009
rect 3698 698935 3754 698944
rect 3606 149832 3662 149841
rect 3606 149767 3662 149776
rect 3712 136785 3740 698935
rect 3804 619177 3832 699654
rect 3884 699508 3936 699514
rect 3884 699450 3936 699456
rect 3790 619168 3846 619177
rect 3790 619103 3846 619112
rect 3792 565888 3844 565894
rect 3792 565830 3844 565836
rect 3698 136776 3754 136785
rect 3698 136711 3754 136720
rect 3804 97617 3832 565830
rect 3896 241097 3924 699450
rect 3988 293185 4016 700538
rect 4066 700224 4122 700233
rect 4066 700159 4122 700168
rect 4080 358465 4108 700159
rect 4252 699780 4304 699786
rect 4252 699722 4304 699728
rect 4264 671265 4292 699722
rect 4250 671256 4306 671265
rect 4250 671191 4306 671200
rect 4356 565894 4384 701383
rect 4344 565888 4396 565894
rect 4344 565830 4396 565836
rect 4448 502314 4476 701490
rect 6656 699938 6684 701898
rect 8128 700330 8156 703520
rect 21456 702500 21508 702506
rect 21456 702442 21508 702448
rect 8116 700324 8168 700330
rect 8116 700266 8168 700272
rect 21468 699938 21496 702442
rect 24320 700398 24348 703520
rect 31206 701856 31262 701865
rect 31206 701791 31262 701800
rect 24308 700392 24360 700398
rect 24308 700334 24360 700340
rect 31220 699938 31248 701791
rect 40512 700466 40540 703520
rect 41052 702636 41104 702642
rect 41052 702578 41104 702584
rect 40500 700460 40552 700466
rect 40500 700402 40552 700408
rect 41064 699938 41092 702578
rect 70124 702432 70176 702438
rect 70124 702374 70176 702380
rect 55772 702024 55824 702030
rect 55772 701966 55824 701972
rect 46018 701312 46074 701321
rect 46018 701247 46074 701256
rect 46032 699938 46060 701247
rect 55784 699938 55812 701966
rect 60646 701720 60702 701729
rect 60646 701655 60702 701664
rect 60660 699938 60688 701655
rect 6440 699910 6684 699938
rect 21160 699910 21496 699938
rect 30912 699910 31248 699938
rect 40756 699910 41092 699938
rect 45724 699910 46060 699938
rect 55476 699910 55812 699938
rect 60444 699910 60688 699938
rect 70136 699666 70164 702374
rect 72988 700738 73016 703520
rect 85304 701344 85356 701350
rect 85304 701286 85356 701292
rect 75460 701276 75512 701282
rect 75460 701218 75512 701224
rect 72976 700732 73028 700738
rect 72976 700674 73028 700680
rect 75472 699938 75500 701218
rect 85316 699938 85344 701286
rect 89180 700874 89208 703520
rect 105464 703458 105492 703520
rect 105452 703452 105504 703458
rect 105452 703394 105504 703400
rect 134432 702296 134484 702302
rect 134432 702238 134484 702244
rect 100024 702160 100076 702166
rect 100024 702102 100076 702108
rect 90180 701480 90232 701486
rect 90180 701422 90232 701428
rect 89168 700868 89220 700874
rect 89168 700810 89220 700816
rect 90192 699938 90220 701422
rect 100036 699938 100064 702102
rect 119712 702092 119764 702098
rect 119712 702034 119764 702040
rect 114284 701616 114336 701622
rect 114284 701558 114336 701564
rect 104806 700088 104862 700097
rect 104806 700023 104862 700032
rect 104820 699938 104848 700023
rect 75164 699910 75500 699938
rect 85008 699910 85344 699938
rect 89884 699910 90220 699938
rect 99728 699910 100064 699938
rect 104604 699910 104848 699938
rect 114296 699666 114324 701558
rect 119724 699938 119752 702034
rect 134444 699938 134472 702238
rect 137848 700194 137876 703520
rect 144276 702228 144328 702234
rect 144276 702170 144328 702176
rect 137836 700188 137888 700194
rect 137836 700130 137888 700136
rect 144288 699938 144316 702170
rect 154028 701888 154080 701894
rect 154028 701830 154080 701836
rect 148968 701752 149020 701758
rect 148968 701694 149020 701700
rect 148980 699938 149008 701694
rect 154040 699938 154068 701830
rect 154132 700126 154160 703520
rect 170324 703474 170352 703520
rect 170508 703474 170536 703530
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 227628 703520 227680 703526
rect 235142 703520 235254 704960
rect 235448 703792 235500 703798
rect 235448 703734 235500 703740
rect 235460 703610 235488 703734
rect 235368 703582 235488 703610
rect 242440 703656 242492 703662
rect 242440 703598 242492 703604
rect 170324 703446 170536 703474
rect 198280 703180 198332 703186
rect 198280 703122 198332 703128
rect 183376 703044 183428 703050
rect 183376 702986 183428 702992
rect 163872 701820 163924 701826
rect 163872 701762 163924 701768
rect 154120 700120 154172 700126
rect 154120 700062 154172 700068
rect 163884 699938 163912 701762
rect 183388 699938 183416 702986
rect 198292 699938 198320 703122
rect 202800 702434 202828 703520
rect 213000 703316 213052 703322
rect 213000 703258 213052 703264
rect 119416 699910 119752 699938
rect 134136 699910 134472 699938
rect 143980 699910 144316 699938
rect 148856 699910 149008 699938
rect 153732 699910 154068 699938
rect 163576 699910 163912 699938
rect 183264 699910 183416 699938
rect 197984 699910 198320 699938
rect 202708 702406 202828 702434
rect 202708 699922 202736 702406
rect 213012 699938 213040 703258
rect 202696 699916 202748 699922
rect 212704 699910 213040 699938
rect 202696 699858 202748 699864
rect 218992 699854 219020 703520
rect 227628 703462 227680 703468
rect 235184 703474 235212 703520
rect 235368 703474 235396 703582
rect 227640 699938 227668 703462
rect 235184 703446 235396 703474
rect 237104 702364 237156 702370
rect 237104 702306 237156 702312
rect 232688 700528 232740 700534
rect 232688 700470 232740 700476
rect 232700 699938 232728 700470
rect 227424 699910 227668 699938
rect 232392 699910 232728 699938
rect 218980 699848 219032 699854
rect 217874 699816 217930 699825
rect 217580 699774 217874 699802
rect 218980 699790 219032 699796
rect 217874 699751 217930 699760
rect 237116 699666 237144 702306
rect 242452 699938 242480 703598
rect 251426 703520 251538 704960
rect 257252 703724 257304 703730
rect 257252 703666 257304 703672
rect 252284 700936 252336 700942
rect 252284 700878 252336 700884
rect 247408 700256 247460 700262
rect 247408 700198 247460 700204
rect 247420 699938 247448 700198
rect 252296 699938 252324 700878
rect 257264 699938 257292 703666
rect 267618 703520 267730 704960
rect 271788 703860 271840 703866
rect 271788 703802 271840 703808
rect 266360 702296 266412 702302
rect 266360 702238 266412 702244
rect 262862 701992 262918 702001
rect 259368 701956 259420 701962
rect 262862 701927 262918 701936
rect 259368 701898 259420 701904
rect 242144 699910 242480 699938
rect 247112 699910 247448 699938
rect 251988 699910 252324 699938
rect 256956 699910 257292 699938
rect 70136 699638 70288 699666
rect 114296 699638 114448 699666
rect 237116 699638 237268 699666
rect 208124 699440 208176 699446
rect 11610 699408 11666 699417
rect 11316 699366 11610 699394
rect 16394 699408 16450 699417
rect 16192 699366 16394 699394
rect 11610 699343 11666 699352
rect 65614 699408 65670 699417
rect 26036 699378 26188 699394
rect 35880 699378 36032 699394
rect 50600 699378 50936 699394
rect 26036 699372 26200 699378
rect 26036 699366 26148 699372
rect 16394 699343 16450 699352
rect 35880 699372 36044 699378
rect 35880 699366 35992 699372
rect 26148 699314 26200 699320
rect 50600 699372 50948 699378
rect 50600 699366 50896 699372
rect 35992 699314 36044 699320
rect 65320 699366 65614 699394
rect 80150 699408 80206 699417
rect 80040 699366 80150 699394
rect 65614 699343 65670 699352
rect 94852 699378 95188 699394
rect 109572 699378 109908 699394
rect 124292 699378 124628 699394
rect 129168 699378 129504 699394
rect 139012 699378 139348 699394
rect 158700 699378 158852 699394
rect 168544 699378 168880 699394
rect 173420 699378 173756 699394
rect 178296 699378 178632 699394
rect 188140 699378 188476 699394
rect 193108 699378 193260 699394
rect 202860 699378 203012 699394
rect 207828 699388 208124 699394
rect 222844 699440 222896 699446
rect 207828 699382 208176 699388
rect 222548 699388 222844 699394
rect 259380 699417 259408 701898
rect 262876 700806 262904 701927
rect 262864 700800 262916 700806
rect 262864 700742 262916 700748
rect 262128 700052 262180 700058
rect 262128 699994 262180 700000
rect 262140 699938 262168 699994
rect 261832 699910 262168 699938
rect 266372 699582 266400 702238
rect 267004 701072 267056 701078
rect 267004 701014 267056 701020
rect 267016 699938 267044 701014
rect 267660 701010 267688 703520
rect 267648 701004 267700 701010
rect 267648 700946 267700 700952
rect 271800 699938 271828 703802
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 300860 703792 300912 703798
rect 300860 703734 300912 703740
rect 277400 702296 277452 702302
rect 277400 702238 277452 702244
rect 276848 700664 276900 700670
rect 276848 700606 276900 700612
rect 276860 699938 276888 700606
rect 266708 699910 267044 699938
rect 271676 699910 271828 699938
rect 276552 699910 276888 699938
rect 277308 699984 277360 699990
rect 277308 699926 277360 699932
rect 277320 699802 277348 699926
rect 277412 699802 277440 702238
rect 280896 701956 280948 701962
rect 280896 701898 280948 701904
rect 278596 701072 278648 701078
rect 278596 701014 278648 701020
rect 278608 699990 278636 701014
rect 280908 700602 280936 701898
rect 281356 700800 281408 700806
rect 281356 700742 281408 700748
rect 280896 700596 280948 700602
rect 280896 700538 280948 700544
rect 278596 699984 278648 699990
rect 278596 699926 278648 699932
rect 277320 699774 277440 699802
rect 281368 699802 281396 700742
rect 283852 700602 283880 703520
rect 291844 702364 291896 702370
rect 291844 702306 291896 702312
rect 291856 701010 291884 702306
rect 292488 701072 292540 701078
rect 292488 701014 292540 701020
rect 295892 701072 295944 701078
rect 295892 701014 295944 701020
rect 291384 701004 291436 701010
rect 291384 700946 291436 700952
rect 291844 701004 291896 701010
rect 291844 700946 291896 700952
rect 283840 700596 283892 700602
rect 283840 700538 283892 700544
rect 286690 699816 286746 699825
rect 281368 699774 281520 699802
rect 286396 699774 286690 699802
rect 286690 699751 286746 699760
rect 291396 699666 291424 700946
rect 292500 700602 292528 701014
rect 292488 700596 292540 700602
rect 292488 700538 292540 700544
rect 295904 699938 295932 701014
rect 300136 700602 300164 703520
rect 298100 700596 298152 700602
rect 298100 700538 298152 700544
rect 300124 700596 300176 700602
rect 300124 700538 300176 700544
rect 295904 699910 296240 699938
rect 298112 699825 298140 700538
rect 300872 699938 300900 703734
rect 315488 703588 315540 703594
rect 315488 703530 315540 703536
rect 311992 702160 312044 702166
rect 311992 702102 312044 702108
rect 305000 702024 305052 702030
rect 305000 701966 305052 701972
rect 305012 700602 305040 701966
rect 311900 701072 311952 701078
rect 311900 701014 311952 701020
rect 305000 700596 305052 700602
rect 305000 700538 305052 700544
rect 300872 699910 301116 699938
rect 305748 699922 306084 699938
rect 305736 699916 306084 699922
rect 305788 699910 306084 699916
rect 305736 699858 305788 699864
rect 310612 699848 310664 699854
rect 298098 699816 298154 699825
rect 310664 699796 310960 699802
rect 310612 699790 310960 699796
rect 310624 699774 310960 699790
rect 298098 699751 298154 699760
rect 291272 699638 291424 699666
rect 311912 699650 311940 701014
rect 312004 699922 312032 702102
rect 315500 699938 315528 703530
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364708 703860 364760 703866
rect 364708 703802 364760 703808
rect 364720 703610 364748 703802
rect 364720 703582 364840 703610
rect 330300 703452 330352 703458
rect 330300 703394 330352 703400
rect 324320 702228 324372 702234
rect 324320 702170 324372 702176
rect 324332 700194 324360 702170
rect 320778 700188 320830 700194
rect 320778 700130 320830 700136
rect 324320 700188 324372 700194
rect 324320 700130 324372 700136
rect 311992 699916 312044 699922
rect 315500 699910 315836 699938
rect 320790 699924 320818 700130
rect 325654 700120 325706 700126
rect 325654 700062 325706 700068
rect 325666 699924 325694 700062
rect 330312 699938 330340 703394
rect 332520 700670 332548 703520
rect 340144 702092 340196 702098
rect 340144 702034 340196 702040
rect 338028 702024 338080 702030
rect 338028 701966 338080 701972
rect 336646 701856 336702 701865
rect 336646 701791 336702 701800
rect 336660 700738 336688 701791
rect 335360 700732 335412 700738
rect 335360 700674 335412 700680
rect 336648 700732 336700 700738
rect 336648 700674 336700 700680
rect 332508 700664 332560 700670
rect 332508 700606 332560 700612
rect 330312 699910 330648 699938
rect 311992 699858 312044 699864
rect 335372 699802 335400 700674
rect 335372 699774 335524 699802
rect 311900 699644 311952 699650
rect 311900 699586 311952 699592
rect 266360 699576 266412 699582
rect 266360 699518 266412 699524
rect 338040 699514 338068 701966
rect 340156 700874 340184 702034
rect 340052 700868 340104 700874
rect 340052 700810 340104 700816
rect 340144 700868 340196 700874
rect 340144 700810 340196 700816
rect 340064 699938 340092 700810
rect 348804 700806 348832 703520
rect 364812 703474 364840 703582
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 394700 703724 394752 703730
rect 394700 703666 394752 703672
rect 364996 703474 365024 703520
rect 364812 703446 365024 703474
rect 359740 703384 359792 703390
rect 359740 703326 359792 703332
rect 348792 700800 348844 700806
rect 348792 700742 348844 700748
rect 345204 700460 345256 700466
rect 345204 700402 345256 700408
rect 345216 699938 345244 700402
rect 354956 700392 355008 700398
rect 354956 700334 355008 700340
rect 349896 700324 349948 700330
rect 349896 700266 349948 700272
rect 349908 699938 349936 700266
rect 354968 699938 354996 700334
rect 359752 699938 359780 703326
rect 374460 703248 374512 703254
rect 374460 703190 374512 703196
rect 364616 701072 364668 701078
rect 364616 701014 364668 701020
rect 364628 699938 364656 701014
rect 374472 699938 374500 703190
rect 389180 703112 389232 703118
rect 389180 703054 389232 703060
rect 389192 699938 389220 703054
rect 394148 702976 394200 702982
rect 394148 702918 394200 702924
rect 394160 699938 394188 702918
rect 394712 700398 394740 703666
rect 397430 703520 397542 704960
rect 400864 703656 400916 703662
rect 400864 703598 400916 703604
rect 394700 700392 394752 700398
rect 394700 700334 394752 700340
rect 397472 700058 397500 703520
rect 399022 700632 399078 700641
rect 399022 700567 399078 700576
rect 397460 700052 397512 700058
rect 397460 699994 397512 700000
rect 399036 699938 399064 700567
rect 400876 700466 400904 703598
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 468484 703520 468536 703526
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 403900 702908 403952 702914
rect 403900 702850 403952 702856
rect 400864 700460 400916 700466
rect 400864 700402 400916 700408
rect 403912 699938 403940 702850
rect 408866 700496 408922 700505
rect 408866 700431 408922 700440
rect 408880 699938 408908 700431
rect 413664 699990 413692 703520
rect 428464 702296 428516 702302
rect 428464 702238 428516 702244
rect 414202 700360 414258 700369
rect 414202 700295 414258 700304
rect 413652 699984 413704 699990
rect 340064 699910 340400 699938
rect 345216 699910 345368 699938
rect 349908 699910 350244 699938
rect 354968 699910 355212 699938
rect 359752 699910 360088 699938
rect 364628 699910 364964 699938
rect 374472 699910 374808 699938
rect 389192 699910 389528 699938
rect 394160 699910 394496 699938
rect 399036 699910 399372 699938
rect 403912 699910 404248 699938
rect 408880 699910 409216 699938
rect 413652 699926 413704 699932
rect 369780 699786 369932 699802
rect 369768 699780 369932 699786
rect 369820 699774 369932 699780
rect 369768 699722 369820 699728
rect 384304 699712 384356 699718
rect 414216 699666 414244 700295
rect 428476 699938 428504 702238
rect 429856 700398 429884 703520
rect 443276 701684 443328 701690
rect 443276 701626 443328 701632
rect 429844 700392 429896 700398
rect 429844 700334 429896 700340
rect 443288 699938 443316 701626
rect 462332 700262 462360 703520
rect 468484 703462 468536 703468
rect 462872 702840 462924 702846
rect 462872 702782 462924 702788
rect 462320 700256 462372 700262
rect 458316 700224 458372 700233
rect 462320 700198 462372 700204
rect 458316 700159 458372 700168
rect 428476 699910 428812 699938
rect 443288 699910 443624 699938
rect 458330 699924 458358 700159
rect 462884 699938 462912 702782
rect 467840 701956 467892 701962
rect 467840 701898 467892 701904
rect 467852 699938 467880 701898
rect 468496 700806 468524 703462
rect 472716 701548 472768 701554
rect 472716 701490 472768 701496
rect 468576 701072 468628 701078
rect 468576 701014 468628 701020
rect 468484 700800 468536 700806
rect 468484 700742 468536 700748
rect 462884 699910 463220 699938
rect 467852 699910 468188 699938
rect 384356 699660 384652 699666
rect 384304 699654 384652 699660
rect 384316 699638 384652 699654
rect 414092 699638 414244 699666
rect 379532 699514 379776 699530
rect 438320 699514 438656 699530
rect 453040 699514 453376 699530
rect 338028 699508 338080 699514
rect 338028 699450 338080 699456
rect 379520 699508 379776 699514
rect 379572 699502 379776 699508
rect 438308 699508 438656 699514
rect 379520 699450 379572 699456
rect 438360 699502 438656 699508
rect 453028 699508 453376 699514
rect 438308 699450 438360 699456
rect 453080 699502 453376 699508
rect 453028 699450 453080 699456
rect 468588 699417 468616 701014
rect 472728 699938 472756 701490
rect 478524 700942 478552 703520
rect 492680 702772 492732 702778
rect 492680 702714 492732 702720
rect 482560 702024 482612 702030
rect 482560 701966 482612 701972
rect 478512 700936 478564 700942
rect 478512 700878 478564 700884
rect 482572 699938 482600 701966
rect 487436 701412 487488 701418
rect 487436 701354 487488 701360
rect 487448 699938 487476 701354
rect 492692 700210 492720 702714
rect 494808 700466 494836 703520
rect 507124 702704 507176 702710
rect 507124 702646 507176 702652
rect 497280 701208 497332 701214
rect 497280 701150 497332 701156
rect 494796 700460 494848 700466
rect 494796 700402 494848 700408
rect 492692 700182 492766 700210
rect 472728 699910 473064 699938
rect 482572 699910 482908 699938
rect 487448 699910 487784 699938
rect 492738 699924 492766 700182
rect 497292 699938 497320 701150
rect 502340 701140 502392 701146
rect 502340 701082 502392 701088
rect 502352 699938 502380 701082
rect 507136 699938 507164 702646
rect 526718 701584 526774 701593
rect 526718 701519 526774 701528
rect 512000 701072 512052 701078
rect 512000 701014 512052 701020
rect 512012 699938 512040 701014
rect 516966 699952 517022 699961
rect 497292 699910 497628 699938
rect 502352 699910 502504 699938
rect 507136 699910 507472 699938
rect 512012 699910 512348 699938
rect 526732 699938 526760 701519
rect 527192 700534 527220 703520
rect 531686 701448 531742 701457
rect 531686 701383 531742 701392
rect 527180 700528 527232 700534
rect 527180 700470 527232 700476
rect 531700 699938 531728 701383
rect 543476 701010 543504 703520
rect 551284 702568 551336 702574
rect 551284 702510 551336 702516
rect 546498 702128 546554 702137
rect 546498 702063 546554 702072
rect 543464 701004 543516 701010
rect 543464 700946 543516 700952
rect 537022 700768 537078 700777
rect 537022 700703 537078 700712
rect 517022 699910 517316 699938
rect 526732 699910 527068 699938
rect 531700 699910 532036 699938
rect 516966 699887 517022 699896
rect 537036 699666 537064 700703
rect 546512 699938 546540 702063
rect 551296 699938 551324 702510
rect 556896 701140 556948 701146
rect 556896 701082 556948 701088
rect 556908 699938 556936 701082
rect 559668 700806 559696 703520
rect 576308 703316 576360 703322
rect 576308 703258 576360 703264
rect 575020 703180 575072 703186
rect 575020 703122 575072 703128
rect 573640 703044 573692 703050
rect 573640 702986 573692 702992
rect 573456 702432 573508 702438
rect 573456 702374 573508 702380
rect 561126 701992 561182 702001
rect 561126 701927 561182 701936
rect 559656 700800 559708 700806
rect 559656 700742 559708 700748
rect 546512 699910 546756 699938
rect 551296 699910 551632 699938
rect 556600 699910 556936 699938
rect 561140 699938 561168 701927
rect 565360 701888 565412 701894
rect 565360 701830 565412 701836
rect 564440 701140 564492 701146
rect 564440 701082 564492 701088
rect 561140 699910 561476 699938
rect 536912 699638 537064 699666
rect 521856 699514 522192 699530
rect 521844 699508 522192 699514
rect 521896 699502 522192 699508
rect 521844 699450 521896 699456
rect 222548 699382 222896 699388
rect 259366 699408 259422 699417
rect 94852 699372 95200 699378
rect 94852 699366 95148 699372
rect 80150 699343 80206 699352
rect 50896 699314 50948 699320
rect 109572 699372 109920 699378
rect 109572 699366 109868 699372
rect 95148 699314 95200 699320
rect 124292 699372 124640 699378
rect 124292 699366 124588 699372
rect 109868 699314 109920 699320
rect 129168 699372 129516 699378
rect 129168 699366 129464 699372
rect 124588 699314 124640 699320
rect 139012 699372 139360 699378
rect 139012 699366 139308 699372
rect 129464 699314 129516 699320
rect 158700 699372 158864 699378
rect 158700 699366 158812 699372
rect 139308 699314 139360 699320
rect 168544 699372 168892 699378
rect 168544 699366 168840 699372
rect 158812 699314 158864 699320
rect 173420 699372 173768 699378
rect 173420 699366 173716 699372
rect 168840 699314 168892 699320
rect 178296 699372 178644 699378
rect 178296 699366 178592 699372
rect 173716 699314 173768 699320
rect 188140 699372 188488 699378
rect 188140 699366 188436 699372
rect 178592 699314 178644 699320
rect 193108 699372 193272 699378
rect 193108 699366 193220 699372
rect 188436 699314 188488 699320
rect 202860 699372 203024 699378
rect 202860 699366 202972 699372
rect 193220 699314 193272 699320
rect 207828 699366 208164 699382
rect 222548 699366 222884 699382
rect 259366 699343 259422 699352
rect 418710 699408 418766 699417
rect 423678 699408 423734 699417
rect 418766 699366 419060 699394
rect 418710 699343 418766 699352
rect 433430 699408 433486 699417
rect 423734 699366 423936 699394
rect 423678 699343 423734 699352
rect 448150 699408 448206 699417
rect 433486 699366 433780 699394
rect 433430 699343 433486 699352
rect 468574 699408 468630 699417
rect 448206 699366 448500 699394
rect 448150 699343 448206 699352
rect 468574 699343 468630 699352
rect 477590 699408 477646 699417
rect 541530 699408 541586 699417
rect 477646 699366 477940 699394
rect 477590 699343 477646 699352
rect 541586 699366 541880 699394
rect 563704 699372 563756 699378
rect 541530 699343 541586 699352
rect 202972 699314 203024 699320
rect 563704 699314 563756 699320
rect 563716 644434 563744 699314
rect 563704 644428 563756 644434
rect 563704 644370 563756 644376
rect 4436 502308 4488 502314
rect 4436 502250 4488 502256
rect 4066 358456 4122 358465
rect 4066 358391 4122 358400
rect 3974 293176 4030 293185
rect 3974 293111 4030 293120
rect 3882 241088 3938 241097
rect 3882 241023 3938 241032
rect 3790 97608 3846 97617
rect 3790 97543 3846 97552
rect 3514 45520 3570 45529
rect 3514 45455 3570 45464
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 3054 6488 3110 6497
rect 3054 6423 3110 6432
rect 3068 1358 3096 6423
rect 563612 3188 563664 3194
rect 563612 3130 563664 3136
rect 563520 2916 563572 2922
rect 563520 2858 563572 2864
rect 3056 1352 3108 1358
rect 3056 1294 3108 1300
rect 563532 1086 563560 2858
rect 563520 1080 563572 1086
rect 563520 1022 563572 1028
rect 563624 950 563652 3130
rect 563704 3052 563756 3058
rect 563704 2994 563756 3000
rect 563612 944 563664 950
rect 563612 886 563664 892
rect 563716 762 563744 2994
rect 564452 1358 564480 701082
rect 565266 698728 565322 698737
rect 565266 698663 565322 698672
rect 565082 698456 565138 698465
rect 565082 698391 565138 698400
rect 565096 20670 565124 698391
rect 565176 698352 565228 698358
rect 565176 698294 565228 698300
rect 565188 245614 565216 698294
rect 565176 245608 565228 245614
rect 565176 245550 565228 245556
rect 565280 167006 565308 698663
rect 565372 458182 565400 701830
rect 569314 701720 569370 701729
rect 569314 701655 569370 701664
rect 566556 701480 566608 701486
rect 566556 701422 566608 701428
rect 566462 698320 566518 698329
rect 566462 698255 566518 698264
rect 565360 458176 565412 458182
rect 565360 458118 565412 458124
rect 565268 167000 565320 167006
rect 565268 166942 565320 166948
rect 566476 33114 566504 698255
rect 566568 219434 566596 701422
rect 567844 699236 567896 699242
rect 567844 699178 567896 699184
rect 566646 698864 566702 698873
rect 566646 698799 566702 698808
rect 566556 219428 566608 219434
rect 566556 219370 566608 219376
rect 566660 206990 566688 698799
rect 566740 698692 566792 698698
rect 566740 698634 566792 698640
rect 566752 379506 566780 698634
rect 567856 578202 567884 699178
rect 569224 697604 569276 697610
rect 569224 697546 569276 697552
rect 567844 578196 567896 578202
rect 567844 578138 567896 578144
rect 566740 379500 566792 379506
rect 566740 379442 566792 379448
rect 566648 206984 566700 206990
rect 566648 206926 566700 206932
rect 569236 73166 569264 697546
rect 569328 139398 569356 701655
rect 570696 701344 570748 701350
rect 570696 701286 570748 701292
rect 570604 701276 570656 701282
rect 570604 701218 570656 701224
rect 569592 699032 569644 699038
rect 569592 698974 569644 698980
rect 569500 698896 569552 698902
rect 569500 698838 569552 698844
rect 569408 698420 569460 698426
rect 569408 698362 569460 698368
rect 569420 299470 569448 698362
rect 569512 511970 569540 698838
rect 569604 525774 569632 698974
rect 569592 525768 569644 525774
rect 569592 525710 569644 525716
rect 569500 511964 569552 511970
rect 569500 511906 569552 511912
rect 569408 299464 569460 299470
rect 569408 299406 569460 299412
rect 570616 179382 570644 701218
rect 570708 233238 570736 701286
rect 571982 700088 572038 700097
rect 571982 700023 572038 700032
rect 570880 699304 570932 699310
rect 570880 699246 570932 699252
rect 570788 698556 570840 698562
rect 570788 698498 570840 698504
rect 570800 353258 570828 698498
rect 570892 632058 570920 699246
rect 570880 632052 570932 632058
rect 570880 631994 570932 632000
rect 570788 353252 570840 353258
rect 570788 353194 570840 353200
rect 571996 259418 572024 700023
rect 572168 699440 572220 699446
rect 572168 699382 572220 699388
rect 572076 698828 572128 698834
rect 572076 698770 572128 698776
rect 572088 485790 572116 698770
rect 572180 684486 572208 699382
rect 573364 697740 573416 697746
rect 573364 697682 573416 697688
rect 572168 684480 572220 684486
rect 572168 684422 572220 684428
rect 572076 485784 572128 485790
rect 572076 485726 572128 485732
rect 571984 259412 572036 259418
rect 571984 259354 572036 259360
rect 570696 233232 570748 233238
rect 570696 233174 570748 233180
rect 570604 179376 570656 179382
rect 570604 179318 570656 179324
rect 569316 139392 569368 139398
rect 569316 139334 569368 139340
rect 573376 126954 573404 697682
rect 573468 193186 573496 702374
rect 573548 698964 573600 698970
rect 573548 698906 573600 698912
rect 573560 538218 573588 698906
rect 573652 564398 573680 702986
rect 574928 701752 574980 701758
rect 574928 701694 574980 701700
rect 574836 701616 574888 701622
rect 574836 701558 574888 701564
rect 574744 697672 574796 697678
rect 574744 697614 574796 697620
rect 573640 564392 573692 564398
rect 573640 564334 573692 564340
rect 573548 538212 573600 538218
rect 573548 538154 573600 538160
rect 573456 193180 573508 193186
rect 573456 193122 573508 193128
rect 573364 126948 573416 126954
rect 573364 126890 573416 126896
rect 574756 86970 574784 697614
rect 574848 325650 574876 701558
rect 574940 419490 574968 701694
rect 575032 618254 575060 703122
rect 576124 702500 576176 702506
rect 576124 702442 576176 702448
rect 575020 618248 575072 618254
rect 575020 618190 575072 618196
rect 574928 419484 574980 419490
rect 574928 419426 574980 419432
rect 574836 325644 574888 325650
rect 574836 325586 574888 325592
rect 574744 86964 574796 86970
rect 574744 86906 574796 86912
rect 569224 73160 569276 73166
rect 569224 73102 569276 73108
rect 576136 46918 576164 702442
rect 576216 699100 576268 699106
rect 576216 699042 576268 699048
rect 576228 592006 576256 699042
rect 576320 672042 576348 703258
rect 578884 702636 578936 702642
rect 578884 702578 578936 702584
rect 577596 701820 577648 701826
rect 577596 701762 577648 701768
rect 577502 701312 577558 701321
rect 577502 701247 577558 701256
rect 576308 672036 576360 672042
rect 576308 671978 576360 671984
rect 576216 592000 576268 592006
rect 576216 591942 576268 591948
rect 577516 100706 577544 701247
rect 577608 471986 577636 701762
rect 577596 471980 577648 471986
rect 577596 471922 577648 471928
rect 578896 112849 578924 702578
rect 580632 700868 580684 700874
rect 580632 700810 580684 700816
rect 580356 700732 580408 700738
rect 580356 700674 580408 700680
rect 580262 699136 580318 699145
rect 580262 699071 580318 699080
rect 578976 698624 579028 698630
rect 578976 698566 579028 698572
rect 578988 404977 579016 698566
rect 580172 684480 580224 684486
rect 580172 684422 580224 684428
rect 580184 683913 580212 684422
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580172 672036 580224 672042
rect 580172 671978 580224 671984
rect 580184 670721 580212 671978
rect 580170 670712 580226 670721
rect 580170 670647 580226 670656
rect 580172 644428 580224 644434
rect 580172 644370 580224 644376
rect 580184 644065 580212 644370
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580172 632052 580224 632058
rect 580172 631994 580224 632000
rect 580184 630873 580212 631994
rect 580170 630864 580226 630873
rect 580170 630799 580226 630808
rect 580172 618248 580224 618254
rect 580172 618190 580224 618196
rect 580184 617545 580212 618190
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 579988 592000 580040 592006
rect 579988 591942 580040 591948
rect 580000 591025 580028 591942
rect 579986 591016 580042 591025
rect 579986 590951 580042 590960
rect 579804 578196 579856 578202
rect 579804 578138 579856 578144
rect 579816 577697 579844 578138
rect 579802 577688 579858 577697
rect 579802 577623 579858 577632
rect 580172 564392 580224 564398
rect 580170 564360 580172 564369
rect 580224 564360 580226 564369
rect 580170 564295 580226 564304
rect 580172 538212 580224 538218
rect 580172 538154 580224 538160
rect 580184 537849 580212 538154
rect 580170 537840 580226 537849
rect 580170 537775 580226 537784
rect 580172 525768 580224 525774
rect 580172 525710 580224 525716
rect 580184 524521 580212 525710
rect 580170 524512 580226 524521
rect 580170 524447 580226 524456
rect 580172 511964 580224 511970
rect 580172 511906 580224 511912
rect 580184 511329 580212 511906
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 580172 485784 580224 485790
rect 580172 485726 580224 485732
rect 580184 484673 580212 485726
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 580172 458176 580224 458182
rect 580170 458144 580172 458153
rect 580224 458144 580226 458153
rect 580170 458079 580226 458088
rect 580172 419484 580224 419490
rect 580172 419426 580224 419432
rect 580184 418305 580212 419426
rect 580170 418296 580226 418305
rect 580170 418231 580226 418240
rect 578974 404968 579030 404977
rect 578974 404903 579030 404912
rect 580172 379500 580224 379506
rect 580172 379442 580224 379448
rect 580184 378457 580212 379442
rect 580170 378448 580226 378457
rect 580170 378383 580226 378392
rect 580172 353252 580224 353258
rect 580172 353194 580224 353200
rect 580184 351937 580212 353194
rect 580170 351928 580226 351937
rect 580170 351863 580226 351872
rect 579988 325644 580040 325650
rect 579988 325586 580040 325592
rect 580000 325281 580028 325586
rect 579986 325272 580042 325281
rect 579986 325207 580042 325216
rect 580172 299464 580224 299470
rect 580172 299406 580224 299412
rect 580184 298761 580212 299406
rect 580170 298752 580226 298761
rect 580170 298687 580226 298696
rect 580172 259412 580224 259418
rect 580172 259354 580224 259360
rect 580184 258913 580212 259354
rect 580170 258904 580226 258913
rect 580170 258839 580226 258848
rect 580172 245608 580224 245614
rect 580170 245576 580172 245585
rect 580224 245576 580226 245585
rect 580170 245511 580226 245520
rect 579620 233232 579672 233238
rect 579620 233174 579672 233180
rect 579632 232393 579660 233174
rect 579618 232384 579674 232393
rect 579618 232319 579674 232328
rect 580172 219428 580224 219434
rect 580172 219370 580224 219376
rect 580184 219065 580212 219370
rect 580170 219056 580226 219065
rect 580170 218991 580226 219000
rect 580172 206984 580224 206990
rect 580172 206926 580224 206932
rect 580184 205737 580212 206926
rect 580170 205728 580226 205737
rect 580170 205663 580226 205672
rect 580172 193180 580224 193186
rect 580172 193122 580224 193128
rect 580184 192545 580212 193122
rect 580170 192536 580226 192545
rect 580170 192471 580226 192480
rect 580172 179376 580224 179382
rect 580172 179318 580224 179324
rect 580184 179217 580212 179318
rect 580170 179208 580226 179217
rect 580170 179143 580226 179152
rect 580172 167000 580224 167006
rect 580172 166942 580224 166948
rect 580184 165889 580212 166942
rect 580170 165880 580226 165889
rect 580170 165815 580226 165824
rect 580172 139392 580224 139398
rect 580170 139360 580172 139369
rect 580224 139360 580226 139369
rect 580170 139295 580226 139304
rect 580172 126948 580224 126954
rect 580172 126890 580224 126896
rect 580184 126041 580212 126890
rect 580170 126032 580226 126041
rect 580170 125967 580226 125976
rect 578882 112840 578938 112849
rect 578882 112775 578938 112784
rect 577504 100700 577556 100706
rect 577504 100642 577556 100648
rect 579804 100700 579856 100706
rect 579804 100642 579856 100648
rect 579816 99521 579844 100642
rect 579802 99512 579858 99521
rect 579802 99447 579858 99456
rect 579620 86964 579672 86970
rect 579620 86906 579672 86912
rect 579632 86193 579660 86906
rect 579618 86184 579674 86193
rect 579618 86119 579674 86128
rect 580172 73160 580224 73166
rect 580172 73102 580224 73108
rect 580184 73001 580212 73102
rect 580170 72992 580226 73001
rect 580170 72927 580226 72936
rect 576124 46912 576176 46918
rect 576124 46854 576176 46860
rect 580172 46912 580224 46918
rect 580172 46854 580224 46860
rect 580184 46345 580212 46854
rect 580170 46336 580226 46345
rect 580170 46271 580226 46280
rect 580170 33144 580226 33153
rect 566464 33108 566516 33114
rect 580170 33079 580172 33088
rect 566464 33050 566516 33056
rect 580224 33079 580226 33088
rect 580172 33050 580224 33056
rect 565084 20664 565136 20670
rect 565084 20606 565136 20612
rect 580172 20664 580224 20670
rect 580172 20606 580224 20612
rect 580184 19825 580212 20606
rect 580170 19816 580226 19825
rect 580170 19751 580226 19760
rect 580276 6633 580304 699071
rect 580368 59673 580396 700674
rect 580448 700596 580500 700602
rect 580448 700538 580500 700544
rect 580460 152697 580488 700538
rect 580540 699916 580592 699922
rect 580540 699858 580592 699864
rect 580552 272241 580580 699858
rect 580644 312089 580672 700810
rect 580816 700188 580868 700194
rect 580816 700130 580868 700136
rect 580724 699576 580776 699582
rect 580724 699518 580776 699524
rect 580736 365129 580764 699518
rect 580828 431633 580856 700130
rect 580908 471980 580960 471986
rect 580908 471922 580960 471928
rect 580920 471481 580948 471922
rect 580906 471472 580962 471481
rect 580906 471407 580962 471416
rect 580814 431624 580870 431633
rect 580814 431559 580870 431568
rect 580722 365120 580778 365129
rect 580722 365055 580778 365064
rect 580630 312080 580686 312089
rect 580630 312015 580686 312024
rect 580538 272232 580594 272241
rect 580538 272167 580594 272176
rect 580446 152688 580502 152697
rect 580446 152623 580502 152632
rect 580354 59664 580410 59673
rect 580354 59599 580410 59608
rect 580262 6624 580318 6633
rect 580262 6559 580318 6568
rect 569132 3188 569184 3194
rect 569132 3130 569184 3136
rect 565912 3120 565964 3126
rect 565912 3062 565964 3068
rect 564440 1352 564492 1358
rect 564440 1294 564492 1300
rect 565924 882 565952 3062
rect 566832 1216 566884 1222
rect 566832 1158 566884 1164
rect 565912 876 565964 882
rect 565912 818 565964 824
rect 1676 672 1728 678
rect 5356 672 5408 678
rect 1676 614 1728 620
rect 4066 640 4122 649
rect 572 604 624 610
rect 572 546 624 552
rect 584 480 612 546
rect 1688 480 1716 614
rect 2884 564 3096 592
rect 4356 610 4600 626
rect 6460 672 6512 678
rect 5408 620 5704 626
rect 5356 614 5704 620
rect 10048 672 10100 678
rect 7838 640 7894 649
rect 6460 614 6512 620
rect 4066 575 4122 584
rect 4344 604 4600 610
rect 2884 480 2912 564
rect 3068 490 3096 564
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 3068 474 3280 490
rect 4080 480 4108 575
rect 4396 598 4600 604
rect 5264 604 5316 610
rect 4344 546 4396 552
rect 5368 598 5704 614
rect 5264 546 5316 552
rect 5276 480 5304 546
rect 6472 480 6500 614
rect 7484 598 7696 626
rect 7484 542 7512 598
rect 7472 536 7524 542
rect 3068 468 3292 474
rect 3068 462 3240 468
rect 3240 410 3292 416
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 6656 474 6808 490
rect 7472 478 7524 484
rect 7668 480 7696 598
rect 9954 640 10010 649
rect 7894 598 8004 626
rect 8588 598 8800 626
rect 8864 610 9108 626
rect 7838 575 7894 584
rect 8588 542 8616 598
rect 8576 536 8628 542
rect 6644 468 6808 474
rect 6696 462 6808 468
rect 6644 410 6696 416
rect 7626 -960 7738 480
rect 8576 478 8628 484
rect 8772 480 8800 598
rect 8852 604 9108 610
rect 8904 598 9108 604
rect 11520 672 11572 678
rect 10100 620 10212 626
rect 10048 614 10212 620
rect 10060 598 10212 614
rect 11408 620 11520 626
rect 19432 672 19484 678
rect 11408 614 11572 620
rect 13266 640 13322 649
rect 11152 604 11204 610
rect 9954 575 10010 584
rect 8852 546 8904 552
rect 9968 480 9996 575
rect 11408 598 11560 614
rect 12348 604 12400 610
rect 11152 546 11204 552
rect 13322 598 13616 626
rect 14476 598 14812 626
rect 15580 610 15916 626
rect 15568 604 15916 610
rect 13266 575 13322 584
rect 12348 546 12400 552
rect 11164 480 11192 546
rect 12360 480 12388 546
rect 12624 536 12676 542
rect 12512 484 12624 490
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 12512 478 12676 484
rect 13360 536 13412 542
rect 13360 478 13412 484
rect 12512 462 12664 478
rect 13372 354 13400 478
rect 13514 354 13626 480
rect 14476 474 14504 598
rect 15620 598 15916 604
rect 16684 598 17020 626
rect 17880 598 18216 626
rect 22376 672 22428 678
rect 19432 614 19484 620
rect 20626 640 20682 649
rect 15568 546 15620 552
rect 16684 542 16712 598
rect 16672 536 16724 542
rect 14464 468 14516 474
rect 14464 410 14516 416
rect 14556 468 14608 474
rect 14556 410 14608 416
rect 13372 326 13626 354
rect 14568 354 14596 410
rect 14710 354 14822 480
rect 14568 326 14822 354
rect 13514 -960 13626 326
rect 14710 -960 14822 326
rect 15906 82 16018 480
rect 16672 478 16724 484
rect 17408 536 17460 542
rect 17010 354 17122 480
rect 17408 478 17460 484
rect 17420 354 17448 478
rect 17880 474 17908 598
rect 18510 504 18566 513
rect 17868 468 17920 474
rect 17868 410 17920 416
rect 17010 326 17448 354
rect 16304 128 16356 134
rect 15906 76 16304 82
rect 15906 70 16356 76
rect 15906 54 16344 70
rect 15906 -960 16018 54
rect 17010 -960 17122 326
rect 18206 218 18318 480
rect 19444 480 19472 614
rect 24860 672 24912 678
rect 23478 640 23534 649
rect 22428 620 22724 626
rect 22376 614 22724 620
rect 20626 575 20682 584
rect 21824 604 21876 610
rect 20076 536 20128 542
rect 20128 484 20424 490
rect 18510 439 18566 448
rect 18524 218 18552 439
rect 18206 190 18552 218
rect 18206 -960 18318 190
rect 18972 128 19024 134
rect 19024 76 19320 82
rect 18972 70 19320 76
rect 18984 54 19320 70
rect 19402 -960 19514 480
rect 20076 478 20424 484
rect 20640 480 20668 575
rect 22388 598 22724 614
rect 23020 604 23072 610
rect 21824 546 21876 552
rect 23534 598 23828 626
rect 25320 672 25372 678
rect 24912 620 25024 626
rect 24860 614 25024 620
rect 28080 672 28132 678
rect 26514 640 26570 649
rect 25320 614 25372 620
rect 24872 598 25024 614
rect 23478 575 23534 584
rect 23020 546 23072 552
rect 24228 564 24440 592
rect 21270 504 21326 513
rect 20088 462 20424 478
rect 20598 -960 20710 480
rect 21326 462 21620 490
rect 21836 480 21864 546
rect 23032 480 23060 546
rect 24228 480 24256 564
rect 21270 439 21326 448
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 24412 474 24440 564
rect 25332 480 25360 614
rect 25792 610 26128 626
rect 25780 604 26128 610
rect 25832 598 26128 604
rect 28724 672 28776 678
rect 28722 640 28724 649
rect 29184 672 29236 678
rect 28776 640 28778 649
rect 28132 620 28428 626
rect 28080 614 28428 620
rect 28092 598 28428 614
rect 26514 575 26570 584
rect 25780 546 25832 552
rect 26528 480 26556 575
rect 27724 564 27936 592
rect 31300 672 31352 678
rect 30286 640 30342 649
rect 29236 620 29532 626
rect 29184 614 29532 620
rect 28722 575 28778 584
rect 28816 604 28868 610
rect 24400 468 24452 474
rect 24400 410 24452 416
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 26896 474 27232 490
rect 27724 480 27752 564
rect 27908 513 27936 564
rect 29196 598 29532 614
rect 30104 604 30156 610
rect 28868 564 28948 592
rect 28816 546 28868 552
rect 27894 504 27950 513
rect 26884 468 27232 474
rect 26936 462 27232 468
rect 26884 410 26936 416
rect 27682 -960 27794 480
rect 28920 480 28948 564
rect 30342 598 30636 626
rect 33784 672 33836 678
rect 31300 614 31352 620
rect 32402 640 32458 649
rect 30286 575 30342 584
rect 30104 546 30156 552
rect 30116 480 30144 546
rect 31312 480 31340 614
rect 33230 640 33286 649
rect 32600 610 32936 626
rect 32402 575 32458 584
rect 32588 604 32936 610
rect 31668 536 31720 542
rect 31720 484 31832 490
rect 27894 439 27950 448
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 31668 478 31832 484
rect 32416 480 32444 575
rect 32640 598 32936 604
rect 34796 672 34848 678
rect 33836 620 34132 626
rect 33784 614 34132 620
rect 37280 672 37332 678
rect 34796 614 34848 620
rect 35990 640 36046 649
rect 33230 575 33286 584
rect 33600 604 33652 610
rect 32588 546 32640 552
rect 33244 542 33272 575
rect 33796 598 34132 614
rect 33600 546 33652 552
rect 33232 536 33284 542
rect 31680 462 31832 478
rect 32374 -960 32486 480
rect 33232 478 33284 484
rect 33612 480 33640 546
rect 34808 480 34836 614
rect 36096 610 36340 626
rect 38384 672 38436 678
rect 37332 620 37536 626
rect 37280 614 37536 620
rect 40684 672 40736 678
rect 38384 614 38436 620
rect 38474 640 38530 649
rect 35990 575 36046 584
rect 36084 604 36340 610
rect 34980 536 35032 542
rect 35032 484 35236 490
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 34980 478 35236 484
rect 36004 480 36032 575
rect 36136 598 36340 604
rect 37188 604 37240 610
rect 36084 546 36136 552
rect 37292 598 37536 614
rect 37188 546 37240 552
rect 37200 480 37228 546
rect 38396 480 38424 614
rect 38530 598 38640 626
rect 39316 598 39620 626
rect 42800 672 42852 678
rect 40684 614 40736 620
rect 38474 575 38530 584
rect 34992 462 35236 478
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39316 406 39344 598
rect 39592 480 39620 598
rect 39304 400 39356 406
rect 39304 342 39356 348
rect 39550 -960 39662 480
rect 39744 474 39896 490
rect 40696 480 40724 614
rect 40788 610 40940 626
rect 46664 672 46716 678
rect 42852 620 43148 626
rect 42800 614 43148 620
rect 40776 604 40940 610
rect 40828 598 40940 604
rect 41880 604 41932 610
rect 40776 546 40828 552
rect 42812 598 43148 614
rect 44008 610 44344 626
rect 43996 604 44344 610
rect 41880 546 41932 552
rect 44048 598 44344 604
rect 45112 598 45448 626
rect 46664 614 46716 620
rect 48504 672 48556 678
rect 48964 672 49016 678
rect 48556 620 48852 626
rect 48504 614 48852 620
rect 50804 672 50856 678
rect 48964 614 49016 620
rect 43996 546 44048 552
rect 41892 480 41920 546
rect 39744 468 39908 474
rect 39744 462 39856 468
rect 39856 410 39908 416
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 42156 400 42208 406
rect 42044 348 42156 354
rect 42044 342 42208 348
rect 42892 400 42944 406
rect 43046 354 43158 480
rect 42944 348 43158 354
rect 42892 342 43158 348
rect 42044 326 42196 342
rect 42904 326 43158 342
rect 43046 -960 43158 326
rect 44242 82 44354 480
rect 45112 406 45140 598
rect 46676 480 46704 614
rect 47860 604 47912 610
rect 48516 598 48852 614
rect 47860 546 47912 552
rect 47872 480 47900 546
rect 48976 480 49004 614
rect 49620 610 49956 626
rect 53748 672 53800 678
rect 52550 640 52606 649
rect 50856 620 51152 626
rect 50804 614 51152 620
rect 49608 604 49956 610
rect 49660 598 49956 604
rect 50160 604 50212 610
rect 49608 546 49660 552
rect 50816 598 51152 614
rect 51356 604 51408 610
rect 50160 546 50212 552
rect 53024 610 53360 626
rect 53748 614 53800 620
rect 55404 672 55456 678
rect 64328 672 64380 678
rect 56046 640 56102 649
rect 55456 620 55660 626
rect 55404 614 55660 620
rect 52550 575 52606 584
rect 53012 604 53360 610
rect 51356 546 51408 552
rect 50172 480 50200 546
rect 51368 480 51396 546
rect 51908 536 51960 542
rect 51960 484 52256 490
rect 45100 400 45152 406
rect 45100 342 45152 348
rect 44100 66 44354 82
rect 44088 60 44354 66
rect 44140 54 44354 60
rect 44088 2 44140 8
rect 44242 -960 44354 54
rect 45438 82 45550 480
rect 45744 128 45796 134
rect 45438 76 45744 82
rect 45438 70 45796 76
rect 45438 54 45784 70
rect 46216 66 46552 82
rect 46204 60 46552 66
rect 45438 -960 45550 54
rect 46256 54 46552 60
rect 46204 2 46256 8
rect 46634 -960 46746 480
rect 47400 128 47452 134
rect 47452 76 47748 82
rect 47400 70 47748 76
rect 47412 54 47748 70
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 51908 478 52256 484
rect 52564 480 52592 575
rect 53064 598 53360 604
rect 53012 546 53064 552
rect 53760 480 53788 614
rect 54944 604 54996 610
rect 55416 598 55660 614
rect 57610 640 57666 649
rect 56428 610 56764 626
rect 56046 575 56102 584
rect 56416 604 56764 610
rect 54944 546 54996 552
rect 54206 504 54262 513
rect 51920 462 52256 478
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54262 462 54556 490
rect 54956 480 54984 546
rect 56060 480 56088 575
rect 56468 598 56764 604
rect 56416 546 56468 552
rect 57256 564 57468 592
rect 58438 640 58494 649
rect 57666 598 57960 626
rect 57610 575 57666 584
rect 59818 640 59874 649
rect 58438 575 58494 584
rect 57256 480 57284 564
rect 57440 513 57468 564
rect 57426 504 57482 513
rect 54206 439 54262 448
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58452 480 58480 575
rect 59464 564 59676 592
rect 62026 640 62082 649
rect 59874 598 60168 626
rect 60832 604 60884 610
rect 59818 575 59874 584
rect 59464 513 59492 564
rect 58806 504 58862 513
rect 57426 439 57482 448
rect 58410 -960 58522 480
rect 59450 504 59506 513
rect 58862 462 59064 490
rect 58806 439 58862 448
rect 59648 480 59676 564
rect 63498 640 63554 649
rect 62132 610 62468 626
rect 62026 575 62082 584
rect 62120 604 62468 610
rect 60832 546 60884 552
rect 60844 480 60872 546
rect 61106 504 61162 513
rect 59450 439 59506 448
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61162 462 61364 490
rect 62040 480 62068 575
rect 62172 598 62468 604
rect 62120 546 62172 552
rect 63236 564 63448 592
rect 63554 598 63664 626
rect 64328 614 64380 620
rect 65616 672 65668 678
rect 66720 672 66772 678
rect 65668 620 65872 626
rect 65616 614 65872 620
rect 68008 672 68060 678
rect 66720 614 66772 620
rect 63498 575 63554 584
rect 63236 480 63264 564
rect 63420 490 63448 564
rect 63500 536 63552 542
rect 63420 484 63500 490
rect 61106 439 61162 448
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 63420 478 63552 484
rect 64340 480 64368 614
rect 65524 604 65576 610
rect 65628 598 65872 614
rect 65524 546 65576 552
rect 64512 536 64564 542
rect 64564 484 64768 490
rect 63420 462 63540 478
rect 64298 -960 64410 480
rect 64512 478 64768 484
rect 65536 480 65564 546
rect 66732 480 66760 614
rect 66824 610 67068 626
rect 66812 604 67068 610
rect 66864 598 67068 604
rect 67744 598 67956 626
rect 69112 672 69164 678
rect 68060 620 68172 626
rect 68008 614 68172 620
rect 70584 672 70636 678
rect 69112 614 69164 620
rect 70472 620 70584 626
rect 133236 672 133288 678
rect 70472 614 70636 620
rect 68020 598 68172 614
rect 66812 546 66864 552
rect 67744 542 67772 598
rect 67732 536 67784 542
rect 64524 462 64768 478
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67732 478 67784 484
rect 67928 480 67956 598
rect 69124 480 69152 614
rect 70308 604 70360 610
rect 70472 598 70624 614
rect 71240 610 71576 626
rect 71228 604 71576 610
rect 70308 546 70360 552
rect 71280 598 71576 604
rect 72344 598 72680 626
rect 73540 598 73876 626
rect 74644 598 74980 626
rect 76944 610 77280 626
rect 78048 610 78384 626
rect 79152 610 79488 626
rect 80348 610 80684 626
rect 81452 610 81788 626
rect 82740 610 82892 626
rect 76196 604 76248 610
rect 71228 546 71280 552
rect 69388 536 69440 542
rect 69276 484 69388 490
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 69276 478 69440 484
rect 70320 480 70348 546
rect 69276 462 69428 478
rect 70278 -960 70390 480
rect 71320 400 71372 406
rect 71474 354 71586 480
rect 72344 406 72372 598
rect 71372 348 71586 354
rect 71320 342 71586 348
rect 72332 400 72384 406
rect 72332 342 72384 348
rect 72424 400 72476 406
rect 72578 354 72690 480
rect 73540 406 73568 598
rect 72476 348 72690 354
rect 72424 342 72690 348
rect 73528 400 73580 406
rect 73528 342 73580 348
rect 73620 400 73672 406
rect 73774 354 73886 480
rect 74644 406 74672 598
rect 76196 546 76248 552
rect 76932 604 77280 610
rect 76984 598 77280 604
rect 77392 604 77444 610
rect 76932 546 76984 552
rect 77392 546 77444 552
rect 78036 604 78384 610
rect 78088 598 78384 604
rect 78588 604 78640 610
rect 78036 546 78088 552
rect 78588 546 78640 552
rect 79140 604 79488 610
rect 79192 598 79488 604
rect 79692 604 79744 610
rect 79140 546 79192 552
rect 79692 546 79744 552
rect 80336 604 80684 610
rect 80388 598 80684 604
rect 80888 604 80940 610
rect 80336 546 80388 552
rect 80888 546 80940 552
rect 81440 604 81788 610
rect 81492 598 81788 604
rect 82084 604 82136 610
rect 81440 546 81492 552
rect 82084 546 82136 552
rect 82728 604 82892 610
rect 82780 598 82892 604
rect 83292 598 83504 626
rect 82728 546 82780 552
rect 76208 480 76236 546
rect 77404 480 77432 546
rect 78600 480 78628 546
rect 79704 480 79732 546
rect 80900 480 80928 546
rect 82096 480 82124 546
rect 83292 480 83320 598
rect 83476 490 83504 598
rect 84488 598 85192 626
rect 85684 598 85896 626
rect 73672 348 73886 354
rect 73620 342 73886 348
rect 74632 400 74684 406
rect 74632 342 74684 348
rect 71332 326 71586 342
rect 72436 326 72690 342
rect 73632 326 73886 342
rect 71474 -960 71586 326
rect 72578 -960 72690 326
rect 73774 -960 73886 326
rect 74970 82 75082 480
rect 74970 54 76084 82
rect 74970 -960 75082 54
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 83476 462 84088 490
rect 84488 480 84516 598
rect 85684 480 85712 598
rect 85868 490 85896 598
rect 86880 598 87492 626
rect 87984 598 88596 626
rect 89180 598 89392 626
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 85868 462 86296 490
rect 86880 480 86908 598
rect 87984 480 88012 598
rect 89180 480 89208 598
rect 89364 490 89392 598
rect 90376 598 90896 626
rect 91572 598 92000 626
rect 92768 598 93196 626
rect 93964 598 94300 626
rect 95160 598 95404 626
rect 96264 598 96600 626
rect 97460 598 97704 626
rect 98656 598 98808 626
rect 99852 598 100004 626
rect 105616 598 105768 626
rect 106812 598 106964 626
rect 107916 598 108160 626
rect 109020 598 109356 626
rect 110216 598 110552 626
rect 111320 598 111656 626
rect 112424 598 112852 626
rect 113620 598 114048 626
rect 114724 598 115244 626
rect 115828 598 116440 626
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 89364 462 89792 490
rect 90376 480 90404 598
rect 91572 480 91600 598
rect 92768 480 92796 598
rect 93964 480 93992 598
rect 95160 480 95188 598
rect 96264 480 96292 598
rect 97460 480 97488 598
rect 98656 480 98684 598
rect 99852 480 99880 598
rect 105740 480 105768 598
rect 106936 480 106964 598
rect 108132 480 108160 598
rect 109328 480 109356 598
rect 110524 480 110552 598
rect 111628 480 111656 598
rect 112824 480 112852 598
rect 114020 480 114048 598
rect 115216 480 115244 598
rect 116412 480 116440 598
rect 117424 598 117636 626
rect 118128 598 118832 626
rect 119324 598 119936 626
rect 117424 490 117452 598
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117024 462 117452 490
rect 117608 480 117636 598
rect 118804 480 118832 598
rect 119908 480 119936 598
rect 120920 598 121132 626
rect 121532 610 121868 626
rect 121532 604 121880 610
rect 121532 598 121828 604
rect 120920 490 120948 598
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 120428 462 120948 490
rect 121104 480 121132 598
rect 121828 546 121880 552
rect 122288 604 122340 610
rect 122288 546 122340 552
rect 123312 598 123524 626
rect 123832 610 124168 626
rect 124936 610 125272 626
rect 126132 610 126468 626
rect 127236 610 127572 626
rect 128340 610 128676 626
rect 123832 604 124180 610
rect 123832 598 124128 604
rect 122300 480 122328 546
rect 123312 490 123340 598
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 122728 462 123340 490
rect 123496 480 123524 598
rect 124128 546 124180 552
rect 124680 604 124732 610
rect 124936 604 125284 610
rect 124936 598 125232 604
rect 124680 546 124732 552
rect 125232 546 125284 552
rect 125876 604 125928 610
rect 126132 604 126480 610
rect 126132 598 126428 604
rect 125876 546 125928 552
rect 126428 546 126480 552
rect 126980 604 127032 610
rect 127236 604 127584 610
rect 127236 598 127532 604
rect 126980 546 127032 552
rect 127532 546 127584 552
rect 128176 604 128228 610
rect 128340 604 128688 610
rect 128340 598 128636 604
rect 128176 546 128228 552
rect 128636 546 128688 552
rect 129372 604 129424 610
rect 130640 598 130976 626
rect 131744 598 132080 626
rect 132940 620 133236 626
rect 134156 672 134208 678
rect 132940 614 133288 620
rect 132940 598 133276 614
rect 133892 610 134044 626
rect 134156 614 134208 620
rect 136180 672 136232 678
rect 137652 672 137704 678
rect 136232 620 136344 626
rect 136180 614 136344 620
rect 133880 604 134044 610
rect 129372 546 129424 552
rect 124692 480 124720 546
rect 125888 480 125916 546
rect 126992 480 127020 546
rect 128188 480 128216 546
rect 129384 480 129412 546
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 129832 128 129884 134
rect 129536 76 129832 82
rect 129536 70 129884 76
rect 130292 128 130344 134
rect 130538 82 130650 480
rect 130948 406 130976 598
rect 130936 400 130988 406
rect 130936 342 130988 348
rect 131734 354 131846 480
rect 132052 406 132080 598
rect 133932 598 134044 604
rect 133880 546 133932 552
rect 134168 480 134196 614
rect 135260 604 135312 610
rect 136192 598 136344 614
rect 137448 610 137600 626
rect 138756 672 138808 678
rect 137652 614 137704 620
rect 138552 620 138756 626
rect 140044 672 140096 678
rect 138552 614 138808 620
rect 136456 604 136508 610
rect 135260 546 135312 552
rect 137448 604 137612 610
rect 137448 598 137560 604
rect 136456 546 136508 552
rect 137560 546 137612 552
rect 134984 536 135036 542
rect 135036 484 135148 490
rect 131948 400 132000 406
rect 131734 348 131948 354
rect 131734 342 132000 348
rect 132040 400 132092 406
rect 132040 342 132092 348
rect 132930 354 133042 480
rect 133144 400 133196 406
rect 132930 348 133144 354
rect 132930 342 133196 348
rect 130344 76 130650 82
rect 130292 70 130650 76
rect 129536 54 129872 70
rect 130304 54 130650 70
rect 130538 -960 130650 54
rect 131734 326 131988 342
rect 132930 326 133184 342
rect 131734 -960 131846 326
rect 132930 -960 133042 326
rect 134126 -960 134238 480
rect 134984 478 135148 484
rect 135272 480 135300 546
rect 136468 480 136496 546
rect 137664 480 137692 614
rect 138552 598 138796 614
rect 139748 610 139992 626
rect 151360 672 151412 678
rect 142066 640 142122 649
rect 140044 614 140096 620
rect 138848 604 138900 610
rect 139748 604 140004 610
rect 139748 598 139952 604
rect 138848 546 138900 552
rect 139952 546 140004 552
rect 138860 480 138888 546
rect 140056 480 140084 614
rect 141240 604 141292 610
rect 141956 598 142066 626
rect 143446 640 143502 649
rect 142066 575 142122 584
rect 142264 598 142476 626
rect 143152 598 143446 626
rect 141240 546 141292 552
rect 141056 536 141108 542
rect 140852 484 141056 490
rect 134996 462 135148 478
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 140852 478 141108 484
rect 141252 480 141280 546
rect 142068 536 142120 542
rect 142264 490 142292 598
rect 142120 484 142292 490
rect 140852 462 141096 478
rect 141210 -960 141322 480
rect 142068 478 142292 484
rect 142448 480 142476 598
rect 144734 640 144790 649
rect 143446 575 143502 584
rect 143552 598 143764 626
rect 144256 610 144592 626
rect 144256 604 144604 610
rect 144256 598 144552 604
rect 143552 480 143580 598
rect 143736 513 143764 598
rect 145746 640 145802 649
rect 145452 598 145746 626
rect 144734 575 144790 584
rect 147126 640 147182 649
rect 146556 610 146892 626
rect 145746 575 145802 584
rect 145932 604 145984 610
rect 144552 546 144604 552
rect 143722 504 143778 513
rect 142080 462 142292 478
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144748 480 144776 575
rect 146556 604 146904 610
rect 146556 598 146852 604
rect 145932 546 145984 552
rect 148966 640 149022 649
rect 147126 575 147182 584
rect 148324 604 148376 610
rect 146852 546 146904 552
rect 145944 480 145972 546
rect 147140 480 147168 575
rect 148856 598 148966 626
rect 150622 640 150678 649
rect 148966 575 149022 584
rect 149348 598 149560 626
rect 148324 546 148376 552
rect 147770 504 147826 513
rect 143722 439 143778 448
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 147660 462 147770 490
rect 148336 480 148364 546
rect 149348 513 149376 598
rect 149334 504 149390 513
rect 147770 439 147826 448
rect 148294 -960 148406 480
rect 149532 480 149560 598
rect 151064 620 151360 626
rect 153016 672 153068 678
rect 151064 614 151412 620
rect 151818 640 151874 649
rect 151064 598 151400 614
rect 150622 575 150678 584
rect 152260 610 152596 626
rect 153660 672 153712 678
rect 153016 614 153068 620
rect 153364 620 153660 626
rect 155408 672 155460 678
rect 153364 614 153712 620
rect 152260 604 152608 610
rect 152260 598 152556 604
rect 151818 575 151874 584
rect 150254 504 150310 513
rect 149334 439 149390 448
rect 149490 -960 149602 480
rect 149960 462 150254 490
rect 150636 480 150664 575
rect 151832 480 151860 575
rect 152556 546 152608 552
rect 153028 480 153056 614
rect 153364 598 153700 614
rect 154468 610 154804 626
rect 162768 672 162820 678
rect 155408 614 155460 620
rect 154212 604 154264 610
rect 154468 604 154816 610
rect 154468 598 154764 604
rect 154212 546 154264 552
rect 154764 546 154816 552
rect 154224 480 154252 546
rect 155420 480 155448 614
rect 156768 610 157104 626
rect 156604 604 156656 610
rect 156768 604 157116 610
rect 156768 598 157064 604
rect 156604 546 156656 552
rect 157872 598 158208 626
rect 157064 546 157116 552
rect 156616 480 156644 546
rect 158180 542 158208 598
rect 158904 604 158956 610
rect 160172 598 160508 626
rect 161276 610 161612 626
rect 162472 620 162768 626
rect 164884 672 164936 678
rect 164790 640 164846 649
rect 162472 614 162820 620
rect 161276 604 161624 610
rect 161276 598 161572 604
rect 158904 546 158956 552
rect 158168 536 158220 542
rect 150254 439 150310 448
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 155960 128 156012 134
rect 155664 76 155960 82
rect 155664 70 156012 76
rect 155664 54 156000 70
rect 156574 -960 156686 480
rect 157524 128 157576 134
rect 157770 82 157882 480
rect 158168 478 158220 484
rect 158916 480 158944 546
rect 159732 536 159784 542
rect 157576 76 157882 82
rect 157524 70 157882 76
rect 157536 54 157882 70
rect 157770 -960 157882 54
rect 158874 -960 158986 480
rect 159732 478 159784 484
rect 159744 354 159772 478
rect 160070 354 160182 480
rect 160480 406 160508 598
rect 162472 598 162808 614
rect 163688 604 163740 610
rect 161572 546 161624 552
rect 164680 598 164790 626
rect 166080 672 166132 678
rect 164884 614 164936 620
rect 164790 575 164846 584
rect 163688 546 163740 552
rect 159744 326 160182 354
rect 160468 400 160520 406
rect 160468 342 160520 348
rect 159364 128 159416 134
rect 159068 76 159364 82
rect 159068 70 159416 76
rect 159068 54 159404 70
rect 160070 -960 160182 326
rect 161266 82 161378 480
rect 162462 354 162574 480
rect 163424 474 163576 490
rect 163700 480 163728 546
rect 164896 480 164924 614
rect 165876 610 166028 626
rect 167092 672 167144 678
rect 166080 614 166132 620
rect 166980 620 167092 626
rect 169576 672 169628 678
rect 167366 640 167422 649
rect 166980 614 167144 620
rect 165876 604 166040 610
rect 165876 598 165988 604
rect 165988 546 166040 552
rect 166092 480 166120 614
rect 166980 598 167132 614
rect 167196 598 167366 626
rect 167196 480 167224 598
rect 169482 640 169538 649
rect 167366 575 167422 584
rect 168380 604 168432 610
rect 169280 598 169482 626
rect 180892 672 180944 678
rect 171966 640 172022 649
rect 169576 614 169628 620
rect 169482 575 169538 584
rect 168380 546 168432 552
rect 168392 480 168420 546
rect 169588 480 169616 614
rect 170384 610 170720 626
rect 170384 604 170732 610
rect 170384 598 170680 604
rect 170680 546 170732 552
rect 170784 598 170996 626
rect 170784 480 170812 598
rect 163412 468 163576 474
rect 163464 462 163576 468
rect 163412 410 163464 416
rect 162676 400 162728 406
rect 162462 348 162676 354
rect 162462 342 162728 348
rect 162462 326 162716 342
rect 161480 128 161532 134
rect 161266 76 161480 82
rect 161266 70 161532 76
rect 161266 54 161520 70
rect 161266 -960 161378 54
rect 162462 -960 162574 326
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168194 368 168250 377
rect 168084 326 168194 354
rect 168194 303 168250 312
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 170968 377 170996 598
rect 172978 640 173034 649
rect 172684 598 172978 626
rect 171966 575 172022 584
rect 175462 640 175518 649
rect 172978 575 173034 584
rect 173164 604 173216 610
rect 171980 480 172008 575
rect 173164 546 173216 552
rect 174096 598 174308 626
rect 173176 480 173204 546
rect 173898 504 173954 513
rect 170954 368 171010 377
rect 171690 368 171746 377
rect 171488 326 171690 354
rect 170954 303 171010 312
rect 171690 303 171746 312
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 173788 462 173898 490
rect 174096 490 174124 598
rect 173898 439 173954 448
rect 174004 462 174124 490
rect 174280 480 174308 598
rect 176382 640 176438 649
rect 176088 598 176382 626
rect 175462 575 175518 584
rect 179050 640 179106 649
rect 176382 575 176438 584
rect 176672 598 176884 626
rect 175476 480 175504 575
rect 176672 480 176700 598
rect 176856 513 176884 598
rect 177684 598 177896 626
rect 176842 504 176898 513
rect 174004 377 174032 462
rect 173990 368 174046 377
rect 173990 303 174046 312
rect 174238 -960 174350 480
rect 175186 368 175242 377
rect 174984 326 175186 354
rect 175186 303 175242 312
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177486 504 177542 513
rect 177192 462 177486 490
rect 176842 439 176898 448
rect 177486 439 177542 448
rect 177684 377 177712 598
rect 177868 480 177896 598
rect 180246 640 180302 649
rect 179492 610 179828 626
rect 179492 604 179840 610
rect 179492 598 179788 604
rect 179050 575 179106 584
rect 179064 480 179092 575
rect 180596 620 180892 626
rect 183744 672 183796 678
rect 182086 640 182142 649
rect 180596 614 180944 620
rect 180596 598 180932 614
rect 181272 598 181484 626
rect 181792 598 182086 626
rect 180246 575 180302 584
rect 179788 546 179840 552
rect 180260 480 180288 575
rect 177670 368 177726 377
rect 177670 303 177726 312
rect 177826 -960 177938 480
rect 178682 368 178738 377
rect 178388 326 178682 354
rect 178682 303 178738 312
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181272 377 181300 598
rect 181456 480 181484 598
rect 182896 610 183232 626
rect 186136 672 186188 678
rect 183744 614 183796 620
rect 184938 640 184994 649
rect 182086 575 182142 584
rect 182548 604 182600 610
rect 182896 604 183244 610
rect 182896 598 183192 604
rect 182548 546 182600 552
rect 183192 546 183244 552
rect 182560 480 182588 546
rect 183756 480 183784 614
rect 191104 672 191156 678
rect 186136 614 186188 620
rect 184938 575 184994 584
rect 184952 480 184980 575
rect 186148 480 186176 614
rect 187404 598 187740 626
rect 188600 598 188844 626
rect 189704 610 190040 626
rect 190808 620 191104 626
rect 194416 672 194468 678
rect 190808 614 191156 620
rect 189704 604 190052 610
rect 189704 598 190000 604
rect 186596 536 186648 542
rect 186300 484 186596 490
rect 181258 368 181314 377
rect 181258 303 181314 312
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184296 128 184348 134
rect 184000 76 184296 82
rect 184000 70 184348 76
rect 184000 54 184336 70
rect 184910 -960 185022 480
rect 185492 128 185544 134
rect 185196 76 185492 82
rect 185196 70 185544 76
rect 185196 54 185532 70
rect 186106 -960 186218 480
rect 186300 478 186648 484
rect 186300 462 186636 478
rect 187302 218 187414 480
rect 187712 474 187740 598
rect 187700 468 187752 474
rect 187700 410 187752 416
rect 186976 202 187414 218
rect 186964 196 187414 202
rect 187016 190 187414 196
rect 186964 138 187016 144
rect 187302 -960 187414 190
rect 188252 128 188304 134
rect 188498 82 188610 480
rect 188816 377 188844 598
rect 190808 598 191144 614
rect 192004 598 192340 626
rect 211620 672 211672 678
rect 196714 640 196770 649
rect 194416 614 194468 620
rect 190000 546 190052 552
rect 192312 542 192340 598
rect 193220 604 193272 610
rect 193220 546 193272 552
rect 189908 536 189960 542
rect 188802 368 188858 377
rect 188802 303 188858 312
rect 189694 354 189806 480
rect 189908 478 189960 484
rect 192300 536 192352 542
rect 189920 354 189948 478
rect 189694 326 189948 354
rect 190798 354 190910 480
rect 191012 468 191064 474
rect 191012 410 191064 416
rect 191024 354 191052 410
rect 190798 326 191052 354
rect 191994 354 192106 480
rect 192300 478 192352 484
rect 193232 480 193260 546
rect 192944 400 192996 406
rect 192206 368 192262 377
rect 191994 326 192206 354
rect 188304 76 188610 82
rect 188252 70 188610 76
rect 188264 54 188610 70
rect 188498 -960 188610 54
rect 189694 -960 189806 326
rect 190798 -960 190910 326
rect 191994 -960 192106 326
rect 192996 348 193108 354
rect 192944 342 193108 348
rect 192956 326 193108 342
rect 192206 303 192262 312
rect 193190 -960 193302 480
rect 194060 474 194212 490
rect 194428 480 194456 614
rect 195612 604 195664 610
rect 196512 598 196714 626
rect 200302 640 200358 649
rect 196714 575 196770 584
rect 196808 604 196860 610
rect 195612 546 195664 552
rect 196808 546 196860 552
rect 197912 604 197964 610
rect 197912 546 197964 552
rect 198936 598 199148 626
rect 195624 480 195652 546
rect 196820 480 196848 546
rect 197924 480 197952 546
rect 194048 468 194212 474
rect 194100 462 194212 468
rect 194048 410 194100 416
rect 194386 -960 194498 480
rect 195242 232 195298 241
rect 195298 190 195408 218
rect 195242 167 195298 176
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197726 368 197782 377
rect 197616 326 197726 354
rect 197726 303 197782 312
rect 197882 -960 197994 480
rect 198936 241 198964 598
rect 199120 480 199148 598
rect 200302 575 200358 584
rect 201498 640 201554 649
rect 203614 640 203670 649
rect 203320 598 203614 626
rect 201498 575 201554 584
rect 200316 480 200344 575
rect 201512 480 201540 575
rect 202524 564 202736 592
rect 207386 640 207442 649
rect 205620 610 205772 626
rect 205620 604 205784 610
rect 205620 598 205732 604
rect 203614 575 203670 584
rect 202418 504 202474 513
rect 198922 232 198978 241
rect 198922 167 198978 176
rect 198922 96 198978 105
rect 198812 54 198922 82
rect 198922 31 198978 40
rect 199078 -960 199190 480
rect 200026 368 200082 377
rect 199916 326 200026 354
rect 200026 303 200082 312
rect 200274 -960 200386 480
rect 201314 368 201370 377
rect 201112 326 201314 354
rect 201314 303 201370 312
rect 201470 -960 201582 480
rect 202216 462 202418 490
rect 202418 439 202474 448
rect 202524 105 202552 564
rect 202708 480 202736 564
rect 203720 564 203932 592
rect 202510 96 202566 105
rect 202510 31 202566 40
rect 202666 -960 202778 480
rect 203720 241 203748 564
rect 203904 480 203932 564
rect 204916 564 205128 592
rect 203706 232 203762 241
rect 203706 167 203762 176
rect 203862 -960 203974 480
rect 204916 377 204944 564
rect 205100 480 205128 564
rect 205732 546 205784 552
rect 206020 564 206232 592
rect 208214 640 208270 649
rect 207920 598 208214 626
rect 207386 575 207442 584
rect 208214 575 208270 584
rect 208398 640 208454 649
rect 209318 640 209374 649
rect 208398 575 208454 584
rect 208596 598 208808 626
rect 209024 598 209318 626
rect 206020 513 206048 564
rect 206006 504 206062 513
rect 204902 368 204958 377
rect 204902 303 204958 312
rect 204810 232 204866 241
rect 204516 190 204810 218
rect 204810 167 204866 176
rect 205058 -960 205170 480
rect 206204 480 206232 564
rect 206926 504 206982 513
rect 206006 439 206062 448
rect 206162 -960 206274 480
rect 206724 462 206926 490
rect 207400 480 207428 575
rect 208412 542 208440 575
rect 208400 536 208452 542
rect 206926 439 206982 448
rect 207358 -960 207470 480
rect 208400 478 208452 484
rect 208596 480 208624 598
rect 208554 -960 208666 480
rect 208780 241 208808 598
rect 210128 610 210464 626
rect 209318 575 209374 584
rect 209780 604 209832 610
rect 210128 604 210476 610
rect 210128 598 210424 604
rect 209780 546 209832 552
rect 210424 546 210476 552
rect 210804 598 211016 626
rect 211324 620 211620 626
rect 215668 672 215720 678
rect 211324 614 211672 620
rect 213366 640 213422 649
rect 211324 598 211660 614
rect 212172 604 212224 610
rect 209792 480 209820 546
rect 210804 513 210832 598
rect 210790 504 210846 513
rect 208766 232 208822 241
rect 208766 167 208822 176
rect 209750 -960 209862 480
rect 210988 480 211016 598
rect 220176 672 220228 678
rect 216126 640 216182 649
rect 215668 614 215720 620
rect 213366 575 213422 584
rect 214472 604 214524 610
rect 212172 546 212224 552
rect 212184 480 212212 546
rect 212724 536 212776 542
rect 212428 484 212724 490
rect 210790 439 210846 448
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 212428 478 212776 484
rect 213380 480 213408 575
rect 214472 546 214524 552
rect 214484 480 214512 546
rect 215680 480 215708 614
rect 215832 598 216126 626
rect 219990 640 220046 649
rect 216936 598 217272 626
rect 216126 575 216182 584
rect 216588 536 216640 542
rect 212428 462 212764 478
rect 213338 -960 213450 480
rect 213828 128 213880 134
rect 213532 76 213828 82
rect 213532 70 213880 76
rect 213532 54 213868 70
rect 214442 -960 214554 480
rect 214728 66 215064 82
rect 214728 60 215076 66
rect 214728 54 215024 60
rect 215024 2 215076 8
rect 215638 -960 215750 480
rect 216588 478 216640 484
rect 216600 218 216628 478
rect 216834 218 216946 480
rect 217244 406 217272 598
rect 217888 598 218054 626
rect 218132 598 218468 626
rect 219236 598 219572 626
rect 217232 400 217284 406
rect 217232 342 217284 348
rect 216600 190 216946 218
rect 216834 -960 216946 190
rect 217888 134 217916 598
rect 218026 480 218054 598
rect 218026 326 218142 480
rect 218440 474 218468 598
rect 219544 542 219572 598
rect 225328 672 225380 678
rect 221830 640 221886 649
rect 220228 620 220340 626
rect 220176 614 220340 620
rect 220188 598 220340 614
rect 220452 604 220504 610
rect 219990 575 219992 584
rect 220044 575 220046 584
rect 219992 546 220044 552
rect 221536 598 221830 626
rect 224940 610 225092 626
rect 225156 620 225328 626
rect 226156 672 226208 678
rect 225156 614 225380 620
rect 226044 620 226156 626
rect 231032 672 231084 678
rect 226044 614 226208 620
rect 226338 640 226394 649
rect 223948 604 224000 610
rect 221830 575 221886 584
rect 220452 546 220504 552
rect 222764 564 222976 592
rect 219532 536 219584 542
rect 218428 468 218480 474
rect 218428 410 218480 416
rect 217876 128 217928 134
rect 217876 70 217928 76
rect 218030 -960 218142 326
rect 219226 82 219338 480
rect 219532 478 219584 484
rect 220464 480 220492 546
rect 222764 480 222792 564
rect 219226 66 219480 82
rect 219226 60 219492 66
rect 219226 54 219440 60
rect 219226 -960 219338 54
rect 219440 2 219492 8
rect 220422 -960 220534 480
rect 221526 354 221638 480
rect 221740 400 221792 406
rect 221526 348 221740 354
rect 221526 342 221792 348
rect 222476 400 222528 406
rect 222528 348 222640 354
rect 222476 342 222640 348
rect 221526 326 221780 342
rect 222488 326 222640 342
rect 221526 -960 221638 326
rect 222722 -960 222834 480
rect 222948 474 222976 564
rect 224940 604 225104 610
rect 224940 598 225052 604
rect 223948 546 224000 552
rect 225052 546 225104 552
rect 225156 598 225368 614
rect 226044 598 226196 614
rect 223578 504 223634 513
rect 222936 468 222988 474
rect 223634 462 223744 490
rect 223960 480 223988 546
rect 225156 480 225184 598
rect 228730 640 228786 649
rect 226338 575 226394 584
rect 227364 598 227576 626
rect 226352 480 226380 575
rect 227364 542 227392 598
rect 227352 536 227404 542
rect 223578 439 223634 448
rect 222936 410 222988 416
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227352 478 227404 484
rect 227548 480 227576 598
rect 230938 640 230994 649
rect 228730 575 228786 584
rect 229836 604 229888 610
rect 228744 480 228772 575
rect 230644 598 230938 626
rect 234620 672 234672 678
rect 231032 614 231084 620
rect 230938 575 230994 584
rect 229836 546 229888 552
rect 229652 536 229704 542
rect 229448 484 229652 490
rect 227352 264 227404 270
rect 227148 212 227352 218
rect 227148 206 227404 212
rect 227148 190 227392 206
rect 227506 -960 227618 480
rect 228344 202 228588 218
rect 228344 196 228600 202
rect 228344 190 228548 196
rect 228548 138 228600 144
rect 228702 -960 228814 480
rect 229448 478 229704 484
rect 229848 480 229876 546
rect 231044 480 231072 614
rect 231748 610 231900 626
rect 231748 604 231912 610
rect 231748 598 231860 604
rect 231860 546 231912 552
rect 232056 598 232268 626
rect 229448 462 229692 478
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232056 270 232084 598
rect 232240 480 232268 598
rect 233252 598 233464 626
rect 235448 672 235500 678
rect 234620 614 234672 620
rect 235152 620 235448 626
rect 237748 672 237800 678
rect 235152 614 235500 620
rect 235814 640 235870 649
rect 233148 536 233200 542
rect 232852 484 233148 490
rect 232044 264 232096 270
rect 232044 206 232096 212
rect 232198 -960 232310 480
rect 232852 478 233200 484
rect 232852 462 233188 478
rect 233252 270 233280 598
rect 233436 480 233464 598
rect 233240 264 233292 270
rect 233240 206 233292 212
rect 233394 -960 233506 480
rect 234048 474 234384 490
rect 234632 480 234660 614
rect 235152 598 235488 614
rect 237452 620 237748 626
rect 242900 672 242952 678
rect 239954 640 240010 649
rect 237452 614 237800 620
rect 235814 575 235870 584
rect 237012 604 237064 610
rect 235828 480 235856 575
rect 237452 598 237788 614
rect 238116 604 238168 610
rect 237012 546 237064 552
rect 238116 546 238168 552
rect 239312 604 239364 610
rect 239660 598 239954 626
rect 240856 610 241192 626
rect 246764 672 246816 678
rect 245198 640 245254 649
rect 242900 614 242952 620
rect 239954 575 240010 584
rect 240508 604 240560 610
rect 239312 546 239364 552
rect 240856 604 241204 610
rect 240856 598 241152 604
rect 240508 546 240560 552
rect 241152 546 241204 552
rect 241532 564 241744 592
rect 237024 480 237052 546
rect 238128 480 238156 546
rect 238852 536 238904 542
rect 238556 484 238852 490
rect 234048 468 234396 474
rect 234048 462 234344 468
rect 234344 410 234396 416
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236256 202 236592 218
rect 236256 196 236604 202
rect 236256 190 236552 196
rect 236552 138 236604 144
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 238556 478 238904 484
rect 239324 480 239352 546
rect 240520 480 240548 546
rect 238556 462 238892 478
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241532 354 241560 564
rect 241716 480 241744 564
rect 242912 480 242940 614
rect 243924 598 244136 626
rect 243924 542 243952 598
rect 243912 536 243964 542
rect 241440 326 241560 354
rect 241440 202 241468 326
rect 241428 196 241480 202
rect 241428 138 241480 144
rect 241674 -960 241786 480
rect 242256 400 242308 406
rect 241960 348 242256 354
rect 241960 342 242308 348
rect 241960 326 242296 342
rect 242870 -960 242982 480
rect 243064 474 243400 490
rect 243912 478 243964 484
rect 244108 480 244136 598
rect 246468 620 246764 626
rect 247960 672 248012 678
rect 246468 614 246816 620
rect 247664 620 247960 626
rect 253480 672 253532 678
rect 249062 640 249118 649
rect 247664 614 248012 620
rect 245198 575 245254 584
rect 246028 604 246080 610
rect 243064 468 243412 474
rect 243064 462 243360 468
rect 243360 410 243412 416
rect 244066 -960 244178 480
rect 244260 474 244596 490
rect 245212 480 245240 575
rect 246468 598 246804 614
rect 247664 598 248000 614
rect 248768 598 249062 626
rect 253276 610 253428 626
rect 257252 672 257304 678
rect 254674 640 254730 649
rect 253480 614 253532 620
rect 249062 575 249118 584
rect 249984 604 250036 610
rect 246028 546 246080 552
rect 249984 546 250036 552
rect 251180 604 251232 610
rect 251180 546 251232 552
rect 252376 604 252428 610
rect 253276 604 253440 610
rect 253276 598 253388 604
rect 252376 546 252428 552
rect 253388 546 253440 552
rect 244260 468 244608 474
rect 244260 462 244556 468
rect 244556 410 244608 416
rect 245170 -960 245282 480
rect 246040 354 246068 546
rect 248972 536 249024 542
rect 246366 354 246478 480
rect 245364 338 245700 354
rect 245364 332 245712 338
rect 245364 326 245660 332
rect 246040 326 246478 354
rect 247316 400 247368 406
rect 247562 354 247674 480
rect 247368 348 247674 354
rect 247316 342 247674 348
rect 247328 326 247674 342
rect 245660 274 245712 280
rect 246366 -960 246478 326
rect 247562 -960 247674 326
rect 248758 354 248870 480
rect 248972 478 249024 484
rect 249706 504 249762 513
rect 248984 354 249012 478
rect 249762 462 249872 490
rect 249996 480 250024 546
rect 251192 480 251220 546
rect 252388 480 252416 546
rect 253492 480 253520 614
rect 254472 610 254624 626
rect 254472 604 254636 610
rect 254472 598 254584 604
rect 254674 575 254730 584
rect 255870 640 255926 649
rect 255870 575 255926 584
rect 256896 598 257108 626
rect 257252 614 257304 620
rect 258264 672 258316 678
rect 260656 672 260708 678
rect 258264 614 258316 620
rect 254584 546 254636 552
rect 254688 480 254716 575
rect 255884 480 255912 575
rect 249706 439 249762 448
rect 248758 326 249012 354
rect 248758 -960 248870 326
rect 249954 -960 250066 480
rect 250904 264 250956 270
rect 250956 212 251068 218
rect 250904 206 251068 212
rect 250916 190 251068 206
rect 251150 -960 251262 480
rect 252020 338 252172 354
rect 252008 332 252172 338
rect 252060 326 252172 332
rect 252008 274 252060 280
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255688 264 255740 270
rect 255576 212 255688 218
rect 255576 206 255740 212
rect 255576 190 255728 206
rect 255842 -960 255954 480
rect 256896 474 256924 598
rect 257080 480 257108 598
rect 256884 468 256936 474
rect 256884 410 256936 416
rect 256772 66 256924 82
rect 256772 60 256936 66
rect 256772 54 256884 60
rect 256884 2 256936 8
rect 257038 -960 257150 480
rect 257264 338 257292 614
rect 257876 474 258028 490
rect 258276 480 258304 614
rect 260176 610 260512 626
rect 262680 672 262732 678
rect 260656 614 260708 620
rect 262384 620 262680 626
rect 268844 672 268896 678
rect 262384 614 262732 620
rect 263138 640 263194 649
rect 259460 604 259512 610
rect 260176 604 260524 610
rect 260176 598 260472 604
rect 259460 546 259512 552
rect 260472 546 260524 552
rect 257876 468 258040 474
rect 257876 462 257988 468
rect 257988 410 258040 416
rect 257252 332 257304 338
rect 257252 274 257304 280
rect 258234 -960 258346 480
rect 258980 474 259316 490
rect 259472 480 259500 546
rect 260668 480 260696 614
rect 262384 598 262720 614
rect 261772 564 261984 592
rect 261576 536 261628 542
rect 261280 484 261576 490
rect 258980 468 259328 474
rect 258980 462 259276 468
rect 259276 410 259328 416
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261280 478 261628 484
rect 261772 480 261800 564
rect 261280 462 261616 478
rect 261730 -960 261842 480
rect 261956 270 261984 564
rect 262784 564 262996 592
rect 263138 575 263194 584
rect 264150 640 264206 649
rect 267278 640 267334 649
rect 266544 604 266596 610
rect 264150 575 264206 584
rect 261944 264 261996 270
rect 261944 206 261996 212
rect 262784 66 262812 564
rect 262968 480 262996 564
rect 262772 60 262824 66
rect 262772 2 262824 8
rect 262926 -960 263038 480
rect 263152 406 263180 575
rect 264164 480 264192 575
rect 265176 564 265388 592
rect 265176 490 265204 564
rect 263140 400 263192 406
rect 263140 342 263192 348
rect 263692 264 263744 270
rect 263580 212 263692 218
rect 263580 206 263744 212
rect 263580 190 263732 206
rect 264122 -960 264234 480
rect 264992 474 265204 490
rect 265360 480 265388 564
rect 266984 598 267278 626
rect 269488 672 269540 678
rect 268844 614 268896 620
rect 269192 620 269488 626
rect 276204 672 276256 678
rect 273626 640 273682 649
rect 269192 614 269540 620
rect 267278 575 267334 584
rect 267740 604 267792 610
rect 266544 546 266596 552
rect 267740 546 267792 552
rect 264980 468 265204 474
rect 265032 462 265204 468
rect 264980 410 265032 416
rect 264684 66 264928 82
rect 264684 60 264940 66
rect 264684 54 264888 60
rect 264888 2 264940 8
rect 265318 -960 265430 480
rect 265788 474 266124 490
rect 266556 480 266584 546
rect 267752 480 267780 546
rect 268384 536 268436 542
rect 268088 484 268384 490
rect 265788 468 266136 474
rect 265788 462 266084 468
rect 266084 410 266136 416
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268088 478 268436 484
rect 268856 480 268884 614
rect 269192 598 269528 614
rect 270040 604 270092 610
rect 270040 546 270092 552
rect 271064 598 271276 626
rect 271492 610 271828 626
rect 271492 604 271840 610
rect 271492 598 271788 604
rect 270052 480 270080 546
rect 268088 462 268424 478
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 270684 400 270736 406
rect 270388 348 270684 354
rect 270388 342 270736 348
rect 270388 326 270724 342
rect 271064 66 271092 598
rect 271248 480 271276 598
rect 271788 546 271840 552
rect 272168 564 272472 592
rect 275190 640 275246 649
rect 274896 598 275190 626
rect 273626 575 273682 584
rect 275190 575 275246 584
rect 275848 598 276000 626
rect 279240 672 279292 678
rect 276204 614 276256 620
rect 271052 60 271104 66
rect 271052 2 271104 8
rect 271206 -960 271318 480
rect 272168 474 272196 564
rect 272444 480 272472 564
rect 273640 480 273668 575
rect 274548 536 274600 542
rect 272156 468 272208 474
rect 272156 410 272208 416
rect 272402 -960 272514 480
rect 272892 264 272944 270
rect 272596 212 272892 218
rect 272596 206 272944 212
rect 272596 190 272932 206
rect 273598 -960 273710 480
rect 274548 478 274600 484
rect 274560 354 274588 478
rect 274794 354 274906 480
rect 274560 326 274906 354
rect 275848 338 275876 598
rect 273792 202 274128 218
rect 273792 196 274140 202
rect 273792 190 274088 196
rect 274088 138 274140 144
rect 274794 -960 274906 326
rect 275836 332 275888 338
rect 275836 274 275888 280
rect 275990 218 276102 480
rect 276216 218 276244 614
rect 277196 610 277532 626
rect 277196 604 277544 610
rect 277196 598 277492 604
rect 278300 598 278636 626
rect 279516 672 279568 678
rect 279292 620 279404 626
rect 279240 614 279404 620
rect 284300 672 284352 678
rect 279516 614 279568 620
rect 281906 640 281962 649
rect 279252 598 279404 614
rect 277492 546 277544 552
rect 278608 542 278636 598
rect 278504 536 278556 542
rect 276756 400 276808 406
rect 277094 354 277206 480
rect 276808 348 277206 354
rect 276756 342 277206 348
rect 276768 326 277206 342
rect 275990 190 276244 218
rect 275990 -960 276102 190
rect 277094 -960 277206 326
rect 278290 354 278402 480
rect 278504 478 278556 484
rect 278596 536 278648 542
rect 278596 478 278648 484
rect 279528 480 279556 614
rect 280712 604 280764 610
rect 284300 614 284352 620
rect 286600 672 286652 678
rect 291108 672 291160 678
rect 286600 614 286652 620
rect 287058 640 287114 649
rect 281906 575 281962 584
rect 283104 604 283156 610
rect 280712 546 280764 552
rect 278516 354 278544 478
rect 278290 326 278544 354
rect 278290 -960 278402 326
rect 279486 -960 279598 480
rect 280448 474 280600 490
rect 280724 480 280752 546
rect 281920 480 281948 575
rect 283104 546 283156 552
rect 283116 480 283144 546
rect 284312 480 284340 614
rect 285404 604 285456 610
rect 285404 546 285456 552
rect 285218 504 285274 513
rect 280436 468 280600 474
rect 280488 462 280600 468
rect 280436 410 280488 416
rect 280682 -960 280794 480
rect 281540 400 281592 406
rect 281592 348 281704 354
rect 281540 342 281704 348
rect 281552 326 281704 342
rect 281878 -960 281990 480
rect 282808 202 282960 218
rect 282808 196 282972 202
rect 282808 190 282920 196
rect 282920 138 282972 144
rect 283074 -960 283186 480
rect 284004 338 284156 354
rect 284004 332 284168 338
rect 284004 326 284116 332
rect 284116 274 284168 280
rect 284270 -960 284382 480
rect 285108 462 285218 490
rect 285416 480 285444 546
rect 286416 536 286468 542
rect 286304 484 286416 490
rect 285218 439 285274 448
rect 285374 -960 285486 480
rect 286304 478 286468 484
rect 286612 480 286640 614
rect 288990 640 289046 649
rect 287058 575 287114 584
rect 287624 598 287836 626
rect 288512 610 288848 626
rect 288512 604 288860 610
rect 288512 598 288808 604
rect 286304 462 286456 478
rect 286570 -960 286682 480
rect 287072 406 287100 575
rect 287624 490 287652 598
rect 287532 474 287652 490
rect 287808 480 287836 598
rect 288990 575 289046 584
rect 290016 598 290228 626
rect 290812 620 291108 626
rect 298468 672 298520 678
rect 292578 640 292634 649
rect 290812 614 291160 620
rect 290812 598 291148 614
rect 291212 598 291424 626
rect 288808 546 288860 552
rect 289004 480 289032 575
rect 287520 468 287652 474
rect 287572 462 287652 468
rect 287520 410 287572 416
rect 287060 400 287112 406
rect 287612 400 287664 406
rect 287060 342 287112 348
rect 287408 348 287612 354
rect 287408 342 287664 348
rect 287408 326 287652 342
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 289708 474 289860 490
rect 289708 468 289872 474
rect 289708 462 289820 468
rect 289820 410 289872 416
rect 290016 202 290044 598
rect 290200 480 290228 598
rect 290004 196 290056 202
rect 290004 138 290056 144
rect 290158 -960 290270 480
rect 291212 338 291240 598
rect 291396 480 291424 598
rect 293866 640 293922 649
rect 292578 575 292634 584
rect 293512 598 293724 626
rect 292592 480 292620 575
rect 293316 536 293368 542
rect 293512 490 293540 598
rect 293368 484 293540 490
rect 291200 332 291252 338
rect 291200 274 291252 280
rect 291354 -960 291466 480
rect 291916 202 292252 218
rect 291916 196 292264 202
rect 291916 190 292212 196
rect 292212 138 292264 144
rect 292550 -960 292662 480
rect 293316 478 293540 484
rect 293696 480 293724 598
rect 293866 575 293922 584
rect 294878 640 294934 649
rect 295614 640 295670 649
rect 295320 598 295614 626
rect 294878 575 294934 584
rect 304724 672 304776 678
rect 303158 640 303214 649
rect 298468 614 298520 620
rect 295614 575 295670 584
rect 296076 604 296128 610
rect 293328 462 293540 478
rect 293112 66 293448 82
rect 293112 60 293460 66
rect 293112 54 293408 60
rect 293408 2 293460 8
rect 293654 -960 293766 480
rect 293880 406 293908 575
rect 294892 480 294920 575
rect 296076 546 296128 552
rect 297272 604 297324 610
rect 297272 546 297324 552
rect 296088 480 296116 546
rect 296812 536 296864 542
rect 296516 484 296812 490
rect 293868 400 293920 406
rect 294512 400 294564 406
rect 293868 342 293920 348
rect 294216 348 294512 354
rect 294216 342 294564 348
rect 294216 326 294552 342
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 296516 478 296864 484
rect 297284 480 297312 546
rect 298480 480 298508 614
rect 299492 598 299704 626
rect 299920 610 300256 626
rect 299920 604 300268 610
rect 299920 598 300216 604
rect 299492 490 299520 598
rect 296516 462 296852 478
rect 297242 -960 297354 480
rect 297916 264 297968 270
rect 297620 212 297916 218
rect 297620 206 297968 212
rect 297620 190 297956 206
rect 298438 -960 298550 480
rect 299400 462 299520 490
rect 299676 480 299704 598
rect 300216 546 300268 552
rect 300596 598 300808 626
rect 298724 338 299060 354
rect 298724 332 299072 338
rect 298724 326 299020 332
rect 299020 274 299072 280
rect 299400 202 299428 462
rect 299388 196 299440 202
rect 299388 138 299440 144
rect 299634 -960 299746 480
rect 300596 354 300624 598
rect 300780 480 300808 598
rect 301792 564 302004 592
rect 304428 620 304724 626
rect 307668 672 307720 678
rect 305826 640 305882 649
rect 304428 614 304776 620
rect 304428 598 304764 614
rect 305532 598 305826 626
rect 303158 575 303214 584
rect 306728 598 307064 626
rect 309968 672 310020 678
rect 307720 620 307832 626
rect 307668 614 307832 620
rect 312636 672 312688 678
rect 310020 620 310132 626
rect 309968 614 310132 620
rect 315948 672 316000 678
rect 312636 614 312688 620
rect 313830 640 313886 649
rect 307680 598 307832 614
rect 307944 604 307996 610
rect 305826 575 305882 584
rect 300504 326 300624 354
rect 300504 66 300532 326
rect 300492 60 300544 66
rect 300492 2 300544 8
rect 300738 -960 300850 480
rect 301024 474 301360 490
rect 301024 468 301372 474
rect 301024 462 301320 468
rect 301320 410 301372 416
rect 301792 406 301820 564
rect 301976 480 302004 564
rect 303172 480 303200 575
rect 303988 536 304040 542
rect 307036 513 307064 598
rect 307944 546 307996 552
rect 309048 604 309100 610
rect 309980 598 310132 614
rect 310244 604 310296 610
rect 309048 546 309100 552
rect 310244 546 310296 552
rect 311440 604 311492 610
rect 311440 546 311492 552
rect 301780 400 301832 406
rect 301780 342 301832 348
rect 301934 -960 302046 480
rect 302128 338 302464 354
rect 302128 332 302476 338
rect 302128 326 302424 332
rect 302424 274 302476 280
rect 303130 -960 303242 480
rect 303988 478 304040 484
rect 307022 504 307078 513
rect 304000 354 304028 478
rect 304326 354 304438 480
rect 304000 326 304438 354
rect 303324 66 303660 82
rect 303324 60 303672 66
rect 303324 54 303620 60
rect 303620 2 303672 8
rect 304326 -960 304438 326
rect 305522 218 305634 480
rect 306718 354 306830 480
rect 307956 480 307984 546
rect 309060 480 309088 546
rect 310256 480 310284 546
rect 311452 480 311480 546
rect 312452 536 312504 542
rect 312340 484 312452 490
rect 307022 439 307078 448
rect 306932 400 306984 406
rect 306718 348 306932 354
rect 306718 342 306984 348
rect 306718 326 306972 342
rect 305736 264 305788 270
rect 305522 212 305736 218
rect 305522 206 305788 212
rect 305522 190 305776 206
rect 305522 -960 305634 190
rect 306718 -960 306830 326
rect 307914 -960 308026 480
rect 308772 264 308824 270
rect 308824 212 308936 218
rect 308772 206 308936 212
rect 308784 190 308936 206
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311084 66 311236 82
rect 311072 60 311236 66
rect 311124 54 311236 60
rect 311072 2 311124 8
rect 311410 -960 311522 480
rect 312340 478 312504 484
rect 312648 480 312676 614
rect 313830 575 313886 584
rect 315026 640 315082 649
rect 315836 620 315948 626
rect 319720 672 319772 678
rect 315836 614 316000 620
rect 316406 640 316462 649
rect 315836 598 315988 614
rect 316224 604 316276 610
rect 315026 575 315082 584
rect 313844 480 313872 575
rect 315040 480 315068 575
rect 316406 575 316462 584
rect 317326 640 317382 649
rect 320916 672 320968 678
rect 319720 614 319772 620
rect 317326 575 317382 584
rect 316224 546 316276 552
rect 316236 480 316264 546
rect 312340 462 312492 478
rect 312606 -960 312718 480
rect 313536 338 313688 354
rect 313536 332 313700 338
rect 313536 326 313648 332
rect 313648 274 313700 280
rect 313802 -960 313914 480
rect 314752 400 314804 406
rect 314640 348 314752 354
rect 314640 342 314804 348
rect 314640 326 314792 342
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 316420 270 316448 575
rect 317144 536 317196 542
rect 316940 484 317144 490
rect 316940 478 317196 484
rect 317340 480 317368 575
rect 318352 564 318564 592
rect 318352 490 318380 564
rect 316940 462 317184 478
rect 316408 264 316460 270
rect 316408 206 316460 212
rect 317298 -960 317410 480
rect 318168 474 318380 490
rect 318536 480 318564 564
rect 318156 468 318380 474
rect 318208 462 318380 468
rect 318156 410 318208 416
rect 318340 400 318392 406
rect 318044 348 318340 354
rect 318044 342 318392 348
rect 318044 326 318380 342
rect 318494 -960 318606 480
rect 319240 474 319576 490
rect 319732 480 319760 614
rect 320344 610 320680 626
rect 323308 672 323360 678
rect 320916 614 320968 620
rect 320344 604 320692 610
rect 320344 598 320640 604
rect 320640 546 320692 552
rect 320928 480 320956 614
rect 321940 598 322152 626
rect 323308 614 323360 620
rect 324412 672 324464 678
rect 329196 672 329248 678
rect 324412 614 324464 620
rect 321940 490 321968 598
rect 319240 468 319588 474
rect 319240 462 319536 468
rect 319536 410 319588 416
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 321848 462 321968 490
rect 322124 480 322152 598
rect 323320 480 323348 614
rect 324424 480 324452 614
rect 325608 604 325660 610
rect 325608 546 325660 552
rect 326632 598 326844 626
rect 335360 672 335412 678
rect 329196 614 329248 620
rect 325620 480 325648 546
rect 326342 504 326398 513
rect 321448 338 321600 354
rect 321448 332 321612 338
rect 321448 326 321560 332
rect 321560 274 321612 280
rect 321848 202 321876 462
rect 321836 196 321888 202
rect 321836 138 321888 144
rect 322082 -960 322194 480
rect 322644 66 322888 82
rect 322644 60 322900 66
rect 322644 54 322848 60
rect 322848 2 322900 8
rect 323278 -960 323390 480
rect 323748 202 324084 218
rect 323748 196 324096 202
rect 323748 190 324044 196
rect 324044 138 324096 144
rect 324382 -960 324494 480
rect 324852 202 325188 218
rect 324852 196 325200 202
rect 324852 190 325148 196
rect 325148 138 325200 144
rect 325578 -960 325690 480
rect 326048 462 326342 490
rect 326342 439 326398 448
rect 326632 406 326660 598
rect 326816 480 326844 598
rect 328000 604 328052 610
rect 328000 546 328052 552
rect 328012 480 328040 546
rect 329208 480 329236 614
rect 331660 598 331996 626
rect 333960 610 334296 626
rect 335064 620 335360 626
rect 344560 672 344612 678
rect 336554 640 336610 649
rect 335064 614 335412 620
rect 330220 564 330432 592
rect 330220 490 330248 564
rect 326620 400 326672 406
rect 326620 342 326672 348
rect 326774 -960 326886 480
rect 327448 400 327500 406
rect 327152 348 327448 354
rect 327152 342 327500 348
rect 327152 326 327488 342
rect 327970 -960 328082 480
rect 328552 264 328604 270
rect 328256 212 328552 218
rect 328256 206 328604 212
rect 328256 190 328592 206
rect 329166 -960 329278 480
rect 330128 462 330248 490
rect 330404 480 330432 564
rect 330852 536 330904 542
rect 330556 484 330852 490
rect 330128 338 330156 462
rect 330116 332 330168 338
rect 330116 274 330168 280
rect 329748 128 329800 134
rect 329452 76 329748 82
rect 329452 70 329800 76
rect 329452 54 329788 70
rect 330362 -960 330474 480
rect 330556 478 330904 484
rect 330556 462 330892 478
rect 331558 82 331670 480
rect 331968 474 331996 598
rect 332692 604 332744 610
rect 333960 604 334308 610
rect 333960 598 334256 604
rect 332692 546 332744 552
rect 335064 598 335400 614
rect 336260 598 336554 626
rect 343454 640 343510 649
rect 341812 610 341964 626
rect 336554 575 336610 584
rect 337476 604 337528 610
rect 334256 546 334308 552
rect 337476 546 337528 552
rect 338672 604 338724 610
rect 338672 546 338724 552
rect 339868 604 339920 610
rect 339868 546 339920 552
rect 340972 604 341024 610
rect 340972 546 341024 552
rect 341800 604 341964 610
rect 341852 598 341964 604
rect 342168 604 342220 610
rect 341800 546 341852 552
rect 342168 546 342220 552
rect 343364 604 343416 610
rect 347688 672 347740 678
rect 344560 614 344612 620
rect 347576 620 347688 626
rect 357532 672 357584 678
rect 347576 614 347740 620
rect 343454 575 343456 584
rect 343364 546 343416 552
rect 343508 575 343510 584
rect 343456 546 343508 552
rect 332704 480 332732 546
rect 335266 504 335322 513
rect 331956 468 332008 474
rect 331956 410 332008 416
rect 331232 66 331670 82
rect 331220 60 331670 66
rect 331272 54 331670 60
rect 331220 2 331272 8
rect 331558 -960 331670 54
rect 332662 -960 332774 480
rect 333152 400 333204 406
rect 332856 348 333152 354
rect 332856 342 333204 348
rect 332856 326 333192 342
rect 333858 218 333970 480
rect 333624 202 333970 218
rect 333612 196 333970 202
rect 333664 190 333970 196
rect 333612 138 333664 144
rect 333858 -960 333970 190
rect 335054 218 335166 480
rect 337488 480 337516 546
rect 338684 480 338712 546
rect 339880 480 339908 546
rect 340984 480 341012 546
rect 342180 480 342208 546
rect 335266 439 335322 448
rect 335280 218 335308 439
rect 335054 190 335308 218
rect 336250 354 336362 480
rect 336250 338 336504 354
rect 337212 338 337364 354
rect 336250 332 336516 338
rect 336250 326 336464 332
rect 335054 -960 335166 190
rect 336250 -960 336362 326
rect 336464 274 336516 280
rect 337200 332 337364 338
rect 337252 326 337364 332
rect 337200 274 337252 280
rect 337446 -960 337558 480
rect 338316 202 338468 218
rect 338304 196 338468 202
rect 338356 190 338468 196
rect 338304 138 338356 144
rect 338642 -960 338754 480
rect 339500 128 339552 134
rect 339552 76 339664 82
rect 339500 70 339664 76
rect 339512 54 339664 70
rect 339838 -960 339950 480
rect 340604 400 340656 406
rect 340656 348 340768 354
rect 340604 342 340768 348
rect 340616 326 340768 342
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343068 474 343220 490
rect 343376 480 343404 546
rect 344374 504 344430 513
rect 343068 468 343232 474
rect 343068 462 343180 468
rect 343180 410 343232 416
rect 343334 -960 343446 480
rect 344172 462 344374 490
rect 344572 480 344600 614
rect 345756 604 345808 610
rect 347576 598 347728 614
rect 351472 598 351684 626
rect 356684 610 357020 626
rect 367008 672 367060 678
rect 364890 640 364946 649
rect 357532 614 357584 620
rect 345756 546 345808 552
rect 346780 564 346992 592
rect 345768 480 345796 546
rect 346780 490 346808 564
rect 344374 439 344430 448
rect 344530 -960 344642 480
rect 345368 202 345612 218
rect 345368 196 345624 202
rect 345368 190 345572 196
rect 345572 138 345624 144
rect 345726 -960 345838 480
rect 346688 462 346808 490
rect 346964 480 346992 564
rect 347884 564 348096 592
rect 347688 536 347740 542
rect 347686 504 347688 513
rect 347740 504 347742 513
rect 346688 338 346716 462
rect 346676 332 346728 338
rect 346676 274 346728 280
rect 346768 264 346820 270
rect 346472 212 346768 218
rect 346472 206 346820 212
rect 346472 190 346808 206
rect 346922 -960 347034 480
rect 347686 439 347742 448
rect 347884 354 347912 564
rect 348068 480 348096 564
rect 349264 564 349476 592
rect 347700 326 347912 354
rect 347700 134 347728 326
rect 347688 128 347740 134
rect 347688 70 347740 76
rect 348026 -960 348138 480
rect 348772 474 349108 490
rect 349264 480 349292 564
rect 348772 468 349120 474
rect 348772 462 349068 468
rect 349068 410 349120 416
rect 349222 -960 349334 480
rect 349448 134 349476 564
rect 350184 564 350488 592
rect 350184 406 350212 564
rect 350460 480 350488 564
rect 351472 490 351500 598
rect 350172 400 350224 406
rect 350172 342 350224 348
rect 349436 128 349488 134
rect 349436 70 349488 76
rect 349876 66 350212 82
rect 349876 60 350224 66
rect 349876 54 350172 60
rect 350172 2 350224 8
rect 350418 -960 350530 480
rect 351288 462 351500 490
rect 351656 480 351684 598
rect 352840 604 352892 610
rect 352840 546 352892 552
rect 354036 604 354088 610
rect 356336 604 356388 610
rect 354036 546 354088 552
rect 355060 564 355272 592
rect 352852 480 352880 546
rect 354048 480 354076 546
rect 354680 536 354732 542
rect 354384 484 354680 490
rect 355060 490 355088 564
rect 351288 406 351316 462
rect 351276 400 351328 406
rect 351276 342 351328 348
rect 351276 264 351328 270
rect 350980 212 351276 218
rect 350980 206 351328 212
rect 350980 190 351316 206
rect 351614 -960 351726 480
rect 352472 400 352524 406
rect 352176 348 352472 354
rect 352176 342 352524 348
rect 352176 326 352512 342
rect 352810 -960 352922 480
rect 353576 128 353628 134
rect 353280 76 353576 82
rect 353280 70 353628 76
rect 353280 54 353616 70
rect 354006 -960 354118 480
rect 354384 478 354732 484
rect 354384 462 354720 478
rect 354968 462 355088 490
rect 355244 480 355272 564
rect 356684 604 357032 610
rect 356684 598 356980 604
rect 356336 546 356388 552
rect 356980 546 357032 552
rect 356348 480 356376 546
rect 357544 480 357572 614
rect 358556 598 358768 626
rect 358984 610 359320 626
rect 358984 604 359332 610
rect 358984 598 359280 604
rect 358556 542 358584 598
rect 358544 536 358596 542
rect 354968 202 354996 462
rect 354956 196 355008 202
rect 354956 138 355008 144
rect 355202 -960 355314 480
rect 355876 400 355928 406
rect 355580 348 355876 354
rect 355580 342 355928 348
rect 355580 326 355916 342
rect 356306 -960 356418 480
rect 357162 232 357218 241
rect 357162 167 357164 176
rect 357216 167 357218 176
rect 357164 138 357216 144
rect 357502 -960 357614 480
rect 358544 478 358596 484
rect 358740 480 358768 598
rect 359280 546 359332 552
rect 359752 598 359964 626
rect 361192 598 361528 626
rect 362388 610 362724 626
rect 362388 604 362736 610
rect 362388 598 362684 604
rect 358084 264 358136 270
rect 357788 212 358084 218
rect 357788 206 358136 212
rect 357788 190 358124 206
rect 358698 -960 358810 480
rect 359752 66 359780 598
rect 359936 480 359964 598
rect 360384 536 360436 542
rect 360088 484 360384 490
rect 359740 60 359792 66
rect 359740 2 359792 8
rect 359894 -960 360006 480
rect 360088 478 360436 484
rect 360088 462 360424 478
rect 361090 218 361202 480
rect 360856 202 361202 218
rect 360844 196 361202 202
rect 360896 190 361202 196
rect 360844 138 360896 144
rect 361090 -960 361202 190
rect 361500 66 361528 598
rect 363492 598 363828 626
rect 364596 598 364890 626
rect 362684 546 362736 552
rect 361946 232 362002 241
rect 361946 167 362002 176
rect 361960 82 361988 167
rect 362286 82 362398 480
rect 361488 60 361540 66
rect 361960 54 362398 82
rect 361488 2 361540 8
rect 362286 -960 362398 54
rect 363482 82 363594 480
rect 363800 474 363828 598
rect 365792 598 366128 626
rect 367008 614 367060 620
rect 368204 672 368256 678
rect 368204 614 368256 620
rect 369400 672 369452 678
rect 370412 672 370464 678
rect 369400 614 369452 620
rect 370300 620 370412 626
rect 372896 672 372948 678
rect 370300 614 370464 620
rect 364890 575 364946 584
rect 366100 513 366128 598
rect 366086 504 366142 513
rect 363788 468 363840 474
rect 363788 410 363840 416
rect 364586 354 364698 480
rect 365782 354 365894 480
rect 367020 480 367048 614
rect 368216 480 368244 614
rect 369412 480 369440 614
rect 370300 598 370452 614
rect 371496 610 371648 626
rect 381176 672 381228 678
rect 372896 614 372948 620
rect 375286 640 375342 649
rect 370688 604 370740 610
rect 370608 564 370688 592
rect 370608 480 370636 564
rect 371496 604 371660 610
rect 371496 598 371608 604
rect 370688 546 370740 552
rect 371608 546 371660 552
rect 371712 564 371924 592
rect 371712 480 371740 564
rect 366086 439 366142 448
rect 365996 400 366048 406
rect 364586 338 364840 354
rect 365782 348 365996 354
rect 365782 342 366048 348
rect 364586 332 364852 338
rect 364586 326 364800 332
rect 363696 128 363748 134
rect 363482 76 363696 82
rect 363482 70 363748 76
rect 363482 54 363736 70
rect 363482 -960 363594 54
rect 364586 -960 364698 326
rect 364800 274 364852 280
rect 365782 326 366036 342
rect 365782 -960 365894 326
rect 366744 202 366896 218
rect 366732 196 366896 202
rect 366784 190 366896 196
rect 366732 138 366784 144
rect 366978 -960 367090 480
rect 367848 202 368000 218
rect 367836 196 368000 202
rect 367888 190 368000 196
rect 367836 138 367888 144
rect 368174 -960 368286 480
rect 369044 338 369196 354
rect 369032 332 369196 338
rect 369084 326 369196 332
rect 369032 274 369084 280
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 371896 66 371924 564
rect 372436 536 372488 542
rect 372488 484 372600 490
rect 372436 478 372600 484
rect 372908 480 372936 614
rect 373920 564 374132 592
rect 375286 575 375342 584
rect 376482 640 376538 649
rect 379702 640 379758 649
rect 376482 575 376538 584
rect 372448 462 372600 478
rect 371884 60 371936 66
rect 371884 2 371936 8
rect 372866 -960 372978 480
rect 373920 270 373948 564
rect 374104 480 374132 564
rect 373908 264 373960 270
rect 373704 202 373856 218
rect 373908 206 373960 212
rect 373704 196 373868 202
rect 373704 190 373816 196
rect 373816 138 373868 144
rect 374062 -960 374174 480
rect 374900 474 375144 490
rect 375300 480 375328 575
rect 376496 480 376524 575
rect 377416 564 377720 592
rect 374900 468 375156 474
rect 374900 462 375104 468
rect 375104 410 375156 416
rect 375258 -960 375370 480
rect 376004 66 376340 82
rect 376004 60 376352 66
rect 376004 54 376300 60
rect 376300 2 376352 8
rect 376454 -960 376566 480
rect 377416 406 377444 564
rect 377692 480 377720 564
rect 378704 564 378916 592
rect 382372 672 382424 678
rect 381176 614 381228 620
rect 379702 575 379758 584
rect 377404 400 377456 406
rect 377404 342 377456 348
rect 377404 264 377456 270
rect 377108 212 377404 218
rect 377108 206 377456 212
rect 377108 190 377444 206
rect 377650 -960 377762 480
rect 378600 400 378652 406
rect 378304 348 378600 354
rect 378304 342 378652 348
rect 378304 326 378640 342
rect 378704 134 378732 564
rect 378888 480 378916 564
rect 378692 128 378744 134
rect 378692 70 378744 76
rect 378846 -960 378958 480
rect 379716 474 379744 575
rect 379808 564 380020 592
rect 379704 468 379756 474
rect 379704 410 379756 416
rect 379808 338 379836 564
rect 379992 480 380020 564
rect 381188 480 381216 614
rect 381708 610 382044 626
rect 384212 672 384264 678
rect 382372 614 382424 620
rect 383916 620 384212 626
rect 386512 672 386564 678
rect 385958 640 386014 649
rect 383916 614 384264 620
rect 381708 604 382056 610
rect 381708 598 382004 604
rect 382004 546 382056 552
rect 382384 480 382412 614
rect 383568 604 383620 610
rect 383916 598 384252 614
rect 385112 610 385448 626
rect 385112 604 385460 610
rect 385112 598 385408 604
rect 383568 546 383620 552
rect 384592 564 384804 592
rect 379796 332 379848 338
rect 379796 274 379848 280
rect 379520 128 379572 134
rect 379408 76 379520 82
rect 379408 70 379572 76
rect 379408 54 379560 70
rect 379950 -960 380062 480
rect 380512 338 380848 354
rect 380512 332 380860 338
rect 380512 326 380808 332
rect 380808 274 380860 280
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 382812 474 383148 490
rect 383580 480 383608 546
rect 382812 468 383160 474
rect 382812 462 383108 468
rect 383108 410 383160 416
rect 383538 -960 383650 480
rect 384592 202 384620 564
rect 384776 480 384804 564
rect 386216 620 386512 626
rect 400128 672 400180 678
rect 392214 640 392270 649
rect 386216 614 386564 620
rect 386216 598 386552 614
rect 389620 610 389956 626
rect 390724 610 391060 626
rect 388260 604 388312 610
rect 385958 575 386014 584
rect 385408 546 385460 552
rect 385972 480 386000 575
rect 386984 564 387196 592
rect 384580 196 384632 202
rect 384580 138 384632 144
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 386984 66 387012 564
rect 387168 480 387196 564
rect 388260 546 388312 552
rect 389456 604 389508 610
rect 389620 604 389968 610
rect 389620 598 389916 604
rect 389456 546 389508 552
rect 390724 604 391072 610
rect 390724 598 391020 604
rect 389916 546 389968 552
rect 391920 598 392214 626
rect 393024 598 393360 626
rect 392214 575 392270 584
rect 391020 546 391072 552
rect 388272 480 388300 546
rect 386972 60 387024 66
rect 386972 2 387024 8
rect 387126 -960 387238 480
rect 387320 66 387656 82
rect 387320 60 387668 66
rect 387320 54 387616 60
rect 387616 2 387668 8
rect 388230 -960 388342 480
rect 388516 474 388852 490
rect 389468 480 389496 546
rect 388516 468 388864 474
rect 388516 462 388812 468
rect 388812 410 388864 416
rect 389426 -960 389538 480
rect 390284 128 390336 134
rect 390622 82 390734 480
rect 391818 354 391930 480
rect 391584 338 391930 354
rect 391572 332 391930 338
rect 391624 326 391930 332
rect 391572 274 391624 280
rect 390336 76 390734 82
rect 390284 70 390734 76
rect 390296 54 390734 70
rect 390622 -960 390734 54
rect 391818 -960 391930 326
rect 393014 354 393126 480
rect 393228 400 393280 406
rect 393014 348 393228 354
rect 393014 342 393280 348
rect 393014 326 393268 342
rect 393014 -960 393126 326
rect 393332 134 393360 598
rect 394252 598 394464 626
rect 395324 598 395660 626
rect 398728 610 398880 626
rect 400128 614 400180 620
rect 401324 672 401376 678
rect 402428 672 402480 678
rect 401324 614 401376 620
rect 402132 620 402428 626
rect 405648 672 405700 678
rect 403622 640 403678 649
rect 402132 614 402480 620
rect 394252 480 394280 598
rect 394436 542 394464 598
rect 394424 536 394476 542
rect 393976 202 394128 218
rect 393964 196 394128 202
rect 394016 190 394128 196
rect 393964 138 394016 144
rect 393320 128 393372 134
rect 393320 70 393372 76
rect 394210 -960 394322 480
rect 394424 478 394476 484
rect 395314 354 395426 480
rect 395632 474 395660 598
rect 396540 604 396592 610
rect 396540 546 396592 552
rect 397736 604 397788 610
rect 398728 604 398892 610
rect 398728 598 398840 604
rect 397736 546 397788 552
rect 398840 546 398892 552
rect 398944 564 399156 592
rect 396264 536 396316 542
rect 396316 484 396428 490
rect 396264 478 396428 484
rect 396552 480 396580 546
rect 397748 480 397776 546
rect 398944 480 398972 564
rect 395620 468 395672 474
rect 396276 462 396428 478
rect 395620 410 395672 416
rect 395528 400 395580 406
rect 395314 348 395528 354
rect 395314 342 395580 348
rect 395314 326 395568 342
rect 395314 -960 395426 326
rect 396510 -960 396622 480
rect 397472 202 397624 218
rect 397460 196 397624 202
rect 397512 190 397624 196
rect 397460 138 397512 144
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 399128 66 399156 564
rect 400140 480 400168 614
rect 401336 480 401364 614
rect 402132 598 402468 614
rect 402532 598 402744 626
rect 402532 480 402560 598
rect 402716 542 402744 598
rect 404432 598 404584 626
rect 405536 620 405648 626
rect 407212 672 407264 678
rect 405536 614 405700 620
rect 405536 598 405688 614
rect 405844 598 406056 626
rect 407212 614 407264 620
rect 408316 672 408368 678
rect 410800 672 410852 678
rect 408368 620 408448 626
rect 408316 614 408448 620
rect 403622 575 403678 584
rect 402704 536 402756 542
rect 399832 66 399984 82
rect 399116 60 399168 66
rect 399832 60 399996 66
rect 399832 54 399944 60
rect 399116 2 399168 8
rect 399944 2 399996 8
rect 400098 -960 400210 480
rect 401140 264 401192 270
rect 401028 212 401140 218
rect 401028 206 401192 212
rect 401028 190 401180 206
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 402704 478 402756 484
rect 403236 474 403480 490
rect 403636 480 403664 575
rect 404556 542 404584 598
rect 404648 564 404860 592
rect 404544 536 404596 542
rect 403236 468 403492 474
rect 403236 462 403440 468
rect 403440 410 403492 416
rect 403594 -960 403706 480
rect 404544 478 404596 484
rect 404648 218 404676 564
rect 404832 480 404860 564
rect 405844 490 405872 598
rect 404556 190 404676 218
rect 404556 134 404584 190
rect 404544 128 404596 134
rect 404544 70 404596 76
rect 404790 -960 404902 480
rect 405752 462 405872 490
rect 406028 480 406056 598
rect 407224 480 407252 614
rect 408328 598 408448 614
rect 408420 480 408448 598
rect 409432 598 409644 626
rect 414296 672 414348 678
rect 410800 614 410852 620
rect 409236 536 409288 542
rect 408940 484 409236 490
rect 405752 134 405780 462
rect 405740 128 405792 134
rect 405740 70 405792 76
rect 405986 -960 406098 480
rect 406936 400 406988 406
rect 406640 348 406936 354
rect 406640 342 406988 348
rect 406640 326 406976 342
rect 407182 -960 407294 480
rect 408132 264 408184 270
rect 407836 212 408132 218
rect 407836 206 408184 212
rect 407836 190 408172 206
rect 408378 -960 408490 480
rect 408940 478 409288 484
rect 408940 462 409276 478
rect 409432 338 409460 598
rect 409616 480 409644 598
rect 410812 480 410840 614
rect 411640 598 411944 626
rect 409420 332 409472 338
rect 409420 274 409472 280
rect 409574 -960 409686 480
rect 410044 338 410380 354
rect 410044 332 410392 338
rect 410044 326 410340 332
rect 410340 274 410392 280
rect 410770 -960 410882 480
rect 411640 134 411668 598
rect 411916 480 411944 598
rect 412928 598 413140 626
rect 414940 672 414992 678
rect 414296 614 414348 620
rect 414644 620 414940 626
rect 415216 672 415268 678
rect 414644 614 414992 620
rect 415214 640 415216 649
rect 416044 672 416096 678
rect 415268 640 415270 649
rect 411628 128 411680 134
rect 411240 66 411576 82
rect 411628 70 411680 76
rect 411240 60 411588 66
rect 411240 54 411536 60
rect 411536 2 411588 8
rect 411874 -960 411986 480
rect 412928 202 412956 598
rect 413112 480 413140 598
rect 414308 480 414336 614
rect 414644 598 414980 614
rect 415214 575 415270 584
rect 415320 598 415532 626
rect 415748 620 416044 626
rect 424968 672 425020 678
rect 415748 614 416096 620
rect 417882 640 417938 649
rect 415748 598 416084 614
rect 416688 604 416740 610
rect 412916 196 412968 202
rect 412916 138 412968 144
rect 412640 128 412692 134
rect 412344 76 412640 82
rect 412344 70 412692 76
rect 412344 54 412680 70
rect 413070 -960 413182 480
rect 413448 202 413784 218
rect 413448 196 413796 202
rect 413448 190 413744 196
rect 413744 138 413796 144
rect 414266 -960 414378 480
rect 415320 474 415348 598
rect 415504 480 415532 598
rect 418342 640 418398 649
rect 418048 598 418342 626
rect 417882 575 417938 584
rect 420256 598 420592 626
rect 421452 598 421788 626
rect 418342 575 418398 584
rect 416688 546 416740 552
rect 416700 480 416728 546
rect 415308 468 415360 474
rect 415308 410 415360 416
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 416852 474 417188 490
rect 417896 480 417924 575
rect 418816 564 419028 592
rect 416852 468 417200 474
rect 416852 462 417148 468
rect 417148 410 417200 416
rect 417854 -960 417966 480
rect 418816 406 418844 564
rect 419000 480 419028 564
rect 418804 400 418856 406
rect 418804 342 418856 348
rect 418958 -960 419070 480
rect 419908 264 419960 270
rect 420154 218 420266 480
rect 420564 406 420592 598
rect 421012 536 421064 542
rect 421012 478 421064 484
rect 420552 400 420604 406
rect 420552 342 420604 348
rect 421024 354 421052 478
rect 421350 354 421462 480
rect 421024 326 421462 354
rect 419960 212 420266 218
rect 419908 206 420266 212
rect 419920 190 420266 206
rect 419448 128 419500 134
rect 419152 76 419448 82
rect 419152 70 419500 76
rect 419152 54 419488 70
rect 420154 -960 420266 190
rect 421350 -960 421462 326
rect 421760 270 421788 598
rect 422404 598 422556 626
rect 424968 614 425020 620
rect 426992 672 427044 678
rect 428464 672 428516 678
rect 427044 620 427156 626
rect 426992 614 427156 620
rect 423772 604 423824 610
rect 422404 542 422432 598
rect 423772 546 423824 552
rect 422392 536 422444 542
rect 422392 478 422444 484
rect 423784 480 423812 546
rect 424980 480 425008 614
rect 426164 604 426216 610
rect 427004 598 427156 614
rect 428016 610 428260 626
rect 431868 672 431920 678
rect 430854 640 430910 649
rect 428464 614 428516 620
rect 427268 604 427320 610
rect 426164 546 426216 552
rect 427268 546 427320 552
rect 428004 604 428260 610
rect 428056 598 428260 604
rect 428004 546 428056 552
rect 426176 480 426204 546
rect 427280 480 427308 546
rect 428476 480 428504 614
rect 429488 598 429700 626
rect 421748 264 421800 270
rect 421748 206 421800 212
rect 422546 218 422658 480
rect 423508 338 423660 354
rect 422760 332 422812 338
rect 422760 274 422812 280
rect 423496 332 423660 338
rect 423548 326 423660 332
rect 423496 274 423548 280
rect 422772 218 422800 274
rect 422546 190 422800 218
rect 422546 -960 422658 190
rect 423742 -960 423854 480
rect 424704 338 424856 354
rect 424692 332 424856 338
rect 424744 326 424856 332
rect 424692 274 424744 280
rect 424938 -960 425050 480
rect 425796 264 425848 270
rect 425848 212 425960 218
rect 425796 206 425960 212
rect 425808 190 425960 206
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429488 474 429516 598
rect 429672 480 429700 598
rect 431664 620 431868 626
rect 434444 672 434496 678
rect 431664 614 431920 620
rect 431664 598 431908 614
rect 432052 604 432104 610
rect 430854 575 430910 584
rect 430672 536 430724 542
rect 430560 484 430672 490
rect 429476 468 429528 474
rect 429476 410 429528 416
rect 429364 66 429516 82
rect 429364 60 429528 66
rect 429364 54 429476 60
rect 429476 2 429528 8
rect 429630 -960 429742 480
rect 430560 478 430724 484
rect 430868 480 430896 575
rect 432052 546 432104 552
rect 432984 598 433288 626
rect 434720 672 434772 678
rect 434444 614 434496 620
rect 434718 640 434720 649
rect 435364 672 435416 678
rect 434772 640 434774 649
rect 432064 480 432092 546
rect 430560 462 430712 478
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 432984 474 433012 598
rect 433260 480 433288 598
rect 434456 480 434484 614
rect 435068 620 435364 626
rect 435068 614 435416 620
rect 435548 672 435600 678
rect 437480 672 437532 678
rect 435548 614 435600 620
rect 436742 640 436798 649
rect 435068 598 435404 614
rect 434718 575 434774 584
rect 435560 480 435588 614
rect 437368 620 437480 626
rect 449624 672 449676 678
rect 437368 614 437532 620
rect 437368 598 437520 614
rect 437768 598 437980 626
rect 436742 575 436798 584
rect 436756 480 436784 575
rect 437768 490 437796 598
rect 432972 468 433024 474
rect 432972 410 433024 416
rect 432768 66 433104 82
rect 432768 60 433116 66
rect 432768 54 433064 60
rect 433064 2 433116 8
rect 433218 -960 433330 480
rect 434260 128 434312 134
rect 433964 76 434260 82
rect 433964 70 434312 76
rect 433964 54 434300 70
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436172 202 436508 218
rect 436172 196 436520 202
rect 436172 190 436468 196
rect 436468 138 436520 144
rect 436714 -960 436826 480
rect 437584 462 437796 490
rect 437952 480 437980 598
rect 438872 598 439176 626
rect 442980 610 443316 626
rect 438768 536 438820 542
rect 438472 484 438768 490
rect 437584 406 437612 462
rect 437572 400 437624 406
rect 437572 342 437624 348
rect 437910 -960 438022 480
rect 438472 478 438820 484
rect 438472 462 438808 478
rect 438872 354 438900 598
rect 439148 480 439176 598
rect 440332 604 440384 610
rect 440332 546 440384 552
rect 441528 604 441580 610
rect 441528 546 441580 552
rect 442632 604 442684 610
rect 442980 604 443328 610
rect 442980 598 443276 604
rect 442632 546 442684 552
rect 443276 546 443328 552
rect 443656 598 443868 626
rect 446384 610 446720 626
rect 440344 480 440372 546
rect 441540 480 441568 546
rect 442644 480 442672 546
rect 438780 326 438900 354
rect 438780 270 438808 326
rect 438768 264 438820 270
rect 438768 206 438820 212
rect 439106 -960 439218 480
rect 439576 66 439912 82
rect 439576 60 439924 66
rect 439576 54 439872 60
rect 439872 2 439924 8
rect 440302 -960 440414 480
rect 440772 202 441108 218
rect 440772 196 441120 202
rect 440772 190 441068 196
rect 441068 138 441120 144
rect 441498 -960 441610 480
rect 442172 400 442224 406
rect 441876 348 442172 354
rect 441876 342 442224 348
rect 441876 326 442212 342
rect 442602 -960 442714 480
rect 443656 474 443684 598
rect 443840 480 443868 598
rect 445024 604 445076 610
rect 445024 546 445076 552
rect 446220 604 446272 610
rect 446384 604 446732 610
rect 446384 598 446680 604
rect 446220 546 446272 552
rect 446680 546 446732 552
rect 447416 604 447468 610
rect 448684 598 449020 626
rect 451280 672 451332 678
rect 449676 620 449788 626
rect 449624 614 449788 620
rect 449636 598 449788 614
rect 449866 598 450032 626
rect 450984 620 451280 626
rect 454224 672 454276 678
rect 450984 614 451332 620
rect 450984 598 451320 614
rect 452088 598 452424 626
rect 453284 598 453528 626
rect 455696 672 455748 678
rect 454276 620 454388 626
rect 454224 614 454388 620
rect 456800 672 456852 678
rect 455696 614 455748 620
rect 456688 620 456800 626
rect 461952 672 462004 678
rect 459558 640 459614 649
rect 456688 614 456852 620
rect 454236 598 454388 614
rect 454500 604 454552 610
rect 447416 546 447468 552
rect 443644 468 443696 474
rect 443644 410 443696 416
rect 443798 -960 443910 480
rect 444176 474 444512 490
rect 445036 480 445064 546
rect 446232 480 446260 546
rect 447428 480 447456 546
rect 448244 536 448296 542
rect 444176 468 444524 474
rect 444176 462 444472 468
rect 444472 410 444524 416
rect 444994 -960 445106 480
rect 445280 338 445616 354
rect 445280 332 445628 338
rect 445280 326 445576 332
rect 445576 274 445628 280
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448244 478 448296 484
rect 448256 218 448284 478
rect 448582 218 448694 480
rect 448256 190 448694 218
rect 448992 202 449020 598
rect 449866 480 449894 598
rect 449778 326 449894 480
rect 450004 338 450032 598
rect 450636 536 450688 542
rect 450636 478 450688 484
rect 450648 354 450676 478
rect 450882 354 450994 480
rect 449992 332 450044 338
rect 447876 128 447928 134
rect 447580 76 447876 82
rect 447580 70 447928 76
rect 447580 54 447916 70
rect 448582 -960 448694 190
rect 448980 196 449032 202
rect 448980 138 449032 144
rect 449778 -960 449890 326
rect 450648 326 450994 354
rect 449992 274 450044 280
rect 450882 -960 450994 326
rect 452078 218 452190 480
rect 452396 338 452424 598
rect 453500 513 453528 598
rect 454500 546 454552 552
rect 453486 504 453542 513
rect 452292 332 452344 338
rect 452292 274 452344 280
rect 452384 332 452436 338
rect 452384 274 452436 280
rect 452304 218 452332 274
rect 452078 190 452332 218
rect 452078 -960 452190 190
rect 453274 82 453386 480
rect 454512 480 454540 546
rect 455708 480 455736 614
rect 456688 598 456840 614
rect 456904 598 457208 626
rect 456904 480 456932 598
rect 453486 439 453542 448
rect 453274 66 453528 82
rect 453274 60 453540 66
rect 453274 54 453488 60
rect 453274 -960 453386 54
rect 453488 2 453540 8
rect 454470 -960 454582 480
rect 455340 66 455492 82
rect 455328 60 455492 66
rect 455380 54 455492 60
rect 455328 2 455380 8
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 457180 474 457208 598
rect 458100 598 458312 626
rect 457792 474 457944 490
rect 458100 480 458128 598
rect 458284 542 458312 598
rect 459204 598 459416 626
rect 458272 536 458324 542
rect 459008 536 459060 542
rect 457168 468 457220 474
rect 457792 468 457956 474
rect 457792 462 457904 468
rect 457168 410 457220 416
rect 457904 410 457956 416
rect 458058 -960 458170 480
rect 458272 478 458324 484
rect 458896 484 459008 490
rect 458896 478 459060 484
rect 459204 480 459232 598
rect 458896 462 459048 478
rect 459162 -960 459274 480
rect 459388 270 459416 598
rect 461582 640 461638 649
rect 459558 575 459614 584
rect 460388 604 460440 610
rect 459376 264 459428 270
rect 459376 206 459428 212
rect 459572 134 459600 575
rect 461950 640 461952 649
rect 463148 672 463200 678
rect 462004 640 462006 649
rect 461582 575 461638 584
rect 461768 604 461820 610
rect 460388 546 460440 552
rect 460400 480 460428 546
rect 461596 480 461624 575
rect 463608 672 463660 678
rect 463148 614 463200 620
rect 463496 620 463608 626
rect 464896 672 464948 678
rect 463496 614 463660 620
rect 463974 640 464030 649
rect 461950 575 462006 584
rect 461768 546 461820 552
rect 462608 564 462820 592
rect 461780 513 461808 546
rect 461766 504 461822 513
rect 460204 400 460256 406
rect 460092 348 460204 354
rect 460092 342 460256 348
rect 460092 326 460244 342
rect 459560 128 459612 134
rect 459560 70 459612 76
rect 460358 -960 460470 480
rect 461196 326 461440 354
rect 461412 270 461440 326
rect 461400 264 461452 270
rect 461400 206 461452 212
rect 461554 -960 461666 480
rect 461766 439 461822 448
rect 462608 218 462636 564
rect 462792 480 462820 564
rect 463160 513 463188 614
rect 463496 598 463648 614
rect 464600 620 464896 626
rect 468392 672 468444 678
rect 464600 614 464948 620
rect 465170 640 465226 649
rect 464600 598 464936 614
rect 463974 575 464030 584
rect 469220 672 469272 678
rect 468392 614 468444 620
rect 469108 620 469220 626
rect 469108 614 469272 620
rect 471060 672 471112 678
rect 471704 672 471756 678
rect 471060 614 471112 620
rect 471408 620 471704 626
rect 474004 672 474056 678
rect 471408 614 471756 620
rect 473708 620 474004 626
rect 476764 672 476816 678
rect 476762 640 476764 649
rect 476948 672 477000 678
rect 476816 640 476818 649
rect 473708 614 474056 620
rect 467472 604 467524 610
rect 465170 575 465226 584
rect 463146 504 463202 513
rect 462516 202 462636 218
rect 462504 196 462636 202
rect 462556 190 462636 196
rect 462504 138 462556 144
rect 462412 128 462464 134
rect 462300 76 462412 82
rect 462300 70 462464 76
rect 462300 54 462452 70
rect 462750 -960 462862 480
rect 463988 480 464016 575
rect 465184 480 465212 575
rect 466104 564 466316 592
rect 466104 490 466132 564
rect 463146 439 463202 448
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 465920 462 466132 490
rect 466288 480 466316 564
rect 467472 546 467524 552
rect 467196 536 467248 542
rect 466900 484 467196 490
rect 465920 338 465948 462
rect 465908 332 465960 338
rect 465908 274 465960 280
rect 465704 202 466040 218
rect 465704 196 466052 202
rect 465704 190 466000 196
rect 466000 138 466052 144
rect 466246 -960 466358 480
rect 466900 478 467248 484
rect 467484 480 467512 546
rect 468300 536 468352 542
rect 468004 484 468300 490
rect 466900 462 467236 478
rect 467442 -960 467554 480
rect 468004 478 468352 484
rect 468404 490 468432 614
rect 469108 598 469260 614
rect 468496 564 468708 592
rect 468496 490 468524 564
rect 468004 462 468340 478
rect 468404 462 468524 490
rect 468680 480 468708 564
rect 469692 564 469904 592
rect 469496 536 469548 542
rect 468638 -960 468750 480
rect 469496 478 469548 484
rect 469508 105 469536 478
rect 469692 354 469720 564
rect 469876 480 469904 564
rect 471072 480 471100 614
rect 471408 598 471744 614
rect 473452 604 473504 610
rect 471992 564 472296 592
rect 469600 326 469720 354
rect 469494 96 469550 105
rect 469600 66 469628 326
rect 469494 31 469550 40
rect 469588 60 469640 66
rect 469588 2 469640 8
rect 469834 -960 469946 480
rect 470304 338 470640 354
rect 470304 332 470652 338
rect 470304 326 470600 332
rect 470600 274 470652 280
rect 471030 -960 471142 480
rect 471992 474 472020 564
rect 472268 480 472296 564
rect 473708 598 474044 614
rect 474812 610 475148 626
rect 474812 604 475160 610
rect 474812 598 475108 604
rect 473452 546 473504 552
rect 474384 564 474596 592
rect 471980 468 472032 474
rect 471980 410 472032 416
rect 472226 -960 472338 480
rect 472512 474 472848 490
rect 473464 480 473492 546
rect 472512 468 472860 474
rect 472512 462 472808 468
rect 472808 410 472860 416
rect 473422 -960 473534 480
rect 474384 406 474412 564
rect 474568 480 474596 564
rect 475108 546 475160 552
rect 475580 564 475792 592
rect 485136 672 485188 678
rect 481730 640 481786 649
rect 476948 614 477000 620
rect 476762 575 476818 584
rect 475580 490 475608 564
rect 474372 400 474424 406
rect 474372 342 474424 348
rect 474526 -960 474638 480
rect 475488 462 475608 490
rect 475764 480 475792 564
rect 476210 504 476266 513
rect 475488 270 475516 462
rect 475476 264 475528 270
rect 475476 206 475528 212
rect 475722 -960 475834 480
rect 475916 462 476210 490
rect 476960 480 476988 614
rect 478216 598 478552 626
rect 479320 610 479656 626
rect 479320 604 479668 610
rect 479320 598 479616 604
rect 476210 439 476266 448
rect 476918 -960 477030 480
rect 477408 128 477460 134
rect 477112 76 477408 82
rect 478114 82 478226 480
rect 477112 70 477460 76
rect 477112 54 477448 70
rect 477880 66 478226 82
rect 478524 66 478552 598
rect 480516 598 480852 626
rect 479616 546 479668 552
rect 480824 542 480852 598
rect 485134 640 485136 649
rect 486608 672 486660 678
rect 485188 640 485190 649
rect 482816 610 483152 626
rect 483768 610 483920 626
rect 482816 604 483164 610
rect 482816 598 483112 604
rect 481730 575 481786 584
rect 480812 536 480864 542
rect 479310 218 479422 480
rect 479524 400 479576 406
rect 479524 342 479576 348
rect 479536 218 479564 342
rect 479310 190 479564 218
rect 477868 60 478226 66
rect 477920 54 478226 60
rect 477868 2 477920 8
rect 478114 -960 478226 54
rect 478512 60 478564 66
rect 478512 2 478564 8
rect 479310 -960 479422 190
rect 480506 82 480618 480
rect 480812 478 480864 484
rect 481744 480 481772 575
rect 483112 546 483164 552
rect 483756 604 483920 610
rect 483808 598 483920 604
rect 484032 604 484084 610
rect 483756 546 483808 552
rect 486220 610 486372 626
rect 486436 620 486608 626
rect 487804 672 487856 678
rect 487724 632 487804 660
rect 486436 614 486660 620
rect 485134 575 485190 584
rect 485228 604 485280 610
rect 484032 546 484084 552
rect 486220 604 486384 610
rect 486220 598 486332 604
rect 485228 546 485280 552
rect 486332 546 486384 552
rect 486436 598 486648 614
rect 487324 610 487568 626
rect 487324 604 487580 610
rect 487324 598 487528 604
rect 484044 480 484072 546
rect 485240 480 485268 546
rect 486436 480 486464 598
rect 487724 592 487752 632
rect 488540 672 488592 678
rect 487804 614 487856 620
rect 488428 620 488540 626
rect 492128 672 492180 678
rect 488428 614 488592 620
rect 489918 640 489974 649
rect 488428 598 488580 614
rect 487528 546 487580 552
rect 487632 564 487752 592
rect 488828 564 489040 592
rect 489918 575 489974 584
rect 491114 640 491170 649
rect 491832 620 492128 626
rect 493324 672 493376 678
rect 491832 614 492180 620
rect 492310 640 492366 649
rect 491832 598 492168 614
rect 491114 575 491170 584
rect 492310 575 492366 584
rect 492678 640 492734 649
rect 493028 620 493324 626
rect 497832 672 497884 678
rect 495898 640 495954 649
rect 493028 614 493376 620
rect 492678 575 492734 584
rect 492864 604 492916 610
rect 487632 480 487660 564
rect 488828 480 488856 564
rect 481456 400 481508 406
rect 481508 348 481620 354
rect 481456 342 481620 348
rect 481468 326 481620 342
rect 480720 196 480772 202
rect 480720 138 480772 144
rect 480732 82 480760 138
rect 480506 54 480760 82
rect 480506 -960 480618 54
rect 481702 -960 481814 480
rect 482806 82 482918 480
rect 483018 96 483074 105
rect 482806 54 483018 82
rect 482806 -960 482918 54
rect 483018 31 483074 40
rect 484002 -960 484114 480
rect 484872 202 485024 218
rect 484860 196 485024 202
rect 484912 190 485024 196
rect 484860 138 484912 144
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489012 474 489040 564
rect 489932 480 489960 575
rect 490194 504 490250 513
rect 489000 468 489052 474
rect 489000 410 489052 416
rect 489736 400 489788 406
rect 489624 348 489736 354
rect 489624 342 489788 348
rect 489624 326 489776 342
rect 489890 -960 490002 480
rect 491128 480 491156 575
rect 491482 504 491538 513
rect 490194 439 490250 448
rect 490208 338 490236 439
rect 490728 338 490972 354
rect 490196 332 490248 338
rect 490728 332 490984 338
rect 490728 326 490932 332
rect 490196 274 490248 280
rect 490932 274 490984 280
rect 490286 96 490342 105
rect 490286 31 490288 40
rect 490340 31 490342 40
rect 490288 2 490340 8
rect 491086 -960 491198 480
rect 492324 480 492352 575
rect 491482 439 491484 448
rect 491536 439 491538 448
rect 491484 410 491536 416
rect 492282 -960 492394 480
rect 492692 270 492720 575
rect 493028 598 493364 614
rect 493508 604 493560 610
rect 492864 546 492916 552
rect 493508 546 493560 552
rect 494532 598 494744 626
rect 492680 264 492732 270
rect 492680 206 492732 212
rect 492876 105 492904 546
rect 493520 480 493548 546
rect 494532 513 494560 598
rect 494518 504 494574 513
rect 492862 96 492918 105
rect 492862 31 492918 40
rect 493478 -960 493590 480
rect 494716 480 494744 598
rect 497536 620 497832 626
rect 497536 614 497884 620
rect 498200 672 498252 678
rect 498936 672 498988 678
rect 498200 614 498252 620
rect 498640 620 498936 626
rect 504180 672 504232 678
rect 498640 614 498988 620
rect 497536 598 497872 614
rect 495898 575 495954 584
rect 494518 439 494574 448
rect 494428 264 494480 270
rect 494132 212 494428 218
rect 494132 206 494480 212
rect 494132 190 494468 206
rect 494674 -960 494786 480
rect 495236 474 495572 490
rect 495912 480 495940 575
rect 496924 564 497136 592
rect 495236 468 495584 474
rect 495236 462 495532 468
rect 495532 410 495584 416
rect 495870 -960 495982 480
rect 496924 354 496952 564
rect 497108 480 497136 564
rect 498212 480 498240 614
rect 498640 598 498976 614
rect 499396 604 499448 610
rect 499396 546 499448 552
rect 500420 598 500632 626
rect 504640 672 504692 678
rect 504180 614 504232 620
rect 504344 620 504640 626
rect 506940 672 506992 678
rect 504344 614 504692 620
rect 499408 480 499436 546
rect 500420 490 500448 598
rect 496832 326 496952 354
rect 496832 134 496860 326
rect 496820 128 496872 134
rect 496432 66 496768 82
rect 496820 70 496872 76
rect 496432 60 496780 66
rect 496432 54 496728 60
rect 496728 2 496780 8
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500328 462 500448 490
rect 500604 480 500632 598
rect 501788 604 501840 610
rect 501788 546 501840 552
rect 502984 604 503036 610
rect 502984 546 503036 552
rect 501800 480 501828 546
rect 502996 480 503024 546
rect 504192 480 504220 614
rect 504344 598 504680 614
rect 505448 598 505784 626
rect 499946 368 500002 377
rect 499946 303 500002 312
rect 499960 270 499988 303
rect 499948 264 500000 270
rect 499948 206 500000 212
rect 500328 202 500356 462
rect 500316 196 500368 202
rect 500316 138 500368 144
rect 500132 128 500184 134
rect 499836 76 500132 82
rect 499836 70 500184 76
rect 499836 54 500172 70
rect 500562 -960 500674 480
rect 500940 66 501276 82
rect 500940 60 501288 66
rect 500940 54 501236 60
rect 501236 2 501288 8
rect 501758 -960 501870 480
rect 502340 264 502392 270
rect 502044 212 502340 218
rect 502044 206 502392 212
rect 502044 190 502380 206
rect 502954 -960 503066 480
rect 503240 202 503576 218
rect 503240 196 503588 202
rect 503240 190 503536 196
rect 503536 138 503588 144
rect 504150 -960 504262 480
rect 505100 400 505152 406
rect 505346 354 505458 480
rect 505152 348 505458 354
rect 505100 342 505458 348
rect 505112 326 505458 342
rect 505346 -960 505458 326
rect 505756 66 505784 598
rect 506308 598 506520 626
rect 506644 620 506940 626
rect 507952 672 508004 678
rect 507826 632 507952 660
rect 507826 626 507854 632
rect 506644 614 506992 620
rect 506644 598 506980 614
rect 507748 598 507854 626
rect 507952 614 508004 620
rect 508596 672 508648 678
rect 509884 672 509936 678
rect 509790 640 509846 649
rect 508596 614 508648 620
rect 506308 490 506336 598
rect 506216 462 506336 490
rect 506492 480 506520 598
rect 506216 338 506244 462
rect 506204 332 506256 338
rect 506204 274 506256 280
rect 505744 60 505796 66
rect 505744 2 505796 8
rect 506450 -960 506562 480
rect 507308 332 507360 338
rect 507308 274 507360 280
rect 507320 218 507348 274
rect 507646 218 507758 480
rect 507320 190 507758 218
rect 508608 218 508636 614
rect 508944 598 509280 626
rect 508842 218 508954 480
rect 509252 338 509280 598
rect 510034 660 510062 748
rect 563408 734 563744 762
rect 565636 808 565688 814
rect 565636 750 565688 756
rect 565820 808 565872 814
rect 565820 750 565872 756
rect 509936 632 510062 660
rect 513288 672 513340 678
rect 509884 614 509936 620
rect 513564 672 513616 678
rect 513340 620 513452 626
rect 513288 614 513452 620
rect 514668 672 514720 678
rect 513564 614 513616 620
rect 514556 620 514668 626
rect 514556 614 514720 620
rect 514760 672 514812 678
rect 518256 672 518308 678
rect 517242 640 517298 649
rect 514760 614 514812 620
rect 509790 575 509846 584
rect 511264 604 511316 610
rect 509804 406 509832 575
rect 511264 546 511316 552
rect 512460 604 512512 610
rect 513300 598 513452 614
rect 512460 546 512512 552
rect 511276 480 511304 546
rect 509792 400 509844 406
rect 509792 342 509844 348
rect 510038 354 510150 480
rect 510988 400 511040 406
rect 510250 368 510306 377
rect 509240 332 509292 338
rect 509240 274 509292 280
rect 510038 326 510250 354
rect 508608 190 508954 218
rect 507646 -960 507758 190
rect 508842 -960 508954 190
rect 510038 -960 510150 326
rect 511040 348 511152 354
rect 510988 342 511152 348
rect 511000 326 511152 342
rect 510250 303 510306 312
rect 511234 -960 511346 480
rect 512196 474 512348 490
rect 512472 480 512500 546
rect 513576 480 513604 614
rect 514556 598 514708 614
rect 514772 480 514800 614
rect 516856 610 517100 626
rect 515956 604 516008 610
rect 516856 604 517112 610
rect 516856 598 517060 604
rect 515956 546 516008 552
rect 517060 546 517112 552
rect 517164 584 517242 592
rect 517960 620 518256 626
rect 519544 672 519596 678
rect 517960 614 518308 620
rect 517960 598 518296 614
rect 518360 598 518572 626
rect 519544 614 519596 620
rect 520096 672 520148 678
rect 520096 614 520148 620
rect 520740 672 520792 678
rect 522856 672 522908 678
rect 520740 614 520792 620
rect 517164 575 517298 584
rect 517164 564 517284 575
rect 515968 480 515996 546
rect 517164 480 517192 564
rect 518360 480 518388 598
rect 518544 490 518572 598
rect 519360 536 519412 542
rect 512184 468 512348 474
rect 512236 462 512348 468
rect 512184 410 512236 416
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515588 128 515640 134
rect 515640 76 515752 82
rect 515588 70 515752 76
rect 515600 54 515752 70
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 518544 462 518664 490
rect 519156 484 519360 490
rect 519156 478 519412 484
rect 519556 480 519584 614
rect 520108 542 520136 614
rect 520096 536 520148 542
rect 519156 462 519400 478
rect 518636 270 518664 462
rect 518624 264 518676 270
rect 518624 206 518676 212
rect 519514 -960 519626 480
rect 520096 478 520148 484
rect 520752 480 520780 614
rect 521672 598 521884 626
rect 522560 620 522856 626
rect 522560 614 522908 620
rect 523040 672 523092 678
rect 523960 672 524012 678
rect 523040 614 523092 620
rect 523664 620 523960 626
rect 523664 614 524012 620
rect 524236 672 524288 678
rect 525064 672 525116 678
rect 524236 614 524288 620
rect 524768 620 525064 626
rect 531872 672 531924 678
rect 529938 640 529994 649
rect 524768 614 525116 620
rect 522560 598 522896 614
rect 520372 264 520424 270
rect 520260 212 520372 218
rect 520260 206 520424 212
rect 520260 190 520412 206
rect 520710 -960 520822 480
rect 521364 202 521608 218
rect 521364 196 521620 202
rect 521364 190 521568 196
rect 521568 138 521620 144
rect 521672 66 521700 598
rect 521856 480 521884 598
rect 523052 480 523080 614
rect 523664 598 524000 614
rect 524248 480 524276 614
rect 524768 598 525104 614
rect 525168 598 525472 626
rect 521660 60 521712 66
rect 521660 2 521712 8
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525168 338 525196 598
rect 525444 480 525472 598
rect 526456 598 526668 626
rect 526456 542 526484 598
rect 526444 536 526496 542
rect 525156 332 525208 338
rect 525156 274 525208 280
rect 525402 -960 525514 480
rect 526444 478 526496 484
rect 526640 480 526668 598
rect 527652 598 527864 626
rect 527180 536 527232 542
rect 527068 484 527180 490
rect 525964 338 526300 354
rect 525964 332 526312 338
rect 525964 326 526260 332
rect 526260 274 526312 280
rect 526598 -960 526710 480
rect 527068 478 527232 484
rect 527068 462 527220 478
rect 527652 406 527680 598
rect 527836 480 527864 598
rect 528848 598 529060 626
rect 527640 400 527692 406
rect 527640 342 527692 348
rect 527794 -960 527906 480
rect 528848 474 528876 598
rect 529032 480 529060 598
rect 531576 620 531872 626
rect 535828 672 535880 678
rect 533710 640 533766 649
rect 531576 614 531924 620
rect 529938 575 529940 584
rect 529992 575 529994 584
rect 530124 604 530176 610
rect 529940 546 529992 552
rect 530124 546 530176 552
rect 531320 604 531372 610
rect 531576 598 531912 614
rect 532344 598 532556 626
rect 531320 546 531372 552
rect 530136 480 530164 546
rect 531332 480 531360 546
rect 528836 468 528888 474
rect 528836 410 528888 416
rect 528172 66 528508 82
rect 528172 60 528520 66
rect 528172 54 528468 60
rect 528468 2 528520 8
rect 528990 -960 529102 480
rect 529664 400 529716 406
rect 529368 348 529664 354
rect 529368 342 529716 348
rect 529368 326 529704 342
rect 530094 -960 530206 480
rect 530766 232 530822 241
rect 530472 190 530766 218
rect 530766 167 530822 176
rect 531290 -960 531402 480
rect 532344 134 532372 598
rect 532528 480 532556 598
rect 534170 640 534226 649
rect 533876 598 534170 626
rect 533710 575 533766 584
rect 534170 575 534226 584
rect 534540 604 534592 610
rect 533724 480 533752 575
rect 534980 598 535316 626
rect 538772 672 538824 678
rect 537574 640 537630 649
rect 535828 614 535880 620
rect 534540 546 534592 552
rect 532332 128 532384 134
rect 532332 70 532384 76
rect 532486 -960 532598 480
rect 533066 368 533122 377
rect 532772 326 533066 354
rect 533066 303 533122 312
rect 533682 -960 533794 480
rect 534552 354 534580 546
rect 534878 354 534990 480
rect 534552 326 534990 354
rect 534878 -960 534990 326
rect 535288 105 535316 598
rect 535840 218 535868 614
rect 536176 598 536512 626
rect 537280 598 537574 626
rect 536074 218 536186 480
rect 536484 406 536512 598
rect 538476 620 538772 626
rect 539140 672 539192 678
rect 538476 614 538824 620
rect 539138 640 539140 649
rect 543740 672 543792 678
rect 539192 640 539194 649
rect 541714 640 541770 649
rect 538476 598 538812 614
rect 537574 575 537630 584
rect 539580 598 539916 626
rect 539138 575 539194 584
rect 536472 400 536524 406
rect 536472 342 536524 348
rect 535840 190 536186 218
rect 536932 264 536984 270
rect 537178 218 537290 480
rect 538374 218 538486 480
rect 538862 368 538918 377
rect 538862 303 538918 312
rect 539570 354 539682 480
rect 539784 468 539836 474
rect 539784 410 539836 416
rect 539796 354 539824 410
rect 539570 326 539824 354
rect 538876 270 538904 303
rect 536984 212 537290 218
rect 536932 206 537290 212
rect 536944 190 537290 206
rect 538048 202 538486 218
rect 538864 264 538916 270
rect 538864 206 538916 212
rect 535274 96 535330 105
rect 535274 31 535330 40
rect 536074 -960 536186 190
rect 537178 -960 537290 190
rect 538036 196 538486 202
rect 538088 190 538486 196
rect 538036 138 538088 144
rect 538374 -960 538486 190
rect 539570 -960 539682 326
rect 539888 202 539916 598
rect 540796 604 540848 610
rect 541770 598 541880 626
rect 541992 604 542044 610
rect 541714 575 541770 584
rect 540796 546 540848 552
rect 541992 546 542044 552
rect 543200 598 543412 626
rect 546684 672 546736 678
rect 543740 614 543792 620
rect 540518 504 540574 513
rect 540574 462 540684 490
rect 540808 480 540836 546
rect 542004 480 542032 546
rect 543200 480 543228 598
rect 543384 490 543412 598
rect 543752 513 543780 614
rect 544212 598 544424 626
rect 544212 542 544240 598
rect 544200 536 544252 542
rect 543738 504 543794 513
rect 540518 439 540574 448
rect 539876 196 539928 202
rect 539876 138 539928 144
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 542820 264 542872 270
rect 542872 212 542984 218
rect 542820 206 542984 212
rect 542832 190 542984 206
rect 543158 -960 543270 480
rect 543384 462 543504 490
rect 543476 338 543504 462
rect 544200 478 544252 484
rect 544396 480 544424 598
rect 545500 598 545712 626
rect 548340 672 548392 678
rect 546684 614 546736 620
rect 548338 640 548340 649
rect 548984 672 549036 678
rect 548392 640 548394 649
rect 545500 480 545528 598
rect 543738 439 543794 448
rect 544088 338 544240 354
rect 543464 332 543516 338
rect 544088 332 544252 338
rect 544088 326 544200 332
rect 543464 274 543516 280
rect 544200 274 544252 280
rect 544354 -960 544466 480
rect 545132 66 545284 82
rect 545120 60 545284 66
rect 545172 54 545284 60
rect 545120 2 545172 8
rect 545458 -960 545570 480
rect 545684 134 545712 598
rect 546696 480 546724 614
rect 547892 564 548104 592
rect 548688 620 548984 626
rect 551192 672 551244 678
rect 548688 614 549036 620
rect 549074 640 549130 649
rect 548688 598 549024 614
rect 548338 575 548394 584
rect 550896 620 551192 626
rect 553308 672 553360 678
rect 550896 614 551244 620
rect 551466 640 551522 649
rect 549074 575 549130 584
rect 550272 604 550324 610
rect 547696 536 547748 542
rect 547492 484 547696 490
rect 545672 128 545724 134
rect 546500 128 546552 134
rect 545672 70 545724 76
rect 546388 76 546500 82
rect 546388 70 546552 76
rect 546388 54 546540 70
rect 546654 -960 546766 480
rect 547492 478 547748 484
rect 547892 480 547920 564
rect 547492 462 547736 478
rect 547850 -960 547962 480
rect 548076 241 548104 564
rect 549088 480 549116 575
rect 550896 598 551232 614
rect 553196 620 553308 626
rect 554596 672 554648 678
rect 553196 614 553360 620
rect 554300 620 554596 626
rect 555884 672 555936 678
rect 554300 614 554648 620
rect 554962 640 555018 649
rect 553196 598 553348 614
rect 554300 598 554636 614
rect 551466 575 551522 584
rect 550272 546 550324 552
rect 548062 232 548118 241
rect 548062 167 548118 176
rect 549046 -960 549158 480
rect 549792 474 550128 490
rect 550284 480 550312 546
rect 551480 480 551508 575
rect 552492 564 552704 592
rect 549792 468 550140 474
rect 549792 462 550088 468
rect 550088 410 550140 416
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552092 338 552428 354
rect 552092 332 552440 338
rect 552092 326 552388 332
rect 552388 274 552440 280
rect 552492 218 552520 564
rect 552676 480 552704 564
rect 553596 564 553808 592
rect 559746 640 559802 649
rect 555936 620 556200 626
rect 555884 614 556200 620
rect 555896 598 556200 614
rect 554962 575 555018 584
rect 552400 190 552520 218
rect 552400 105 552428 190
rect 552386 96 552442 105
rect 552386 31 552442 40
rect 552634 -960 552746 480
rect 553596 406 553624 564
rect 553780 480 553808 564
rect 554976 480 555004 575
rect 553584 400 553636 406
rect 553584 342 553636 348
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 555496 474 555832 490
rect 556172 480 556200 598
rect 558288 598 558592 626
rect 557184 564 557396 592
rect 555496 468 555844 474
rect 555496 462 555792 468
rect 555792 410 555844 416
rect 556130 -960 556242 480
rect 556896 400 556948 406
rect 556600 348 556896 354
rect 556600 342 556948 348
rect 556600 326 556936 342
rect 557184 202 557212 564
rect 557368 480 557396 564
rect 557172 196 557224 202
rect 557172 138 557224 144
rect 557326 -960 557438 480
rect 558288 377 558316 598
rect 558564 480 558592 598
rect 559746 575 559802 584
rect 560680 598 560892 626
rect 561108 610 561444 626
rect 561108 604 561456 610
rect 561108 598 561404 604
rect 559760 480 559788 575
rect 558274 368 558330 377
rect 557704 338 558040 354
rect 557704 332 558052 338
rect 557704 326 558000 332
rect 558274 303 558330 312
rect 558000 274 558052 280
rect 558522 -960 558634 480
rect 558900 338 559052 354
rect 558900 332 559064 338
rect 558900 326 559012 332
rect 559012 274 559064 280
rect 559718 -960 559830 480
rect 560680 270 560708 598
rect 560864 480 560892 598
rect 561404 546 561456 552
rect 562048 604 562100 610
rect 562048 546 562100 552
rect 563072 598 563284 626
rect 562060 480 562088 546
rect 560668 264 560720 270
rect 560004 202 560248 218
rect 560668 206 560720 212
rect 560004 196 560260 202
rect 560004 190 560208 196
rect 560208 138 560260 144
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 562600 264 562652 270
rect 562304 212 562600 218
rect 562304 206 562652 212
rect 562304 190 562640 206
rect 563072 66 563100 598
rect 563256 480 563284 598
rect 564452 598 564664 626
rect 564452 480 564480 598
rect 563060 60 563112 66
rect 563060 2 563112 8
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 564636 134 564664 598
rect 565648 480 565676 750
rect 565832 678 565860 750
rect 565820 672 565872 678
rect 565820 614 565872 620
rect 566844 480 566872 1158
rect 568028 808 568080 814
rect 568028 750 568080 756
rect 568040 480 568068 750
rect 569144 480 569172 3130
rect 571524 3120 571576 3126
rect 571524 3062 571576 3068
rect 569868 2848 569920 2854
rect 569868 2790 569920 2796
rect 569880 1018 569908 2790
rect 569868 1012 569920 1018
rect 569868 954 569920 960
rect 570328 740 570380 746
rect 570328 682 570380 688
rect 570340 480 570368 682
rect 571536 480 571564 3062
rect 583392 3052 583444 3058
rect 583392 2994 583444 3000
rect 572720 2916 572772 2922
rect 572720 2858 572772 2864
rect 572732 480 572760 2858
rect 576308 2848 576360 2854
rect 576308 2790 576360 2796
rect 573916 604 573968 610
rect 573916 546 573968 552
rect 575112 604 575164 610
rect 575112 546 575164 552
rect 573928 480 573956 546
rect 575124 480 575152 546
rect 576320 480 576348 2790
rect 581000 1148 581052 1154
rect 581000 1090 581052 1096
rect 577240 598 577452 626
rect 577240 490 577268 598
rect 564624 128 564676 134
rect 564624 70 564676 76
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 576872 462 577268 490
rect 577424 480 577452 598
rect 578436 598 578648 626
rect 576872 354 576900 462
rect 576780 338 576900 354
rect 576768 332 576900 338
rect 576820 326 576900 332
rect 576768 274 576820 280
rect 577382 -960 577494 480
rect 578436 354 578464 598
rect 578620 480 578648 598
rect 581012 480 581040 1090
rect 582024 598 582236 626
rect 578344 326 578464 354
rect 578344 202 578372 326
rect 578332 196 578384 202
rect 578332 138 578384 144
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582024 354 582052 598
rect 582208 480 582236 598
rect 583404 480 583432 2994
rect 581840 326 582052 354
rect 581840 270 581868 326
rect 581828 264 581880 270
rect 581828 206 581880 212
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 18 700712 74 700768
rect 662 698128 718 698184
rect 846 606056 902 606112
rect 754 553832 810 553888
rect 662 449520 718 449576
rect 570 410488 626 410544
rect 570 397432 626 397488
rect 1490 684256 1546 684312
rect 1582 632032 1638 632088
rect 1766 697720 1822 697776
rect 1674 579944 1730 580000
rect 1950 697992 2006 698048
rect 1858 527856 1914 527912
rect 1766 475632 1822 475688
rect 1950 423544 2006 423600
rect 570 214920 626 214976
rect 570 188808 626 188864
rect 202 163376 258 163432
rect 110 111152 166 111208
rect 18 71848 74 71904
rect 2134 702072 2190 702128
rect 2318 701528 2374 701584
rect 2226 254088 2282 254144
rect 2410 697584 2466 697640
rect 4342 701392 4398 701448
rect 2870 700576 2926 700632
rect 2686 697856 2742 697912
rect 3238 700440 3294 700496
rect 3054 700304 3110 700360
rect 2870 566888 2926 566944
rect 3146 658144 3202 658200
rect 3054 514800 3110 514856
rect 2686 371320 2742 371376
rect 2594 345344 2650 345400
rect 2502 319232 2558 319288
rect 3238 501744 3294 501800
rect 3330 462576 3386 462632
rect 3146 306176 3202 306232
rect 2410 267144 2466 267200
rect 2778 201864 2834 201920
rect 2318 84632 2374 84688
rect 2134 58520 2190 58576
rect 2042 32408 2098 32464
rect 3606 699896 3662 699952
rect 3514 698536 3570 698592
rect 3698 698944 3754 699000
rect 3606 149776 3662 149832
rect 3790 619112 3846 619168
rect 3698 136720 3754 136776
rect 4066 700168 4122 700224
rect 4250 671200 4306 671256
rect 31206 701800 31262 701856
rect 46018 701256 46074 701312
rect 60646 701664 60702 701720
rect 104806 700032 104862 700088
rect 217874 699760 217930 699816
rect 262862 701936 262918 701992
rect 11610 699352 11666 699408
rect 16394 699352 16450 699408
rect 65614 699352 65670 699408
rect 80150 699352 80206 699408
rect 286690 699760 286746 699816
rect 298098 699760 298154 699816
rect 336646 701800 336702 701856
rect 399022 700576 399078 700632
rect 408866 700440 408922 700496
rect 414202 700304 414258 700360
rect 458316 700168 458372 700224
rect 526718 701528 526774 701584
rect 516966 699896 517022 699952
rect 531686 701392 531742 701448
rect 546498 702072 546554 702128
rect 537022 700712 537078 700768
rect 561126 701936 561182 701992
rect 259366 699352 259422 699408
rect 418710 699352 418766 699408
rect 423678 699352 423734 699408
rect 433430 699352 433486 699408
rect 448150 699352 448206 699408
rect 468574 699352 468630 699408
rect 477590 699352 477646 699408
rect 541530 699352 541586 699408
rect 4066 358400 4122 358456
rect 3974 293120 4030 293176
rect 3882 241032 3938 241088
rect 3790 97552 3846 97608
rect 3514 45464 3570 45520
rect 3422 19352 3478 19408
rect 3054 6432 3110 6488
rect 565266 698672 565322 698728
rect 565082 698400 565138 698456
rect 569314 701664 569370 701720
rect 566462 698264 566518 698320
rect 566646 698808 566702 698864
rect 571982 700032 572038 700088
rect 577502 701256 577558 701312
rect 580262 699080 580318 699136
rect 580170 683848 580226 683904
rect 580170 670656 580226 670712
rect 580170 644000 580226 644056
rect 580170 630808 580226 630864
rect 580170 617480 580226 617536
rect 579986 590960 580042 591016
rect 579802 577632 579858 577688
rect 580170 564340 580172 564360
rect 580172 564340 580224 564360
rect 580224 564340 580226 564360
rect 580170 564304 580226 564340
rect 580170 537784 580226 537840
rect 580170 524456 580226 524512
rect 580170 511264 580226 511320
rect 580170 484608 580226 484664
rect 580170 458124 580172 458144
rect 580172 458124 580224 458144
rect 580224 458124 580226 458144
rect 580170 458088 580226 458124
rect 580170 418240 580226 418296
rect 578974 404912 579030 404968
rect 580170 378392 580226 378448
rect 580170 351872 580226 351928
rect 579986 325216 580042 325272
rect 580170 298696 580226 298752
rect 580170 258848 580226 258904
rect 580170 245556 580172 245576
rect 580172 245556 580224 245576
rect 580224 245556 580226 245576
rect 580170 245520 580226 245556
rect 579618 232328 579674 232384
rect 580170 219000 580226 219056
rect 580170 205672 580226 205728
rect 580170 192480 580226 192536
rect 580170 179152 580226 179208
rect 580170 165824 580226 165880
rect 580170 139340 580172 139360
rect 580172 139340 580224 139360
rect 580224 139340 580226 139360
rect 580170 139304 580226 139340
rect 580170 125976 580226 126032
rect 578882 112784 578938 112840
rect 579802 99456 579858 99512
rect 579618 86128 579674 86184
rect 580170 72936 580226 72992
rect 580170 46280 580226 46336
rect 580170 33108 580226 33144
rect 580170 33088 580172 33108
rect 580172 33088 580224 33108
rect 580224 33088 580226 33108
rect 580170 19760 580226 19816
rect 580906 471416 580962 471472
rect 580814 431568 580870 431624
rect 580722 365064 580778 365120
rect 580630 312024 580686 312080
rect 580538 272176 580594 272232
rect 580446 152632 580502 152688
rect 580354 59608 580410 59664
rect 580262 6568 580318 6624
rect 4066 584 4122 640
rect 7838 584 7894 640
rect 9954 584 10010 640
rect 13266 584 13322 640
rect 18510 448 18566 504
rect 20626 584 20682 640
rect 23478 584 23534 640
rect 21270 448 21326 504
rect 26514 584 26570 640
rect 28722 620 28724 640
rect 28724 620 28776 640
rect 28776 620 28778 640
rect 28722 584 28778 620
rect 27894 448 27950 504
rect 30286 584 30342 640
rect 32402 584 32458 640
rect 33230 584 33286 640
rect 35990 584 36046 640
rect 38474 584 38530 640
rect 52550 584 52606 640
rect 56046 584 56102 640
rect 54206 448 54262 504
rect 57610 584 57666 640
rect 58438 584 58494 640
rect 57426 448 57482 504
rect 59818 584 59874 640
rect 58806 448 58862 504
rect 59450 448 59506 504
rect 62026 584 62082 640
rect 61106 448 61162 504
rect 63498 584 63554 640
rect 142066 584 142122 640
rect 143446 584 143502 640
rect 144734 584 144790 640
rect 145746 584 145802 640
rect 143722 448 143778 504
rect 147126 584 147182 640
rect 148966 584 149022 640
rect 147770 448 147826 504
rect 149334 448 149390 504
rect 150622 584 150678 640
rect 151818 584 151874 640
rect 150254 448 150310 504
rect 164790 584 164846 640
rect 167366 584 167422 640
rect 169482 584 169538 640
rect 168194 312 168250 368
rect 171966 584 172022 640
rect 172978 584 173034 640
rect 170954 312 171010 368
rect 171690 312 171746 368
rect 173898 448 173954 504
rect 175462 584 175518 640
rect 176382 584 176438 640
rect 173990 312 174046 368
rect 175186 312 175242 368
rect 176842 448 176898 504
rect 177486 448 177542 504
rect 179050 584 179106 640
rect 180246 584 180302 640
rect 177670 312 177726 368
rect 178682 312 178738 368
rect 182086 584 182142 640
rect 184938 584 184994 640
rect 181258 312 181314 368
rect 188802 312 188858 368
rect 192206 312 192262 368
rect 196714 584 196770 640
rect 195242 176 195298 232
rect 197726 312 197782 368
rect 200302 584 200358 640
rect 201498 584 201554 640
rect 203614 584 203670 640
rect 198922 176 198978 232
rect 198922 40 198978 96
rect 200026 312 200082 368
rect 201314 312 201370 368
rect 202418 448 202474 504
rect 202510 40 202566 96
rect 203706 176 203762 232
rect 207386 584 207442 640
rect 208214 584 208270 640
rect 208398 584 208454 640
rect 204902 312 204958 368
rect 204810 176 204866 232
rect 206006 448 206062 504
rect 206926 448 206982 504
rect 209318 584 209374 640
rect 208766 176 208822 232
rect 210790 448 210846 504
rect 213366 584 213422 640
rect 216126 584 216182 640
rect 219990 604 220046 640
rect 219990 584 219992 604
rect 219992 584 220044 604
rect 220044 584 220046 604
rect 221830 584 221886 640
rect 223578 448 223634 504
rect 226338 584 226394 640
rect 228730 584 228786 640
rect 230938 584 230994 640
rect 235814 584 235870 640
rect 239954 584 240010 640
rect 245198 584 245254 640
rect 249062 584 249118 640
rect 249706 448 249762 504
rect 254674 584 254730 640
rect 255870 584 255926 640
rect 263138 584 263194 640
rect 264150 584 264206 640
rect 267278 584 267334 640
rect 273626 584 273682 640
rect 275190 584 275246 640
rect 281906 584 281962 640
rect 285218 448 285274 504
rect 287058 584 287114 640
rect 288990 584 289046 640
rect 292578 584 292634 640
rect 293866 584 293922 640
rect 294878 584 294934 640
rect 295614 584 295670 640
rect 303158 584 303214 640
rect 305826 584 305882 640
rect 307022 448 307078 504
rect 313830 584 313886 640
rect 315026 584 315082 640
rect 316406 584 316462 640
rect 317326 584 317382 640
rect 326342 448 326398 504
rect 336554 584 336610 640
rect 343454 604 343510 640
rect 343454 584 343456 604
rect 343456 584 343508 604
rect 343508 584 343510 604
rect 335266 448 335322 504
rect 344374 448 344430 504
rect 347686 484 347688 504
rect 347688 484 347740 504
rect 347740 484 347742 504
rect 347686 448 347742 484
rect 357162 196 357218 232
rect 357162 176 357164 196
rect 357164 176 357216 196
rect 357216 176 357218 196
rect 361946 176 362002 232
rect 364890 584 364946 640
rect 366086 448 366142 504
rect 375286 584 375342 640
rect 376482 584 376538 640
rect 379702 584 379758 640
rect 385958 584 386014 640
rect 392214 584 392270 640
rect 403622 584 403678 640
rect 415214 620 415216 640
rect 415216 620 415268 640
rect 415268 620 415270 640
rect 415214 584 415270 620
rect 417882 584 417938 640
rect 418342 584 418398 640
rect 430854 584 430910 640
rect 434718 620 434720 640
rect 434720 620 434772 640
rect 434772 620 434774 640
rect 434718 584 434774 620
rect 436742 584 436798 640
rect 453486 448 453542 504
rect 459558 584 459614 640
rect 461582 584 461638 640
rect 461950 620 461952 640
rect 461952 620 462004 640
rect 462004 620 462006 640
rect 461950 584 462006 620
rect 461766 448 461822 504
rect 463974 584 464030 640
rect 465170 584 465226 640
rect 463146 448 463202 504
rect 469494 40 469550 96
rect 476762 620 476764 640
rect 476764 620 476816 640
rect 476816 620 476818 640
rect 476762 584 476818 620
rect 476210 448 476266 504
rect 481730 584 481786 640
rect 485134 620 485136 640
rect 485136 620 485188 640
rect 485188 620 485190 640
rect 485134 584 485190 620
rect 489918 584 489974 640
rect 491114 584 491170 640
rect 492310 584 492366 640
rect 492678 584 492734 640
rect 483018 40 483074 96
rect 490194 448 490250 504
rect 490286 60 490342 96
rect 490286 40 490288 60
rect 490288 40 490340 60
rect 490340 40 490342 60
rect 491482 468 491538 504
rect 491482 448 491484 468
rect 491484 448 491536 468
rect 491536 448 491538 468
rect 492862 40 492918 96
rect 494518 448 494574 504
rect 495898 584 495954 640
rect 499946 312 500002 368
rect 509790 584 509846 640
rect 510250 312 510306 368
rect 517242 584 517298 640
rect 529938 604 529994 640
rect 529938 584 529940 604
rect 529940 584 529992 604
rect 529992 584 529994 604
rect 530766 176 530822 232
rect 533710 584 533766 640
rect 534170 584 534226 640
rect 533066 312 533122 368
rect 537574 584 537630 640
rect 539138 620 539140 640
rect 539140 620 539192 640
rect 539192 620 539194 640
rect 539138 584 539194 620
rect 538862 312 538918 368
rect 535274 40 535330 96
rect 541714 584 541770 640
rect 540518 448 540574 504
rect 543738 448 543794 504
rect 548338 620 548340 640
rect 548340 620 548392 640
rect 548392 620 548394 640
rect 548338 584 548394 620
rect 549074 584 549130 640
rect 551466 584 551522 640
rect 548062 176 548118 232
rect 554962 584 555018 640
rect 552386 40 552442 96
rect 559746 584 559802 640
rect 558274 312 558330 368
<< metal3 >>
rect 2129 702130 2195 702133
rect 546493 702130 546559 702133
rect 2129 702128 546559 702130
rect 2129 702072 2134 702128
rect 2190 702072 546498 702128
rect 546554 702072 546559 702128
rect 2129 702070 546559 702072
rect 2129 702067 2195 702070
rect 546493 702067 546559 702070
rect 262857 701994 262923 701997
rect 561121 701994 561187 701997
rect 262857 701992 561187 701994
rect 262857 701936 262862 701992
rect 262918 701936 561126 701992
rect 561182 701936 561187 701992
rect 262857 701934 561187 701936
rect 262857 701931 262923 701934
rect 561121 701931 561187 701934
rect 31201 701858 31267 701861
rect 336641 701858 336707 701861
rect 31201 701856 336707 701858
rect 31201 701800 31206 701856
rect 31262 701800 336646 701856
rect 336702 701800 336707 701856
rect 31201 701798 336707 701800
rect 31201 701795 31267 701798
rect 336641 701795 336707 701798
rect 60641 701722 60707 701725
rect 569309 701722 569375 701725
rect 60641 701720 569375 701722
rect 60641 701664 60646 701720
rect 60702 701664 569314 701720
rect 569370 701664 569375 701720
rect 60641 701662 569375 701664
rect 60641 701659 60707 701662
rect 569309 701659 569375 701662
rect 2313 701586 2379 701589
rect 526713 701586 526779 701589
rect 2313 701584 526779 701586
rect 2313 701528 2318 701584
rect 2374 701528 526718 701584
rect 526774 701528 526779 701584
rect 2313 701526 526779 701528
rect 2313 701523 2379 701526
rect 526713 701523 526779 701526
rect 4337 701450 4403 701453
rect 531681 701450 531747 701453
rect 4337 701448 531747 701450
rect 4337 701392 4342 701448
rect 4398 701392 531686 701448
rect 531742 701392 531747 701448
rect 4337 701390 531747 701392
rect 4337 701387 4403 701390
rect 531681 701387 531747 701390
rect 46013 701314 46079 701317
rect 577497 701314 577563 701317
rect 46013 701312 577563 701314
rect 46013 701256 46018 701312
rect 46074 701256 577502 701312
rect 577558 701256 577563 701312
rect 46013 701254 577563 701256
rect 46013 701251 46079 701254
rect 577497 701251 577563 701254
rect 13 700770 79 700773
rect 537017 700770 537083 700773
rect 13 700768 537083 700770
rect 13 700712 18 700768
rect 74 700712 537022 700768
rect 537078 700712 537083 700768
rect 13 700710 537083 700712
rect 13 700707 79 700710
rect 537017 700707 537083 700710
rect 2865 700634 2931 700637
rect 399017 700634 399083 700637
rect 2865 700632 399083 700634
rect 2865 700576 2870 700632
rect 2926 700576 399022 700632
rect 399078 700576 399083 700632
rect 2865 700574 399083 700576
rect 2865 700571 2931 700574
rect 399017 700571 399083 700574
rect 3233 700498 3299 700501
rect 408861 700498 408927 700501
rect 3233 700496 408927 700498
rect 3233 700440 3238 700496
rect 3294 700440 408866 700496
rect 408922 700440 408927 700496
rect 3233 700438 408927 700440
rect 3233 700435 3299 700438
rect 408861 700435 408927 700438
rect 3049 700362 3115 700365
rect 414197 700362 414263 700365
rect 3049 700360 414263 700362
rect 3049 700304 3054 700360
rect 3110 700304 414202 700360
rect 414258 700304 414263 700360
rect 3049 700302 414263 700304
rect 3049 700299 3115 700302
rect 414197 700299 414263 700302
rect 4061 700226 4127 700229
rect 458311 700226 458377 700229
rect 4061 700224 458377 700226
rect 4061 700168 4066 700224
rect 4122 700168 458316 700224
rect 458372 700168 458377 700224
rect 4061 700166 458377 700168
rect 4061 700163 4127 700166
rect 458311 700163 458377 700166
rect 104801 700090 104867 700093
rect 571977 700090 572043 700093
rect 104801 700088 572043 700090
rect 104801 700032 104806 700088
rect 104862 700032 571982 700088
rect 572038 700032 572043 700088
rect 104801 700030 572043 700032
rect 104801 700027 104867 700030
rect 571977 700027 572043 700030
rect 3601 699954 3667 699957
rect 516961 699954 517027 699957
rect 3601 699952 517027 699954
rect 3601 699896 3606 699952
rect 3662 699896 516966 699952
rect 517022 699896 517027 699952
rect 3601 699894 517027 699896
rect 3601 699891 3667 699894
rect 516961 699891 517027 699894
rect 217869 699818 217935 699821
rect 286685 699818 286751 699821
rect 298093 699818 298159 699821
rect 217869 699816 267750 699818
rect 217869 699760 217874 699816
rect 217930 699760 267750 699816
rect 217869 699758 267750 699760
rect 217869 699755 217935 699758
rect 11605 699410 11671 699413
rect 13854 699410 13860 699412
rect 11605 699408 13860 699410
rect 11605 699352 11610 699408
rect 11666 699352 13860 699408
rect 11605 699350 13860 699352
rect 11605 699347 11671 699350
rect 13854 699348 13860 699350
rect 13924 699348 13930 699412
rect 16389 699410 16455 699413
rect 21398 699410 21404 699412
rect 16389 699408 21404 699410
rect 16389 699352 16394 699408
rect 16450 699352 21404 699408
rect 16389 699350 21404 699352
rect 16389 699347 16455 699350
rect 21398 699348 21404 699350
rect 21468 699348 21474 699412
rect 65609 699410 65675 699413
rect 69974 699410 69980 699412
rect 65609 699408 69980 699410
rect 65609 699352 65614 699408
rect 65670 699352 69980 699408
rect 65609 699350 69980 699352
rect 65609 699347 65675 699350
rect 69974 699348 69980 699350
rect 70044 699348 70050 699412
rect 80145 699410 80211 699413
rect 82118 699410 82124 699412
rect 80145 699408 82124 699410
rect 80145 699352 80150 699408
rect 80206 699352 82124 699408
rect 80145 699350 82124 699352
rect 80145 699347 80211 699350
rect 82118 699348 82124 699350
rect 82188 699348 82194 699412
rect 259361 699410 259427 699413
rect 259361 699408 259562 699410
rect 259361 699352 259366 699408
rect 259422 699352 259562 699408
rect 259361 699350 259562 699352
rect 259361 699347 259427 699350
rect 259502 699138 259562 699350
rect 267690 699274 267750 699758
rect 286685 699816 298159 699818
rect 286685 699760 286690 699816
rect 286746 699760 298098 699816
rect 298154 699760 298159 699816
rect 286685 699758 298159 699760
rect 286685 699755 286751 699758
rect 298093 699755 298159 699758
rect 418705 699412 418771 699413
rect 423673 699412 423739 699413
rect 433425 699412 433491 699413
rect 448145 699412 448211 699413
rect 418654 699410 418660 699412
rect 418614 699350 418660 699410
rect 418724 699408 418771 699412
rect 423622 699410 423628 699412
rect 418766 699352 418771 699408
rect 418654 699348 418660 699350
rect 418724 699348 418771 699352
rect 423582 699350 423628 699410
rect 423692 699408 423739 699412
rect 433374 699410 433380 699412
rect 423734 699352 423739 699408
rect 423622 699348 423628 699350
rect 423692 699348 423739 699352
rect 433334 699350 433380 699410
rect 433444 699408 433491 699412
rect 448094 699410 448100 699412
rect 433486 699352 433491 699408
rect 433374 699348 433380 699350
rect 433444 699348 433491 699352
rect 448054 699350 448100 699410
rect 448164 699408 448211 699412
rect 448206 699352 448211 699408
rect 448094 699348 448100 699350
rect 448164 699348 448211 699352
rect 465758 699348 465764 699412
rect 465828 699410 465834 699412
rect 468569 699410 468635 699413
rect 477585 699412 477651 699413
rect 477534 699410 477540 699412
rect 465828 699408 468635 699410
rect 465828 699352 468574 699408
rect 468630 699352 468635 699408
rect 465828 699350 468635 699352
rect 477494 699350 477540 699410
rect 477604 699408 477651 699412
rect 477646 699352 477651 699408
rect 465828 699348 465834 699350
rect 418705 699347 418771 699348
rect 423673 699347 423739 699348
rect 433425 699347 433491 699348
rect 448145 699347 448211 699348
rect 468569 699347 468635 699350
rect 477534 699348 477540 699350
rect 477604 699348 477651 699352
rect 539910 699348 539916 699412
rect 539980 699410 539986 699412
rect 541525 699410 541591 699413
rect 539980 699408 541591 699410
rect 539980 699352 541530 699408
rect 541586 699352 541591 699408
rect 539980 699350 541591 699352
rect 539980 699348 539986 699350
rect 477585 699347 477651 699348
rect 541525 699347 541591 699350
rect 418838 699274 418844 699276
rect 267690 699214 418844 699274
rect 418838 699212 418844 699214
rect 418908 699212 418914 699276
rect 580257 699138 580323 699141
rect 259502 699136 580323 699138
rect 259502 699080 580262 699136
rect 580318 699080 580323 699136
rect 259502 699078 580323 699080
rect 580257 699075 580323 699078
rect 3693 699002 3759 699005
rect 465758 699002 465764 699004
rect 3693 699000 465764 699002
rect 3693 698944 3698 699000
rect 3754 698944 465764 699000
rect 3693 698942 465764 698944
rect 3693 698939 3759 698942
rect 465758 698940 465764 698942
rect 465828 698940 465834 699004
rect 82118 698804 82124 698868
rect 82188 698866 82194 698868
rect 566641 698866 566707 698869
rect 82188 698864 566707 698866
rect 82188 698808 566646 698864
rect 566702 698808 566707 698864
rect 82188 698806 566707 698808
rect 82188 698804 82194 698806
rect 566641 698803 566707 698806
rect 69974 698668 69980 698732
rect 70044 698730 70050 698732
rect 565261 698730 565327 698733
rect 70044 698728 565327 698730
rect 70044 698672 565266 698728
rect 565322 698672 565327 698728
rect 70044 698670 565327 698672
rect 70044 698668 70050 698670
rect 565261 698667 565327 698670
rect 3509 698594 3575 698597
rect 539910 698594 539916 698596
rect 3509 698592 539916 698594
rect 3509 698536 3514 698592
rect 3570 698536 539916 698592
rect 3509 698534 539916 698536
rect 3509 698531 3575 698534
rect 539910 698532 539916 698534
rect 539980 698532 539986 698596
rect 21398 698396 21404 698460
rect 21468 698458 21474 698460
rect 565077 698458 565143 698461
rect 21468 698456 565143 698458
rect 21468 698400 565082 698456
rect 565138 698400 565143 698456
rect 21468 698398 565143 698400
rect 21468 698396 21474 698398
rect 565077 698395 565143 698398
rect 13854 698260 13860 698324
rect 13924 698322 13930 698324
rect 566457 698322 566523 698325
rect 13924 698320 566523 698322
rect 13924 698264 566462 698320
rect 566518 698264 566523 698320
rect 13924 698262 566523 698264
rect 13924 698260 13930 698262
rect 566457 698259 566523 698262
rect 657 698186 723 698189
rect 423622 698186 423628 698188
rect 657 698184 423628 698186
rect 657 698128 662 698184
rect 718 698128 423628 698184
rect 657 698126 423628 698128
rect 657 698123 723 698126
rect 423622 698124 423628 698126
rect 423692 698124 423698 698188
rect 1945 698050 2011 698053
rect 433374 698050 433380 698052
rect 1945 698048 433380 698050
rect 1945 697992 1950 698048
rect 2006 697992 433380 698048
rect 1945 697990 433380 697992
rect 1945 697987 2011 697990
rect 433374 697988 433380 697990
rect 433444 697988 433450 698052
rect 2681 697914 2747 697917
rect 448094 697914 448100 697916
rect 2681 697912 448100 697914
rect 2681 697856 2686 697912
rect 2742 697856 448100 697912
rect 2681 697854 448100 697856
rect 2681 697851 2747 697854
rect 448094 697852 448100 697854
rect 448164 697852 448170 697916
rect 1761 697778 1827 697781
rect 418654 697778 418660 697780
rect 1761 697776 418660 697778
rect 1761 697720 1766 697776
rect 1822 697720 418660 697776
rect 1761 697718 418660 697720
rect 1761 697715 1827 697718
rect 418654 697716 418660 697718
rect 418724 697716 418730 697780
rect 418838 697716 418844 697780
rect 418908 697778 418914 697780
rect 418908 697718 583586 697778
rect 418908 697716 418914 697718
rect 2405 697642 2471 697645
rect 477534 697642 477540 697644
rect 2405 697640 477540 697642
rect 2405 697584 2410 697640
rect 2466 697584 477540 697640
rect 2405 697582 477540 697584
rect 2405 697579 2471 697582
rect 477534 697580 477540 697582
rect 477604 697580 477610 697644
rect -960 697220 480 697460
rect 583526 697370 583586 697718
rect 583342 697324 583586 697370
rect 583342 697310 584960 697324
rect 583342 697234 583402 697310
rect 583520 697234 584960 697310
rect 583342 697174 584960 697234
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 1485 684314 1551 684317
rect -960 684312 1551 684314
rect -960 684256 1490 684312
rect 1546 684256 1551 684312
rect -960 684254 1551 684256
rect -960 684164 480 684254
rect 1485 684251 1551 684254
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 4245 671258 4311 671261
rect -960 671256 4311 671258
rect -960 671200 4250 671256
rect 4306 671200 4311 671256
rect -960 671198 4311 671200
rect -960 671108 480 671198
rect 4245 671195 4311 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3141 658202 3207 658205
rect -960 658200 3207 658202
rect -960 658144 3146 658200
rect 3202 658144 3207 658200
rect -960 658142 3207 658144
rect -960 658052 480 658142
rect 3141 658139 3207 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 1577 632090 1643 632093
rect -960 632088 1643 632090
rect -960 632032 1582 632088
rect 1638 632032 1643 632088
rect -960 632030 1643 632032
rect -960 631940 480 632030
rect 1577 632027 1643 632030
rect 580165 630866 580231 630869
rect 583520 630866 584960 630956
rect 580165 630864 584960 630866
rect 580165 630808 580170 630864
rect 580226 630808 584960 630864
rect 580165 630806 584960 630808
rect 580165 630803 580231 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3785 619170 3851 619173
rect -960 619168 3851 619170
rect -960 619112 3790 619168
rect 3846 619112 3851 619168
rect -960 619110 3851 619112
rect -960 619020 480 619110
rect 3785 619107 3851 619110
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 841 606114 907 606117
rect -960 606112 907 606114
rect -960 606056 846 606112
rect 902 606056 907 606112
rect -960 606054 907 606056
rect -960 605964 480 606054
rect 841 606051 907 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 579981 591018 580047 591021
rect 583520 591018 584960 591108
rect 579981 591016 584960 591018
rect 579981 590960 579986 591016
rect 580042 590960 584960 591016
rect 579981 590958 584960 590960
rect 579981 590955 580047 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 1669 580002 1735 580005
rect -960 580000 1735 580002
rect -960 579944 1674 580000
rect 1730 579944 1735 580000
rect -960 579942 1735 579944
rect -960 579852 480 579942
rect 1669 579939 1735 579942
rect 579797 577690 579863 577693
rect 583520 577690 584960 577780
rect 579797 577688 584960 577690
rect 579797 577632 579802 577688
rect 579858 577632 584960 577688
rect 579797 577630 584960 577632
rect 579797 577627 579863 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 2865 566946 2931 566949
rect -960 566944 2931 566946
rect -960 566888 2870 566944
rect 2926 566888 2931 566944
rect -960 566886 2931 566888
rect -960 566796 480 566886
rect 2865 566883 2931 566886
rect 580165 564362 580231 564365
rect 583520 564362 584960 564452
rect 580165 564360 584960 564362
rect 580165 564304 580170 564360
rect 580226 564304 584960 564360
rect 580165 564302 584960 564304
rect 580165 564299 580231 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 749 553890 815 553893
rect -960 553888 815 553890
rect -960 553832 754 553888
rect 810 553832 815 553888
rect -960 553830 815 553832
rect -960 553740 480 553830
rect 749 553827 815 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 580165 537842 580231 537845
rect 583520 537842 584960 537932
rect 580165 537840 584960 537842
rect 580165 537784 580170 537840
rect 580226 537784 584960 537840
rect 580165 537782 584960 537784
rect 580165 537779 580231 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 1853 527914 1919 527917
rect -960 527912 1919 527914
rect -960 527856 1858 527912
rect 1914 527856 1919 527912
rect -960 527854 1919 527856
rect -960 527764 480 527854
rect 1853 527851 1919 527854
rect 580165 524514 580231 524517
rect 583520 524514 584960 524604
rect 580165 524512 584960 524514
rect 580165 524456 580170 524512
rect 580226 524456 584960 524512
rect 580165 524454 584960 524456
rect 580165 524451 580231 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 3049 514858 3115 514861
rect -960 514856 3115 514858
rect -960 514800 3054 514856
rect 3110 514800 3115 514856
rect -960 514798 3115 514800
rect -960 514708 480 514798
rect 3049 514795 3115 514798
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 3233 501802 3299 501805
rect -960 501800 3299 501802
rect -960 501744 3238 501800
rect 3294 501744 3299 501800
rect -960 501742 3299 501744
rect -960 501652 480 501742
rect 3233 501739 3299 501742
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect 1761 475690 1827 475693
rect -960 475688 1827 475690
rect -960 475632 1766 475688
rect 1822 475632 1827 475688
rect -960 475630 1827 475632
rect -960 475540 480 475630
rect 1761 475627 1827 475630
rect 580901 471474 580967 471477
rect 583520 471474 584960 471564
rect 580901 471472 584960 471474
rect 580901 471416 580906 471472
rect 580962 471416 584960 471472
rect 580901 471414 584960 471416
rect 580901 471411 580967 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 3325 462634 3391 462637
rect -960 462632 3391 462634
rect -960 462576 3330 462632
rect 3386 462576 3391 462632
rect -960 462574 3391 462576
rect -960 462484 480 462574
rect 3325 462571 3391 462574
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 580165 458083 580231 458086
rect 583520 457996 584960 458086
rect -960 449578 480 449668
rect 657 449578 723 449581
rect -960 449576 723 449578
rect -960 449520 662 449576
rect 718 449520 723 449576
rect -960 449518 723 449520
rect -960 449428 480 449518
rect 657 449515 723 449518
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 580809 431626 580875 431629
rect 583520 431626 584960 431716
rect 580809 431624 584960 431626
rect 580809 431568 580814 431624
rect 580870 431568 584960 431624
rect 580809 431566 584960 431568
rect 580809 431563 580875 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 1945 423602 2011 423605
rect -960 423600 2011 423602
rect -960 423544 1950 423600
rect 2006 423544 2011 423600
rect -960 423542 2011 423544
rect -960 423452 480 423542
rect 1945 423539 2011 423542
rect 580165 418298 580231 418301
rect 583520 418298 584960 418388
rect 580165 418296 584960 418298
rect 580165 418240 580170 418296
rect 580226 418240 584960 418296
rect 580165 418238 584960 418240
rect 580165 418235 580231 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 565 410546 631 410549
rect -960 410544 631 410546
rect -960 410488 570 410544
rect 626 410488 631 410544
rect -960 410486 631 410488
rect -960 410396 480 410486
rect 565 410483 631 410486
rect 578969 404970 579035 404973
rect 583520 404970 584960 405060
rect 578969 404968 584960 404970
rect 578969 404912 578974 404968
rect 579030 404912 584960 404968
rect 578969 404910 584960 404912
rect 578969 404907 579035 404910
rect 583520 404820 584960 404910
rect -960 397490 480 397580
rect 565 397490 631 397493
rect -960 397488 631 397490
rect -960 397432 570 397488
rect 626 397432 631 397488
rect -960 397430 631 397432
rect -960 397340 480 397430
rect 565 397427 631 397430
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 580165 378450 580231 378453
rect 583520 378450 584960 378540
rect 580165 378448 584960 378450
rect 580165 378392 580170 378448
rect 580226 378392 584960 378448
rect 580165 378390 584960 378392
rect 580165 378387 580231 378390
rect 583520 378300 584960 378390
rect -960 371378 480 371468
rect 2681 371378 2747 371381
rect -960 371376 2747 371378
rect -960 371320 2686 371376
rect 2742 371320 2747 371376
rect -960 371318 2747 371320
rect -960 371228 480 371318
rect 2681 371315 2747 371318
rect 580717 365122 580783 365125
rect 583520 365122 584960 365212
rect 580717 365120 584960 365122
rect 580717 365064 580722 365120
rect 580778 365064 584960 365120
rect 580717 365062 584960 365064
rect 580717 365059 580783 365062
rect 583520 364972 584960 365062
rect -960 358458 480 358548
rect 4061 358458 4127 358461
rect -960 358456 4127 358458
rect -960 358400 4066 358456
rect 4122 358400 4127 358456
rect -960 358398 4127 358400
rect -960 358308 480 358398
rect 4061 358395 4127 358398
rect 580165 351930 580231 351933
rect 583520 351930 584960 352020
rect 580165 351928 584960 351930
rect 580165 351872 580170 351928
rect 580226 351872 584960 351928
rect 580165 351870 584960 351872
rect 580165 351867 580231 351870
rect 583520 351780 584960 351870
rect -960 345402 480 345492
rect 2589 345402 2655 345405
rect -960 345400 2655 345402
rect -960 345344 2594 345400
rect 2650 345344 2655 345400
rect -960 345342 2655 345344
rect -960 345252 480 345342
rect 2589 345339 2655 345342
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 579981 325274 580047 325277
rect 583520 325274 584960 325364
rect 579981 325272 584960 325274
rect 579981 325216 579986 325272
rect 580042 325216 584960 325272
rect 579981 325214 584960 325216
rect 579981 325211 580047 325214
rect 583520 325124 584960 325214
rect -960 319290 480 319380
rect 2497 319290 2563 319293
rect -960 319288 2563 319290
rect -960 319232 2502 319288
rect 2558 319232 2563 319288
rect -960 319230 2563 319232
rect -960 319140 480 319230
rect 2497 319227 2563 319230
rect 580625 312082 580691 312085
rect 583520 312082 584960 312172
rect 580625 312080 584960 312082
rect 580625 312024 580630 312080
rect 580686 312024 584960 312080
rect 580625 312022 584960 312024
rect 580625 312019 580691 312022
rect 583520 311932 584960 312022
rect -960 306234 480 306324
rect 3141 306234 3207 306237
rect -960 306232 3207 306234
rect -960 306176 3146 306232
rect 3202 306176 3207 306232
rect -960 306174 3207 306176
rect -960 306084 480 306174
rect 3141 306171 3207 306174
rect 580165 298754 580231 298757
rect 583520 298754 584960 298844
rect 580165 298752 584960 298754
rect 580165 298696 580170 298752
rect 580226 298696 584960 298752
rect 580165 298694 584960 298696
rect 580165 298691 580231 298694
rect 583520 298604 584960 298694
rect -960 293178 480 293268
rect 3969 293178 4035 293181
rect -960 293176 4035 293178
rect -960 293120 3974 293176
rect 4030 293120 4035 293176
rect -960 293118 4035 293120
rect -960 293028 480 293118
rect 3969 293115 4035 293118
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 580533 272234 580599 272237
rect 583520 272234 584960 272324
rect 580533 272232 584960 272234
rect 580533 272176 580538 272232
rect 580594 272176 584960 272232
rect 580533 272174 584960 272176
rect 580533 272171 580599 272174
rect 583520 272084 584960 272174
rect -960 267202 480 267292
rect 2405 267202 2471 267205
rect -960 267200 2471 267202
rect -960 267144 2410 267200
rect 2466 267144 2471 267200
rect -960 267142 2471 267144
rect -960 267052 480 267142
rect 2405 267139 2471 267142
rect 580165 258906 580231 258909
rect 583520 258906 584960 258996
rect 580165 258904 584960 258906
rect 580165 258848 580170 258904
rect 580226 258848 584960 258904
rect 580165 258846 584960 258848
rect 580165 258843 580231 258846
rect 583520 258756 584960 258846
rect -960 254146 480 254236
rect 2221 254146 2287 254149
rect -960 254144 2287 254146
rect -960 254088 2226 254144
rect 2282 254088 2287 254144
rect -960 254086 2287 254088
rect -960 253996 480 254086
rect 2221 254083 2287 254086
rect 580165 245578 580231 245581
rect 583520 245578 584960 245668
rect 580165 245576 584960 245578
rect 580165 245520 580170 245576
rect 580226 245520 584960 245576
rect 580165 245518 584960 245520
rect 580165 245515 580231 245518
rect 583520 245428 584960 245518
rect -960 241090 480 241180
rect 3877 241090 3943 241093
rect -960 241088 3943 241090
rect -960 241032 3882 241088
rect 3938 241032 3943 241088
rect -960 241030 3943 241032
rect -960 240940 480 241030
rect 3877 241027 3943 241030
rect 579613 232386 579679 232389
rect 583520 232386 584960 232476
rect 579613 232384 584960 232386
rect 579613 232328 579618 232384
rect 579674 232328 584960 232384
rect 579613 232326 584960 232328
rect 579613 232323 579679 232326
rect 583520 232236 584960 232326
rect -960 227884 480 228124
rect 580165 219058 580231 219061
rect 583520 219058 584960 219148
rect 580165 219056 584960 219058
rect 580165 219000 580170 219056
rect 580226 219000 584960 219056
rect 580165 218998 584960 219000
rect 580165 218995 580231 218998
rect 583520 218908 584960 218998
rect -960 214978 480 215068
rect 565 214978 631 214981
rect -960 214976 631 214978
rect -960 214920 570 214976
rect 626 214920 631 214976
rect -960 214918 631 214920
rect -960 214828 480 214918
rect 565 214915 631 214918
rect 580165 205730 580231 205733
rect 583520 205730 584960 205820
rect 580165 205728 584960 205730
rect 580165 205672 580170 205728
rect 580226 205672 584960 205728
rect 580165 205670 584960 205672
rect 580165 205667 580231 205670
rect 583520 205580 584960 205670
rect -960 201922 480 202012
rect 2773 201922 2839 201925
rect -960 201920 2839 201922
rect -960 201864 2778 201920
rect 2834 201864 2839 201920
rect -960 201862 2839 201864
rect -960 201772 480 201862
rect 2773 201859 2839 201862
rect 580165 192538 580231 192541
rect 583520 192538 584960 192628
rect 580165 192536 584960 192538
rect 580165 192480 580170 192536
rect 580226 192480 584960 192536
rect 580165 192478 584960 192480
rect 580165 192475 580231 192478
rect 583520 192388 584960 192478
rect -960 188866 480 188956
rect 565 188866 631 188869
rect -960 188864 631 188866
rect -960 188808 570 188864
rect 626 188808 631 188864
rect -960 188806 631 188808
rect -960 188716 480 188806
rect 565 188803 631 188806
rect 580165 179210 580231 179213
rect 583520 179210 584960 179300
rect 580165 179208 584960 179210
rect 580165 179152 580170 179208
rect 580226 179152 584960 179208
rect 580165 179150 584960 179152
rect 580165 179147 580231 179150
rect 583520 179060 584960 179150
rect -960 175796 480 176036
rect 580165 165882 580231 165885
rect 583520 165882 584960 165972
rect 580165 165880 584960 165882
rect 580165 165824 580170 165880
rect 580226 165824 584960 165880
rect 580165 165822 584960 165824
rect 580165 165819 580231 165822
rect 583520 165732 584960 165822
rect 197 163434 263 163437
rect 197 163432 306 163434
rect 197 163376 202 163432
rect 258 163376 306 163432
rect 197 163371 306 163376
rect 246 163026 306 163371
rect 246 162980 674 163026
rect -960 162966 674 162980
rect -960 162890 480 162966
rect 614 162890 674 162966
rect -960 162830 674 162890
rect -960 162740 480 162830
rect 580441 152690 580507 152693
rect 583520 152690 584960 152780
rect 580441 152688 584960 152690
rect 580441 152632 580446 152688
rect 580502 152632 584960 152688
rect 580441 152630 584960 152632
rect 580441 152627 580507 152630
rect 583520 152540 584960 152630
rect -960 149834 480 149924
rect 3601 149834 3667 149837
rect -960 149832 3667 149834
rect -960 149776 3606 149832
rect 3662 149776 3667 149832
rect -960 149774 3667 149776
rect -960 149684 480 149774
rect 3601 149771 3667 149774
rect 580165 139362 580231 139365
rect 583520 139362 584960 139452
rect 580165 139360 584960 139362
rect 580165 139304 580170 139360
rect 580226 139304 584960 139360
rect 580165 139302 584960 139304
rect 580165 139299 580231 139302
rect 583520 139212 584960 139302
rect -960 136778 480 136868
rect 3693 136778 3759 136781
rect -960 136776 3759 136778
rect -960 136720 3698 136776
rect 3754 136720 3759 136776
rect -960 136718 3759 136720
rect -960 136628 480 136718
rect 3693 136715 3759 136718
rect 580165 126034 580231 126037
rect 583520 126034 584960 126124
rect 580165 126032 584960 126034
rect 580165 125976 580170 126032
rect 580226 125976 584960 126032
rect 580165 125974 584960 125976
rect 580165 125971 580231 125974
rect 583520 125884 584960 125974
rect -960 123572 480 123812
rect 578877 112842 578943 112845
rect 583520 112842 584960 112932
rect 578877 112840 584960 112842
rect 578877 112784 578882 112840
rect 578938 112784 584960 112840
rect 578877 112782 584960 112784
rect 578877 112779 578943 112782
rect 583520 112692 584960 112782
rect 105 111210 171 111213
rect 105 111208 306 111210
rect 105 111152 110 111208
rect 166 111152 306 111208
rect 105 111150 306 111152
rect 105 111147 171 111150
rect 246 110802 306 111150
rect 246 110756 674 110802
rect -960 110742 674 110756
rect -960 110666 480 110742
rect 614 110666 674 110742
rect -960 110606 674 110666
rect -960 110516 480 110606
rect 579797 99514 579863 99517
rect 583520 99514 584960 99604
rect 579797 99512 584960 99514
rect 579797 99456 579802 99512
rect 579858 99456 584960 99512
rect 579797 99454 584960 99456
rect 579797 99451 579863 99454
rect 583520 99364 584960 99454
rect -960 97610 480 97700
rect 3785 97610 3851 97613
rect -960 97608 3851 97610
rect -960 97552 3790 97608
rect 3846 97552 3851 97608
rect -960 97550 3851 97552
rect -960 97460 480 97550
rect 3785 97547 3851 97550
rect 579613 86186 579679 86189
rect 583520 86186 584960 86276
rect 579613 86184 584960 86186
rect 579613 86128 579618 86184
rect 579674 86128 584960 86184
rect 579613 86126 584960 86128
rect 579613 86123 579679 86126
rect 583520 86036 584960 86126
rect -960 84690 480 84780
rect 2313 84690 2379 84693
rect -960 84688 2379 84690
rect -960 84632 2318 84688
rect 2374 84632 2379 84688
rect -960 84630 2379 84632
rect -960 84540 480 84630
rect 2313 84627 2379 84630
rect 580165 72994 580231 72997
rect 583520 72994 584960 73084
rect 580165 72992 584960 72994
rect 580165 72936 580170 72992
rect 580226 72936 584960 72992
rect 580165 72934 584960 72936
rect 580165 72931 580231 72934
rect 583520 72844 584960 72934
rect 13 71906 79 71909
rect 13 71904 122 71906
rect 13 71848 18 71904
rect 74 71848 122 71904
rect 13 71843 122 71848
rect 62 71770 122 71843
rect 62 71724 674 71770
rect -960 71710 674 71724
rect -960 71634 480 71710
rect 614 71634 674 71710
rect -960 71574 674 71634
rect -960 71484 480 71574
rect 580349 59666 580415 59669
rect 583520 59666 584960 59756
rect 580349 59664 584960 59666
rect 580349 59608 580354 59664
rect 580410 59608 584960 59664
rect 580349 59606 584960 59608
rect 580349 59603 580415 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 2129 58578 2195 58581
rect -960 58576 2195 58578
rect -960 58520 2134 58576
rect 2190 58520 2195 58576
rect -960 58518 2195 58520
rect -960 58428 480 58518
rect 2129 58515 2195 58518
rect 580165 46338 580231 46341
rect 583520 46338 584960 46428
rect 580165 46336 584960 46338
rect 580165 46280 580170 46336
rect 580226 46280 584960 46336
rect 580165 46278 584960 46280
rect 580165 46275 580231 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3509 45522 3575 45525
rect -960 45520 3575 45522
rect -960 45464 3514 45520
rect 3570 45464 3575 45520
rect -960 45462 3575 45464
rect -960 45372 480 45462
rect 3509 45459 3575 45462
rect 580165 33146 580231 33149
rect 583520 33146 584960 33236
rect 580165 33144 584960 33146
rect 580165 33088 580170 33144
rect 580226 33088 584960 33144
rect 580165 33086 584960 33088
rect 580165 33083 580231 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 2037 32466 2103 32469
rect -960 32464 2103 32466
rect -960 32408 2042 32464
rect 2098 32408 2103 32464
rect -960 32406 2103 32408
rect -960 32316 480 32406
rect 2037 32403 2103 32406
rect 580165 19818 580231 19821
rect 583520 19818 584960 19908
rect 580165 19816 584960 19818
rect 580165 19760 580170 19816
rect 580226 19760 584960 19816
rect 580165 19758 584960 19760
rect 580165 19755 580231 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 580257 6626 580323 6629
rect 583520 6626 584960 6716
rect 580257 6624 584960 6626
rect -960 6490 480 6580
rect 580257 6568 580262 6624
rect 580318 6568 584960 6624
rect 580257 6566 584960 6568
rect 580257 6563 580323 6566
rect 3049 6490 3115 6493
rect -960 6488 3115 6490
rect -960 6432 3054 6488
rect 3110 6432 3115 6488
rect 583520 6476 584960 6566
rect -960 6430 3115 6432
rect -960 6340 480 6430
rect 3049 6427 3115 6430
rect 551318 914 551324 916
rect 536790 854 551324 914
rect 4061 642 4127 645
rect 7833 642 7899 645
rect 4061 640 7899 642
rect 4061 584 4066 640
rect 4122 584 7838 640
rect 7894 584 7899 640
rect 4061 582 7899 584
rect 4061 579 4127 582
rect 7833 579 7899 582
rect 9949 642 10015 645
rect 13261 642 13327 645
rect 9949 640 13327 642
rect 9949 584 9954 640
rect 10010 584 13266 640
rect 13322 584 13327 640
rect 9949 582 13327 584
rect 9949 579 10015 582
rect 13261 579 13327 582
rect 20621 642 20687 645
rect 23473 642 23539 645
rect 20621 640 23539 642
rect 20621 584 20626 640
rect 20682 584 23478 640
rect 23534 584 23539 640
rect 20621 582 23539 584
rect 20621 579 20687 582
rect 23473 579 23539 582
rect 26509 642 26575 645
rect 28717 642 28783 645
rect 30281 642 30347 645
rect 26509 640 28783 642
rect 26509 584 26514 640
rect 26570 584 28722 640
rect 28778 584 28783 640
rect 26509 582 28783 584
rect 26509 579 26575 582
rect 28717 579 28783 582
rect 29134 640 30347 642
rect 29134 584 30286 640
rect 30342 584 30347 640
rect 29134 582 30347 584
rect 18505 506 18571 509
rect 21265 506 21331 509
rect 18505 504 21331 506
rect 18505 448 18510 504
rect 18566 448 21270 504
rect 21326 448 21331 504
rect 18505 446 21331 448
rect 18505 443 18571 446
rect 21265 443 21331 446
rect 27889 506 27955 509
rect 29134 506 29194 582
rect 30281 579 30347 582
rect 32397 642 32463 645
rect 33225 642 33291 645
rect 32397 640 33291 642
rect 32397 584 32402 640
rect 32458 584 33230 640
rect 33286 584 33291 640
rect 32397 582 33291 584
rect 32397 579 32463 582
rect 33225 579 33291 582
rect 35985 642 36051 645
rect 38469 642 38535 645
rect 35985 640 38535 642
rect 35985 584 35990 640
rect 36046 584 38474 640
rect 38530 584 38535 640
rect 35985 582 38535 584
rect 35985 579 36051 582
rect 38469 579 38535 582
rect 52545 642 52611 645
rect 56041 642 56107 645
rect 57605 642 57671 645
rect 52545 640 53850 642
rect 52545 584 52550 640
rect 52606 584 53850 640
rect 52545 582 53850 584
rect 52545 579 52611 582
rect 27889 504 29194 506
rect 27889 448 27894 504
rect 27950 448 29194 504
rect 27889 446 29194 448
rect 53790 506 53850 582
rect 56041 640 57671 642
rect 56041 584 56046 640
rect 56102 584 57610 640
rect 57666 584 57671 640
rect 56041 582 57671 584
rect 56041 579 56107 582
rect 57605 579 57671 582
rect 58433 642 58499 645
rect 59813 642 59879 645
rect 58433 640 59879 642
rect 58433 584 58438 640
rect 58494 584 59818 640
rect 59874 584 59879 640
rect 58433 582 59879 584
rect 58433 579 58499 582
rect 59813 579 59879 582
rect 62021 642 62087 645
rect 63493 642 63559 645
rect 62021 640 63559 642
rect 62021 584 62026 640
rect 62082 584 63498 640
rect 63554 584 63559 640
rect 62021 582 63559 584
rect 62021 579 62087 582
rect 63493 579 63559 582
rect 142061 642 142127 645
rect 143441 642 143507 645
rect 144729 642 144795 645
rect 142061 640 142170 642
rect 142061 584 142066 640
rect 142122 584 142170 640
rect 142061 579 142170 584
rect 143441 640 144795 642
rect 143441 584 143446 640
rect 143502 584 144734 640
rect 144790 584 144795 640
rect 143441 582 144795 584
rect 143441 579 143507 582
rect 144729 579 144795 582
rect 145741 642 145807 645
rect 147121 642 147187 645
rect 145741 640 147187 642
rect 145741 584 145746 640
rect 145802 584 147126 640
rect 147182 584 147187 640
rect 145741 582 147187 584
rect 145741 579 145807 582
rect 147121 579 147187 582
rect 148961 642 149027 645
rect 150617 642 150683 645
rect 151813 642 151879 645
rect 148961 640 150683 642
rect 148961 584 148966 640
rect 149022 584 150622 640
rect 150678 584 150683 640
rect 148961 582 150683 584
rect 148961 579 149027 582
rect 150617 579 150683 582
rect 151678 640 151879 642
rect 151678 584 151818 640
rect 151874 584 151879 640
rect 151678 582 151879 584
rect 54201 506 54267 509
rect 53790 504 54267 506
rect 53790 448 54206 504
rect 54262 448 54267 504
rect 53790 446 54267 448
rect 27889 443 27955 446
rect 54201 443 54267 446
rect 57421 506 57487 509
rect 58801 506 58867 509
rect 57421 504 58867 506
rect 57421 448 57426 504
rect 57482 448 58806 504
rect 58862 448 58867 504
rect 57421 446 58867 448
rect 57421 443 57487 446
rect 58801 443 58867 446
rect 59445 506 59511 509
rect 61101 506 61167 509
rect 59445 504 61167 506
rect 59445 448 59450 504
rect 59506 448 61106 504
rect 61162 448 61167 504
rect 59445 446 61167 448
rect 142110 506 142170 579
rect 143717 506 143783 509
rect 142110 504 143783 506
rect 142110 448 143722 504
rect 143778 448 143783 504
rect 142110 446 143783 448
rect 59445 443 59511 446
rect 61101 443 61167 446
rect 143717 443 143783 446
rect 147765 506 147831 509
rect 149329 506 149395 509
rect 147765 504 149395 506
rect 147765 448 147770 504
rect 147826 448 149334 504
rect 149390 448 149395 504
rect 147765 446 149395 448
rect 147765 443 147831 446
rect 149329 443 149395 446
rect 150249 506 150315 509
rect 151678 506 151738 582
rect 151813 579 151879 582
rect 164785 642 164851 645
rect 167361 642 167427 645
rect 164785 640 167427 642
rect 164785 584 164790 640
rect 164846 584 167366 640
rect 167422 584 167427 640
rect 164785 582 167427 584
rect 164785 579 164851 582
rect 167361 579 167427 582
rect 169477 642 169543 645
rect 171961 642 172027 645
rect 169477 640 172027 642
rect 169477 584 169482 640
rect 169538 584 171966 640
rect 172022 584 172027 640
rect 169477 582 172027 584
rect 169477 579 169543 582
rect 171961 579 172027 582
rect 172973 642 173039 645
rect 175457 642 175523 645
rect 172973 640 175523 642
rect 172973 584 172978 640
rect 173034 584 175462 640
rect 175518 584 175523 640
rect 172973 582 175523 584
rect 172973 579 173039 582
rect 175457 579 175523 582
rect 176377 642 176443 645
rect 179045 642 179111 645
rect 180241 642 180307 645
rect 176377 640 179111 642
rect 176377 584 176382 640
rect 176438 584 179050 640
rect 179106 584 179111 640
rect 176377 582 179111 584
rect 176377 579 176443 582
rect 179045 579 179111 582
rect 179370 640 180307 642
rect 179370 584 180246 640
rect 180302 584 180307 640
rect 179370 582 180307 584
rect 150249 504 151738 506
rect 150249 448 150254 504
rect 150310 448 151738 504
rect 150249 446 151738 448
rect 173893 506 173959 509
rect 176837 506 176903 509
rect 173893 504 176903 506
rect 173893 448 173898 504
rect 173954 448 176842 504
rect 176898 448 176903 504
rect 173893 446 176903 448
rect 150249 443 150315 446
rect 173893 443 173959 446
rect 176837 443 176903 446
rect 177481 506 177547 509
rect 179370 506 179430 582
rect 180241 579 180307 582
rect 182081 642 182147 645
rect 184933 642 184999 645
rect 182081 640 184999 642
rect 182081 584 182086 640
rect 182142 584 184938 640
rect 184994 584 184999 640
rect 182081 582 184999 584
rect 182081 579 182147 582
rect 184933 579 184999 582
rect 196709 642 196775 645
rect 200297 642 200363 645
rect 201493 642 201559 645
rect 196709 640 200363 642
rect 196709 584 196714 640
rect 196770 584 200302 640
rect 200358 584 200363 640
rect 196709 582 200363 584
rect 196709 579 196775 582
rect 200297 579 200363 582
rect 201358 640 201559 642
rect 201358 584 201498 640
rect 201554 584 201559 640
rect 201358 582 201559 584
rect 201358 506 201418 582
rect 201493 579 201559 582
rect 203609 642 203675 645
rect 207381 642 207447 645
rect 203609 640 207447 642
rect 203609 584 203614 640
rect 203670 584 207386 640
rect 207442 584 207447 640
rect 203609 582 207447 584
rect 203609 579 203675 582
rect 207381 579 207447 582
rect 208209 642 208275 645
rect 208393 642 208459 645
rect 208209 640 208459 642
rect 208209 584 208214 640
rect 208270 584 208398 640
rect 208454 584 208459 640
rect 208209 582 208459 584
rect 208209 579 208275 582
rect 208393 579 208459 582
rect 209313 642 209379 645
rect 213361 642 213427 645
rect 209313 640 213427 642
rect 209313 584 209318 640
rect 209374 584 213366 640
rect 213422 584 213427 640
rect 209313 582 213427 584
rect 209313 579 209379 582
rect 213361 579 213427 582
rect 216121 642 216187 645
rect 219985 642 220051 645
rect 216121 640 220051 642
rect 216121 584 216126 640
rect 216182 584 219990 640
rect 220046 584 220051 640
rect 216121 582 220051 584
rect 216121 579 216187 582
rect 219985 579 220051 582
rect 221825 642 221891 645
rect 226333 642 226399 645
rect 228725 642 228791 645
rect 221825 640 226399 642
rect 221825 584 221830 640
rect 221886 584 226338 640
rect 226394 584 226399 640
rect 221825 582 226399 584
rect 221825 579 221891 582
rect 226333 579 226399 582
rect 227670 640 228791 642
rect 227670 584 228730 640
rect 228786 584 228791 640
rect 227670 582 228791 584
rect 177481 504 179430 506
rect 177481 448 177486 504
rect 177542 448 179430 504
rect 177481 446 179430 448
rect 198782 446 201418 506
rect 202413 506 202479 509
rect 206001 506 206067 509
rect 202413 504 206067 506
rect 202413 448 202418 504
rect 202474 448 206006 504
rect 206062 448 206067 504
rect 202413 446 206067 448
rect 177481 443 177547 446
rect 168189 370 168255 373
rect 170949 370 171015 373
rect 168189 368 171015 370
rect 168189 312 168194 368
rect 168250 312 170954 368
rect 171010 312 171015 368
rect 168189 310 171015 312
rect 168189 307 168255 310
rect 170949 307 171015 310
rect 171685 370 171751 373
rect 173985 370 174051 373
rect 171685 368 174051 370
rect 171685 312 171690 368
rect 171746 312 173990 368
rect 174046 312 174051 368
rect 171685 310 174051 312
rect 171685 307 171751 310
rect 173985 307 174051 310
rect 175181 370 175247 373
rect 177665 370 177731 373
rect 175181 368 177731 370
rect 175181 312 175186 368
rect 175242 312 177670 368
rect 177726 312 177731 368
rect 175181 310 177731 312
rect 175181 307 175247 310
rect 177665 307 177731 310
rect 178677 370 178743 373
rect 181253 370 181319 373
rect 178677 368 181319 370
rect 178677 312 178682 368
rect 178738 312 181258 368
rect 181314 312 181319 368
rect 178677 310 181319 312
rect 178677 307 178743 310
rect 181253 307 181319 310
rect 188797 370 188863 373
rect 192201 370 192267 373
rect 188797 368 192267 370
rect 188797 312 188802 368
rect 188858 312 192206 368
rect 192262 312 192267 368
rect 188797 310 192267 312
rect 188797 307 188863 310
rect 192201 307 192267 310
rect 197721 370 197787 373
rect 198782 370 198842 446
rect 202413 443 202479 446
rect 206001 443 206067 446
rect 206921 506 206987 509
rect 210785 506 210851 509
rect 206921 504 210851 506
rect 206921 448 206926 504
rect 206982 448 210790 504
rect 210846 448 210851 504
rect 206921 446 210851 448
rect 206921 443 206987 446
rect 210785 443 210851 446
rect 223573 506 223639 509
rect 227670 506 227730 582
rect 228725 579 228791 582
rect 230933 642 230999 645
rect 235809 642 235875 645
rect 230933 640 235875 642
rect 230933 584 230938 640
rect 230994 584 235814 640
rect 235870 584 235875 640
rect 230933 582 235875 584
rect 230933 579 230999 582
rect 235809 579 235875 582
rect 239949 642 240015 645
rect 245193 642 245259 645
rect 239949 640 245259 642
rect 239949 584 239954 640
rect 240010 584 245198 640
rect 245254 584 245259 640
rect 239949 582 245259 584
rect 239949 579 240015 582
rect 245193 579 245259 582
rect 249057 642 249123 645
rect 254669 642 254735 645
rect 255865 642 255931 645
rect 249057 640 254735 642
rect 249057 584 249062 640
rect 249118 584 254674 640
rect 254730 584 254735 640
rect 249057 582 254735 584
rect 249057 579 249123 582
rect 254669 579 254735 582
rect 255822 640 255931 642
rect 255822 584 255870 640
rect 255926 584 255931 640
rect 255822 579 255931 584
rect 263133 642 263199 645
rect 264145 642 264211 645
rect 263133 640 264211 642
rect 263133 584 263138 640
rect 263194 584 264150 640
rect 264206 584 264211 640
rect 263133 582 264211 584
rect 263133 579 263199 582
rect 264145 579 264211 582
rect 267273 642 267339 645
rect 273621 642 273687 645
rect 267273 640 273687 642
rect 267273 584 267278 640
rect 267334 584 273626 640
rect 273682 584 273687 640
rect 267273 582 273687 584
rect 267273 579 267339 582
rect 273621 579 273687 582
rect 275185 642 275251 645
rect 281901 642 281967 645
rect 275185 640 281967 642
rect 275185 584 275190 640
rect 275246 584 281906 640
rect 281962 584 281967 640
rect 275185 582 281967 584
rect 275185 579 275251 582
rect 281901 579 281967 582
rect 287053 642 287119 645
rect 288985 642 289051 645
rect 292573 642 292639 645
rect 287053 640 289051 642
rect 287053 584 287058 640
rect 287114 584 288990 640
rect 289046 584 289051 640
rect 287053 582 289051 584
rect 287053 579 287119 582
rect 288985 579 289051 582
rect 289126 640 292639 642
rect 289126 584 292578 640
rect 292634 584 292639 640
rect 289126 582 292639 584
rect 223573 504 227730 506
rect 223573 448 223578 504
rect 223634 448 227730 504
rect 223573 446 227730 448
rect 249701 506 249767 509
rect 255822 506 255882 579
rect 249701 504 255882 506
rect 249701 448 249706 504
rect 249762 448 255882 504
rect 249701 446 255882 448
rect 285213 506 285279 509
rect 289126 506 289186 582
rect 292573 579 292639 582
rect 293861 642 293927 645
rect 294873 642 294939 645
rect 293861 640 294939 642
rect 293861 584 293866 640
rect 293922 584 294878 640
rect 294934 584 294939 640
rect 293861 582 294939 584
rect 293861 579 293927 582
rect 294873 579 294939 582
rect 295609 642 295675 645
rect 303153 642 303219 645
rect 295609 640 303219 642
rect 295609 584 295614 640
rect 295670 584 303158 640
rect 303214 584 303219 640
rect 295609 582 303219 584
rect 295609 579 295675 582
rect 303153 579 303219 582
rect 305821 642 305887 645
rect 313825 642 313891 645
rect 315021 642 315087 645
rect 305821 640 313891 642
rect 305821 584 305826 640
rect 305882 584 313830 640
rect 313886 584 313891 640
rect 305821 582 313891 584
rect 305821 579 305887 582
rect 313825 579 313891 582
rect 314886 640 315087 642
rect 314886 584 315026 640
rect 315082 584 315087 640
rect 314886 582 315087 584
rect 285213 504 289186 506
rect 285213 448 285218 504
rect 285274 448 289186 504
rect 285213 446 289186 448
rect 307017 506 307083 509
rect 314886 506 314946 582
rect 315021 579 315087 582
rect 316401 642 316467 645
rect 317321 642 317387 645
rect 316401 640 317387 642
rect 316401 584 316406 640
rect 316462 584 317326 640
rect 317382 584 317387 640
rect 316401 582 317387 584
rect 316401 579 316467 582
rect 317321 579 317387 582
rect 336549 642 336615 645
rect 343449 642 343515 645
rect 336549 640 343515 642
rect 336549 584 336554 640
rect 336610 584 343454 640
rect 343510 584 343515 640
rect 336549 582 343515 584
rect 336549 579 336615 582
rect 343449 579 343515 582
rect 364885 642 364951 645
rect 375281 642 375347 645
rect 376477 642 376543 645
rect 364885 640 375347 642
rect 364885 584 364890 640
rect 364946 584 375286 640
rect 375342 584 375347 640
rect 364885 582 375347 584
rect 364885 579 364951 582
rect 375281 579 375347 582
rect 375422 640 376543 642
rect 375422 584 376482 640
rect 376538 584 376543 640
rect 375422 582 376543 584
rect 307017 504 314946 506
rect 307017 448 307022 504
rect 307078 448 314946 504
rect 307017 446 314946 448
rect 326337 506 326403 509
rect 335261 506 335327 509
rect 326337 504 335327 506
rect 326337 448 326342 504
rect 326398 448 335266 504
rect 335322 448 335327 504
rect 326337 446 335327 448
rect 223573 443 223639 446
rect 249701 443 249767 446
rect 285213 443 285279 446
rect 307017 443 307083 446
rect 326337 443 326403 446
rect 335261 443 335327 446
rect 344369 506 344435 509
rect 347681 506 347747 509
rect 344369 504 347747 506
rect 344369 448 344374 504
rect 344430 448 347686 504
rect 347742 448 347747 504
rect 344369 446 347747 448
rect 344369 443 344435 446
rect 347681 443 347747 446
rect 366081 506 366147 509
rect 375422 506 375482 582
rect 376477 579 376543 582
rect 379697 642 379763 645
rect 385953 642 386019 645
rect 379697 640 386019 642
rect 379697 584 379702 640
rect 379758 584 385958 640
rect 386014 584 386019 640
rect 379697 582 386019 584
rect 379697 579 379763 582
rect 385953 579 386019 582
rect 392209 642 392275 645
rect 403617 642 403683 645
rect 392209 640 403683 642
rect 392209 584 392214 640
rect 392270 584 403622 640
rect 403678 584 403683 640
rect 392209 582 403683 584
rect 392209 579 392275 582
rect 403617 579 403683 582
rect 415209 642 415275 645
rect 417877 642 417943 645
rect 415209 640 417943 642
rect 415209 584 415214 640
rect 415270 584 417882 640
rect 417938 584 417943 640
rect 415209 582 417943 584
rect 415209 579 415275 582
rect 417877 579 417943 582
rect 418337 642 418403 645
rect 430849 642 430915 645
rect 418337 640 430915 642
rect 418337 584 418342 640
rect 418398 584 430854 640
rect 430910 584 430915 640
rect 418337 582 430915 584
rect 418337 579 418403 582
rect 430849 579 430915 582
rect 434713 642 434779 645
rect 436737 642 436803 645
rect 434713 640 436803 642
rect 434713 584 434718 640
rect 434774 584 436742 640
rect 436798 584 436803 640
rect 434713 582 436803 584
rect 434713 579 434779 582
rect 436737 579 436803 582
rect 459553 642 459619 645
rect 461577 642 461643 645
rect 459553 640 461643 642
rect 459553 584 459558 640
rect 459614 584 461582 640
rect 461638 584 461643 640
rect 459553 582 461643 584
rect 459553 579 459619 582
rect 461577 579 461643 582
rect 461945 642 462011 645
rect 463969 642 464035 645
rect 465165 642 465231 645
rect 461945 640 464035 642
rect 461945 584 461950 640
rect 462006 584 463974 640
rect 464030 584 464035 640
rect 461945 582 464035 584
rect 461945 579 462011 582
rect 463969 579 464035 582
rect 465030 640 465231 642
rect 465030 584 465170 640
rect 465226 584 465231 640
rect 465030 582 465231 584
rect 366081 504 375482 506
rect 366081 448 366086 504
rect 366142 448 375482 504
rect 366081 446 375482 448
rect 453481 506 453547 509
rect 461761 506 461827 509
rect 453481 504 461827 506
rect 453481 448 453486 504
rect 453542 448 461766 504
rect 461822 448 461827 504
rect 453481 446 461827 448
rect 366081 443 366147 446
rect 453481 443 453547 446
rect 461761 443 461827 446
rect 463141 506 463207 509
rect 465030 506 465090 582
rect 465165 579 465231 582
rect 476757 642 476823 645
rect 481725 642 481791 645
rect 476757 640 481791 642
rect 476757 584 476762 640
rect 476818 584 481730 640
rect 481786 584 481791 640
rect 476757 582 481791 584
rect 476757 579 476823 582
rect 481725 579 481791 582
rect 485129 642 485195 645
rect 489913 642 489979 645
rect 491109 642 491175 645
rect 492305 642 492371 645
rect 485129 640 489979 642
rect 485129 584 485134 640
rect 485190 584 489918 640
rect 489974 584 489979 640
rect 485129 582 489979 584
rect 485129 579 485195 582
rect 489913 579 489979 582
rect 490054 640 491175 642
rect 490054 584 491114 640
rect 491170 584 491175 640
rect 490054 582 491175 584
rect 463141 504 465090 506
rect 463141 448 463146 504
rect 463202 448 465090 504
rect 463141 446 465090 448
rect 476205 506 476271 509
rect 490054 506 490114 582
rect 491109 579 491175 582
rect 491342 640 492371 642
rect 491342 584 492310 640
rect 492366 584 492371 640
rect 491342 582 492371 584
rect 476205 504 490114 506
rect 476205 448 476210 504
rect 476266 448 490114 504
rect 476205 446 490114 448
rect 490189 506 490255 509
rect 491342 506 491402 582
rect 492305 579 492371 582
rect 492673 642 492739 645
rect 495893 642 495959 645
rect 492673 640 495959 642
rect 492673 584 492678 640
rect 492734 584 495898 640
rect 495954 584 495959 640
rect 492673 582 495959 584
rect 492673 579 492739 582
rect 495893 579 495959 582
rect 509785 642 509851 645
rect 517237 642 517303 645
rect 509785 640 517303 642
rect 509785 584 509790 640
rect 509846 584 517242 640
rect 517298 584 517303 640
rect 509785 582 517303 584
rect 509785 579 509851 582
rect 517237 579 517303 582
rect 529933 642 529999 645
rect 533705 642 533771 645
rect 529933 640 533771 642
rect 529933 584 529938 640
rect 529994 584 533710 640
rect 533766 584 533771 640
rect 529933 582 533771 584
rect 529933 579 529999 582
rect 533705 579 533771 582
rect 534165 642 534231 645
rect 536790 642 536850 854
rect 551318 852 551324 854
rect 551388 852 551394 916
rect 546450 718 557550 778
rect 534165 640 536850 642
rect 534165 584 534170 640
rect 534226 584 536850 640
rect 534165 582 536850 584
rect 537569 642 537635 645
rect 539133 642 539199 645
rect 537569 640 539199 642
rect 537569 584 537574 640
rect 537630 584 539138 640
rect 539194 584 539199 640
rect 537569 582 539199 584
rect 534165 579 534231 582
rect 537569 579 537635 582
rect 539133 579 539199 582
rect 541709 642 541775 645
rect 546450 642 546510 718
rect 541709 640 546510 642
rect 541709 584 541714 640
rect 541770 584 546510 640
rect 541709 582 546510 584
rect 548333 642 548399 645
rect 549069 642 549135 645
rect 548333 640 549135 642
rect 548333 584 548338 640
rect 548394 584 549074 640
rect 549130 584 549135 640
rect 548333 582 549135 584
rect 541709 579 541775 582
rect 548333 579 548399 582
rect 549069 579 549135 582
rect 551318 580 551324 644
rect 551388 642 551394 644
rect 551461 642 551527 645
rect 554957 642 555023 645
rect 551388 640 551527 642
rect 551388 584 551466 640
rect 551522 584 551527 640
rect 551388 582 551527 584
rect 551388 580 551394 582
rect 551461 579 551527 582
rect 554822 640 555023 642
rect 554822 584 554962 640
rect 555018 584 555023 640
rect 554822 582 555023 584
rect 557490 642 557550 718
rect 559741 642 559807 645
rect 557490 640 559807 642
rect 557490 584 559746 640
rect 559802 584 559807 640
rect 557490 582 559807 584
rect 490189 504 491402 506
rect 490189 448 490194 504
rect 490250 448 491402 504
rect 490189 446 491402 448
rect 491477 506 491543 509
rect 494513 506 494579 509
rect 491477 504 494579 506
rect 491477 448 491482 504
rect 491538 448 494518 504
rect 494574 448 494579 504
rect 491477 446 494579 448
rect 463141 443 463207 446
rect 476205 443 476271 446
rect 490189 443 490255 446
rect 491477 443 491543 446
rect 494513 443 494579 446
rect 540513 506 540579 509
rect 543733 506 543799 509
rect 554822 506 554882 582
rect 554957 579 555023 582
rect 559741 579 559807 582
rect 540513 504 543658 506
rect 540513 448 540518 504
rect 540574 448 543658 504
rect 540513 446 543658 448
rect 540513 443 540579 446
rect 197721 368 198842 370
rect 197721 312 197726 368
rect 197782 312 198842 368
rect 197721 310 198842 312
rect 200021 370 200087 373
rect 201309 370 201375 373
rect 204897 370 204963 373
rect 200021 368 200130 370
rect 200021 312 200026 368
rect 200082 312 200130 368
rect 197721 307 197787 310
rect 200021 307 200130 312
rect 201309 368 204963 370
rect 201309 312 201314 368
rect 201370 312 204902 368
rect 204958 312 204963 368
rect 201309 310 204963 312
rect 201309 307 201375 310
rect 204897 307 204963 310
rect 499941 370 500007 373
rect 510245 370 510311 373
rect 499941 368 510311 370
rect 499941 312 499946 368
rect 500002 312 510250 368
rect 510306 312 510311 368
rect 499941 310 510311 312
rect 499941 307 500007 310
rect 510245 307 510311 310
rect 533061 370 533127 373
rect 538857 370 538923 373
rect 533061 368 538923 370
rect 533061 312 533066 368
rect 533122 312 538862 368
rect 538918 312 538923 368
rect 533061 310 538923 312
rect 543598 370 543658 446
rect 543733 504 554882 506
rect 543733 448 543738 504
rect 543794 448 554882 504
rect 543733 446 554882 448
rect 543733 443 543799 446
rect 558269 370 558335 373
rect 543598 368 558335 370
rect 543598 312 558274 368
rect 558330 312 558335 368
rect 543598 310 558335 312
rect 533061 307 533127 310
rect 538857 307 538923 310
rect 558269 307 558335 310
rect 195237 234 195303 237
rect 198917 234 198983 237
rect 195237 232 198983 234
rect 195237 176 195242 232
rect 195298 176 198922 232
rect 198978 176 198983 232
rect 195237 174 198983 176
rect 200070 234 200130 307
rect 203701 234 203767 237
rect 200070 232 203767 234
rect 200070 176 203706 232
rect 203762 176 203767 232
rect 200070 174 203767 176
rect 195237 171 195303 174
rect 198917 171 198983 174
rect 203701 171 203767 174
rect 204805 234 204871 237
rect 208761 234 208827 237
rect 204805 232 208827 234
rect 204805 176 204810 232
rect 204866 176 208766 232
rect 208822 176 208827 232
rect 204805 174 208827 176
rect 204805 171 204871 174
rect 208761 171 208827 174
rect 357157 234 357223 237
rect 361941 234 362007 237
rect 357157 232 362007 234
rect 357157 176 357162 232
rect 357218 176 361946 232
rect 362002 176 362007 232
rect 357157 174 362007 176
rect 357157 171 357223 174
rect 361941 171 362007 174
rect 530761 234 530827 237
rect 548057 234 548123 237
rect 530761 232 548123 234
rect 530761 176 530766 232
rect 530822 176 548062 232
rect 548118 176 548123 232
rect 530761 174 548123 176
rect 530761 171 530827 174
rect 548057 171 548123 174
rect 198917 98 198983 101
rect 202505 98 202571 101
rect 198917 96 202571 98
rect 198917 40 198922 96
rect 198978 40 202510 96
rect 202566 40 202571 96
rect 198917 38 202571 40
rect 198917 35 198983 38
rect 202505 35 202571 38
rect 469489 98 469555 101
rect 483013 98 483079 101
rect 469489 96 483079 98
rect 469489 40 469494 96
rect 469550 40 483018 96
rect 483074 40 483079 96
rect 469489 38 483079 40
rect 469489 35 469555 38
rect 483013 35 483079 38
rect 490281 98 490347 101
rect 492857 98 492923 101
rect 490281 96 492923 98
rect 490281 40 490286 96
rect 490342 40 492862 96
rect 492918 40 492923 96
rect 490281 38 492923 40
rect 490281 35 490347 38
rect 492857 35 492923 38
rect 535269 98 535335 101
rect 552381 98 552447 101
rect 535269 96 552447 98
rect 535269 40 535274 96
rect 535330 40 552386 96
rect 552442 40 552447 96
rect 535269 38 552447 40
rect 535269 35 535335 38
rect 552381 35 552447 38
<< via3 >>
rect 13860 699348 13924 699412
rect 21404 699348 21468 699412
rect 69980 699348 70044 699412
rect 82124 699348 82188 699412
rect 418660 699408 418724 699412
rect 418660 699352 418710 699408
rect 418710 699352 418724 699408
rect 418660 699348 418724 699352
rect 423628 699408 423692 699412
rect 423628 699352 423678 699408
rect 423678 699352 423692 699408
rect 423628 699348 423692 699352
rect 433380 699408 433444 699412
rect 433380 699352 433430 699408
rect 433430 699352 433444 699408
rect 433380 699348 433444 699352
rect 448100 699408 448164 699412
rect 448100 699352 448150 699408
rect 448150 699352 448164 699408
rect 448100 699348 448164 699352
rect 465764 699348 465828 699412
rect 477540 699408 477604 699412
rect 477540 699352 477590 699408
rect 477590 699352 477604 699408
rect 477540 699348 477604 699352
rect 539916 699348 539980 699412
rect 418844 699212 418908 699276
rect 465764 698940 465828 699004
rect 82124 698804 82188 698868
rect 69980 698668 70044 698732
rect 539916 698532 539980 698596
rect 21404 698396 21468 698460
rect 13860 698260 13924 698324
rect 423628 698124 423692 698188
rect 433380 697988 433444 698052
rect 448100 697852 448164 697916
rect 418660 697716 418724 697780
rect 418844 697716 418908 697780
rect 477540 697580 477604 697644
rect 551324 852 551388 916
rect 551324 580 551388 644
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 680614 -8106 711002
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 -8106 680614
rect -8726 680294 -8106 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 -8106 680294
rect -8726 644614 -8106 680058
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 -8106 644614
rect -8726 644294 -8106 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 -8106 644294
rect -8726 608614 -8106 644058
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 -8106 608614
rect -8726 608294 -8106 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 -8106 608294
rect -8726 572614 -8106 608058
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 -8106 572614
rect -8726 572294 -8106 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 -8106 572294
rect -8726 536614 -8106 572058
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 -8106 536614
rect -8726 536294 -8106 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 -8106 536294
rect -8726 500614 -8106 536058
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 -8106 500614
rect -8726 500294 -8106 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 -8106 500294
rect -8726 464614 -8106 500058
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 -8106 464614
rect -8726 464294 -8106 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 -8106 464294
rect -8726 428614 -8106 464058
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 -8106 428614
rect -8726 428294 -8106 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 -8106 428294
rect -8726 392614 -8106 428058
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 -8106 392614
rect -8726 392294 -8106 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 -8106 392294
rect -8726 356614 -8106 392058
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 -8106 356614
rect -8726 356294 -8106 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 -8106 356294
rect -8726 320614 -8106 356058
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 -8106 320614
rect -8726 320294 -8106 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 -8106 320294
rect -8726 284614 -8106 320058
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 -8106 284614
rect -8726 284294 -8106 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 -8106 284294
rect -8726 248614 -8106 284058
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 -8106 248614
rect -8726 248294 -8106 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 -8106 248294
rect -8726 212614 -8106 248058
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 -8106 212614
rect -8726 212294 -8106 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 -8106 212294
rect -8726 176614 -8106 212058
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 -8106 176614
rect -8726 176294 -8106 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 -8106 176294
rect -8726 140614 -8106 176058
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 -8106 140614
rect -8726 140294 -8106 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 -8106 140294
rect -8726 104614 -8106 140058
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 -8106 104614
rect -8726 104294 -8106 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 -8106 104294
rect -8726 68614 -8106 104058
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 -8106 68614
rect -8726 68294 -8106 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 -8106 68294
rect -8726 32614 -8106 68058
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 -8106 32614
rect -8726 32294 -8106 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 -8106 32294
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 13574 710598
rect 12954 710278 13574 710362
rect 12954 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 13574 710278
rect -7766 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 -7146 698614
rect -7766 698294 -7146 698378
rect -7766 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 -7146 698294
rect -7766 662614 -7146 698058
rect -7766 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 -7146 662614
rect -7766 662294 -7146 662378
rect -7766 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 -7146 662294
rect -7766 626614 -7146 662058
rect -7766 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 -7146 626614
rect -7766 626294 -7146 626378
rect -7766 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 -7146 626294
rect -7766 590614 -7146 626058
rect -7766 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 -7146 590614
rect -7766 590294 -7146 590378
rect -7766 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 -7146 590294
rect -7766 554614 -7146 590058
rect -7766 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 -7146 554614
rect -7766 554294 -7146 554378
rect -7766 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 -7146 554294
rect -7766 518614 -7146 554058
rect -7766 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 -7146 518614
rect -7766 518294 -7146 518378
rect -7766 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 -7146 518294
rect -7766 482614 -7146 518058
rect -7766 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 -7146 482614
rect -7766 482294 -7146 482378
rect -7766 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 -7146 482294
rect -7766 446614 -7146 482058
rect -7766 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 -7146 446614
rect -7766 446294 -7146 446378
rect -7766 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 -7146 446294
rect -7766 410614 -7146 446058
rect -7766 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 -7146 410614
rect -7766 410294 -7146 410378
rect -7766 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 -7146 410294
rect -7766 374614 -7146 410058
rect -7766 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 -7146 374614
rect -7766 374294 -7146 374378
rect -7766 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 -7146 374294
rect -7766 338614 -7146 374058
rect -7766 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 -7146 338614
rect -7766 338294 -7146 338378
rect -7766 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 -7146 338294
rect -7766 302614 -7146 338058
rect -7766 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 -7146 302614
rect -7766 302294 -7146 302378
rect -7766 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 -7146 302294
rect -7766 266614 -7146 302058
rect -7766 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 -7146 266614
rect -7766 266294 -7146 266378
rect -7766 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 -7146 266294
rect -7766 230614 -7146 266058
rect -7766 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 -7146 230614
rect -7766 230294 -7146 230378
rect -7766 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 -7146 230294
rect -7766 194614 -7146 230058
rect -7766 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 -7146 194614
rect -7766 194294 -7146 194378
rect -7766 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 -7146 194294
rect -7766 158614 -7146 194058
rect -7766 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 -7146 158614
rect -7766 158294 -7146 158378
rect -7766 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 -7146 158294
rect -7766 122614 -7146 158058
rect -7766 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 -7146 122614
rect -7766 122294 -7146 122378
rect -7766 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 -7146 122294
rect -7766 86614 -7146 122058
rect -7766 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 -7146 86614
rect -7766 86294 -7146 86378
rect -7766 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 -7146 86294
rect -7766 50614 -7146 86058
rect -7766 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 -7146 50614
rect -7766 50294 -7146 50378
rect -7766 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 -7146 50294
rect -7766 14614 -7146 50058
rect -7766 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 -7146 14614
rect -7766 14294 -7146 14378
rect -7766 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 -7146 14294
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 676894 -6186 709082
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 -6186 676894
rect -6806 676574 -6186 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 -6186 676574
rect -6806 640894 -6186 676338
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 -6186 640894
rect -6806 640574 -6186 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 -6186 640574
rect -6806 604894 -6186 640338
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 -6186 604894
rect -6806 604574 -6186 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 -6186 604574
rect -6806 568894 -6186 604338
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 -6186 568894
rect -6806 568574 -6186 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 -6186 568574
rect -6806 532894 -6186 568338
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 -6186 532894
rect -6806 532574 -6186 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 -6186 532574
rect -6806 496894 -6186 532338
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 -6186 496894
rect -6806 496574 -6186 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 -6186 496574
rect -6806 460894 -6186 496338
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 -6186 460894
rect -6806 460574 -6186 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 -6186 460574
rect -6806 424894 -6186 460338
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 -6186 424894
rect -6806 424574 -6186 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 -6186 424574
rect -6806 388894 -6186 424338
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 -6186 388894
rect -6806 388574 -6186 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 -6186 388574
rect -6806 352894 -6186 388338
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 -6186 352894
rect -6806 352574 -6186 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 -6186 352574
rect -6806 316894 -6186 352338
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 -6186 316894
rect -6806 316574 -6186 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 -6186 316574
rect -6806 280894 -6186 316338
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 -6186 280894
rect -6806 280574 -6186 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 -6186 280574
rect -6806 244894 -6186 280338
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 -6186 244894
rect -6806 244574 -6186 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 -6186 244574
rect -6806 208894 -6186 244338
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 -6186 208894
rect -6806 208574 -6186 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 -6186 208574
rect -6806 172894 -6186 208338
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 -6186 172894
rect -6806 172574 -6186 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 -6186 172574
rect -6806 136894 -6186 172338
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 -6186 136894
rect -6806 136574 -6186 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 -6186 136574
rect -6806 100894 -6186 136338
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 -6186 100894
rect -6806 100574 -6186 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 -6186 100574
rect -6806 64894 -6186 100338
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 -6186 64894
rect -6806 64574 -6186 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 -6186 64574
rect -6806 28894 -6186 64338
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 -6186 28894
rect -6806 28574 -6186 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 -6186 28574
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 9854 708678
rect 9234 708358 9854 708442
rect 9234 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 9854 708358
rect -5846 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 -5226 694894
rect -5846 694574 -5226 694658
rect -5846 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 -5226 694574
rect -5846 658894 -5226 694338
rect -5846 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 -5226 658894
rect -5846 658574 -5226 658658
rect -5846 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 -5226 658574
rect -5846 622894 -5226 658338
rect -5846 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 -5226 622894
rect -5846 622574 -5226 622658
rect -5846 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 -5226 622574
rect -5846 586894 -5226 622338
rect -5846 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 -5226 586894
rect -5846 586574 -5226 586658
rect -5846 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 -5226 586574
rect -5846 550894 -5226 586338
rect -5846 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 -5226 550894
rect -5846 550574 -5226 550658
rect -5846 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 -5226 550574
rect -5846 514894 -5226 550338
rect -5846 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 -5226 514894
rect -5846 514574 -5226 514658
rect -5846 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 -5226 514574
rect -5846 478894 -5226 514338
rect -5846 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 -5226 478894
rect -5846 478574 -5226 478658
rect -5846 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 -5226 478574
rect -5846 442894 -5226 478338
rect -5846 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 -5226 442894
rect -5846 442574 -5226 442658
rect -5846 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 -5226 442574
rect -5846 406894 -5226 442338
rect -5846 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 -5226 406894
rect -5846 406574 -5226 406658
rect -5846 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 -5226 406574
rect -5846 370894 -5226 406338
rect -5846 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 -5226 370894
rect -5846 370574 -5226 370658
rect -5846 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 -5226 370574
rect -5846 334894 -5226 370338
rect -5846 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 -5226 334894
rect -5846 334574 -5226 334658
rect -5846 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 -5226 334574
rect -5846 298894 -5226 334338
rect -5846 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 -5226 298894
rect -5846 298574 -5226 298658
rect -5846 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 -5226 298574
rect -5846 262894 -5226 298338
rect -5846 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 -5226 262894
rect -5846 262574 -5226 262658
rect -5846 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 -5226 262574
rect -5846 226894 -5226 262338
rect -5846 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 -5226 226894
rect -5846 226574 -5226 226658
rect -5846 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 -5226 226574
rect -5846 190894 -5226 226338
rect -5846 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 -5226 190894
rect -5846 190574 -5226 190658
rect -5846 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 -5226 190574
rect -5846 154894 -5226 190338
rect -5846 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 -5226 154894
rect -5846 154574 -5226 154658
rect -5846 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 -5226 154574
rect -5846 118894 -5226 154338
rect -5846 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 -5226 118894
rect -5846 118574 -5226 118658
rect -5846 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 -5226 118574
rect -5846 82894 -5226 118338
rect -5846 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 -5226 82894
rect -5846 82574 -5226 82658
rect -5846 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 -5226 82574
rect -5846 46894 -5226 82338
rect -5846 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 -5226 46894
rect -5846 46574 -5226 46658
rect -5846 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 -5226 46574
rect -5846 10894 -5226 46338
rect -5846 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 -5226 10894
rect -5846 10574 -5226 10658
rect -5846 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 -5226 10574
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 673174 -4266 707162
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 -4266 673174
rect -4886 672854 -4266 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 -4266 672854
rect -4886 637174 -4266 672618
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 -4266 637174
rect -4886 636854 -4266 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 -4266 636854
rect -4886 601174 -4266 636618
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 -4266 601174
rect -4886 600854 -4266 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 -4266 600854
rect -4886 565174 -4266 600618
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 -4266 565174
rect -4886 564854 -4266 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 -4266 564854
rect -4886 529174 -4266 564618
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 -4266 529174
rect -4886 528854 -4266 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 -4266 528854
rect -4886 493174 -4266 528618
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 -4266 493174
rect -4886 492854 -4266 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 -4266 492854
rect -4886 457174 -4266 492618
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 -4266 457174
rect -4886 456854 -4266 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 -4266 456854
rect -4886 421174 -4266 456618
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 -4266 421174
rect -4886 420854 -4266 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 -4266 420854
rect -4886 385174 -4266 420618
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 -4266 385174
rect -4886 384854 -4266 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 -4266 384854
rect -4886 349174 -4266 384618
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 -4266 349174
rect -4886 348854 -4266 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 -4266 348854
rect -4886 313174 -4266 348618
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 -4266 313174
rect -4886 312854 -4266 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 -4266 312854
rect -4886 277174 -4266 312618
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 -4266 277174
rect -4886 276854 -4266 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 -4266 276854
rect -4886 241174 -4266 276618
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 -4266 241174
rect -4886 240854 -4266 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 -4266 240854
rect -4886 205174 -4266 240618
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 -4266 205174
rect -4886 204854 -4266 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 -4266 204854
rect -4886 169174 -4266 204618
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 -4266 169174
rect -4886 168854 -4266 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 -4266 168854
rect -4886 133174 -4266 168618
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 -4266 133174
rect -4886 132854 -4266 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 -4266 132854
rect -4886 97174 -4266 132618
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 -4266 97174
rect -4886 96854 -4266 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 -4266 96854
rect -4886 61174 -4266 96618
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 -4266 61174
rect -4886 60854 -4266 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 -4266 60854
rect -4886 25174 -4266 60618
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 -4266 25174
rect -4886 24854 -4266 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 -4266 24854
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 6134 706758
rect 5514 706438 6134 706522
rect 5514 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 6134 706438
rect -3926 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 -3306 691174
rect -3926 690854 -3306 690938
rect -3926 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 -3306 690854
rect -3926 655174 -3306 690618
rect -3926 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 -3306 655174
rect -3926 654854 -3306 654938
rect -3926 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 -3306 654854
rect -3926 619174 -3306 654618
rect -3926 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 -3306 619174
rect -3926 618854 -3306 618938
rect -3926 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 -3306 618854
rect -3926 583174 -3306 618618
rect -3926 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 -3306 583174
rect -3926 582854 -3306 582938
rect -3926 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 -3306 582854
rect -3926 547174 -3306 582618
rect -3926 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 -3306 547174
rect -3926 546854 -3306 546938
rect -3926 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 -3306 546854
rect -3926 511174 -3306 546618
rect -3926 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 -3306 511174
rect -3926 510854 -3306 510938
rect -3926 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 -3306 510854
rect -3926 475174 -3306 510618
rect -3926 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 -3306 475174
rect -3926 474854 -3306 474938
rect -3926 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 -3306 474854
rect -3926 439174 -3306 474618
rect -3926 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 -3306 439174
rect -3926 438854 -3306 438938
rect -3926 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 -3306 438854
rect -3926 403174 -3306 438618
rect -3926 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 -3306 403174
rect -3926 402854 -3306 402938
rect -3926 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 -3306 402854
rect -3926 367174 -3306 402618
rect -3926 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 -3306 367174
rect -3926 366854 -3306 366938
rect -3926 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 -3306 366854
rect -3926 331174 -3306 366618
rect -3926 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 -3306 331174
rect -3926 330854 -3306 330938
rect -3926 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 -3306 330854
rect -3926 295174 -3306 330618
rect -3926 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 -3306 295174
rect -3926 294854 -3306 294938
rect -3926 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 -3306 294854
rect -3926 259174 -3306 294618
rect -3926 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 -3306 259174
rect -3926 258854 -3306 258938
rect -3926 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 -3306 258854
rect -3926 223174 -3306 258618
rect -3926 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 -3306 223174
rect -3926 222854 -3306 222938
rect -3926 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 -3306 222854
rect -3926 187174 -3306 222618
rect -3926 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 -3306 187174
rect -3926 186854 -3306 186938
rect -3926 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 -3306 186854
rect -3926 151174 -3306 186618
rect -3926 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 -3306 151174
rect -3926 150854 -3306 150938
rect -3926 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 -3306 150854
rect -3926 115174 -3306 150618
rect -3926 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 -3306 115174
rect -3926 114854 -3306 114938
rect -3926 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 -3306 114854
rect -3926 79174 -3306 114618
rect -3926 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 -3306 79174
rect -3926 78854 -3306 78938
rect -3926 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 -3306 78854
rect -3926 43174 -3306 78618
rect -3926 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 -3306 43174
rect -3926 42854 -3306 42938
rect -3926 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 -3306 42854
rect -3926 7174 -3306 42618
rect -3926 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 -3306 7174
rect -3926 6854 -3306 6938
rect -3926 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 -3306 6854
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 702000 2414 704282
rect 5514 702000 6134 706202
rect 9234 702000 9854 708122
rect 12954 702000 13574 710042
rect 30954 711558 31574 711590
rect 30954 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 31574 711558
rect 30954 711238 31574 711322
rect 30954 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 31574 711238
rect 27234 709638 27854 709670
rect 27234 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 27854 709638
rect 27234 709318 27854 709402
rect 27234 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 27854 709318
rect 23514 707718 24134 707750
rect 23514 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 24134 707718
rect 23514 707398 24134 707482
rect 23514 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 24134 707398
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 19794 702000 20414 705242
rect 23514 702000 24134 707162
rect 27234 702000 27854 709082
rect 30954 702000 31574 711002
rect 48954 710598 49574 711590
rect 48954 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 49574 710598
rect 48954 710278 49574 710362
rect 48954 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 49574 710278
rect 45234 708678 45854 709670
rect 45234 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 45854 708678
rect 45234 708358 45854 708442
rect 45234 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 45854 708358
rect 41514 706758 42134 707750
rect 41514 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 42134 706758
rect 41514 706438 42134 706522
rect 41514 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 42134 706438
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 702000 38414 704282
rect 41514 702000 42134 706202
rect 45234 702000 45854 708122
rect 48954 702000 49574 710042
rect 66954 711558 67574 711590
rect 66954 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 67574 711558
rect 66954 711238 67574 711322
rect 66954 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 67574 711238
rect 63234 709638 63854 709670
rect 63234 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 63854 709638
rect 63234 709318 63854 709402
rect 63234 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 63854 709318
rect 59514 707718 60134 707750
rect 59514 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 60134 707718
rect 59514 707398 60134 707482
rect 59514 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 60134 707398
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 702000 56414 705242
rect 59514 702000 60134 707162
rect 63234 702000 63854 709082
rect 66954 702000 67574 711002
rect 84954 710598 85574 711590
rect 84954 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 85574 710598
rect 84954 710278 85574 710362
rect 84954 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 85574 710278
rect 81234 708678 81854 709670
rect 81234 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 81854 708678
rect 81234 708358 81854 708442
rect 81234 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 81854 708358
rect 77514 706758 78134 707750
rect 77514 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 78134 706758
rect 77514 706438 78134 706522
rect 77514 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 78134 706438
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 702000 74414 704282
rect 77514 702000 78134 706202
rect 81234 702000 81854 708122
rect 84954 702000 85574 710042
rect 102954 711558 103574 711590
rect 102954 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 103574 711558
rect 102954 711238 103574 711322
rect 102954 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 103574 711238
rect 99234 709638 99854 709670
rect 99234 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 99854 709638
rect 99234 709318 99854 709402
rect 99234 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 99854 709318
rect 95514 707718 96134 707750
rect 95514 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 96134 707718
rect 95514 707398 96134 707482
rect 95514 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 96134 707398
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 702000 92414 705242
rect 95514 702000 96134 707162
rect 99234 702000 99854 709082
rect 102954 702000 103574 711002
rect 120954 710598 121574 711590
rect 120954 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 121574 710598
rect 120954 710278 121574 710362
rect 120954 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 121574 710278
rect 117234 708678 117854 709670
rect 117234 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 117854 708678
rect 117234 708358 117854 708442
rect 117234 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 117854 708358
rect 113514 706758 114134 707750
rect 113514 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 114134 706758
rect 113514 706438 114134 706522
rect 113514 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 114134 706438
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 702000 110414 704282
rect 113514 702000 114134 706202
rect 117234 702000 117854 708122
rect 120954 702000 121574 710042
rect 138954 711558 139574 711590
rect 138954 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 139574 711558
rect 138954 711238 139574 711322
rect 138954 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 139574 711238
rect 135234 709638 135854 709670
rect 135234 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 135854 709638
rect 135234 709318 135854 709402
rect 135234 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 135854 709318
rect 131514 707718 132134 707750
rect 131514 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 132134 707718
rect 131514 707398 132134 707482
rect 131514 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 132134 707398
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 127794 702000 128414 705242
rect 131514 702000 132134 707162
rect 135234 702000 135854 709082
rect 138954 702000 139574 711002
rect 156954 710598 157574 711590
rect 156954 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 157574 710598
rect 156954 710278 157574 710362
rect 156954 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 157574 710278
rect 153234 708678 153854 709670
rect 153234 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 153854 708678
rect 153234 708358 153854 708442
rect 153234 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 153854 708358
rect 149514 706758 150134 707750
rect 149514 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 150134 706758
rect 149514 706438 150134 706522
rect 149514 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 150134 706438
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 702000 146414 704282
rect 149514 702000 150134 706202
rect 153234 702000 153854 708122
rect 156954 702000 157574 710042
rect 174954 711558 175574 711590
rect 174954 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 175574 711558
rect 174954 711238 175574 711322
rect 174954 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 175574 711238
rect 171234 709638 171854 709670
rect 171234 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 171854 709638
rect 171234 709318 171854 709402
rect 171234 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 171854 709318
rect 167514 707718 168134 707750
rect 167514 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 168134 707718
rect 167514 707398 168134 707482
rect 167514 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 168134 707398
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 702000 164414 705242
rect 167514 702000 168134 707162
rect 171234 702000 171854 709082
rect 174954 702000 175574 711002
rect 192954 710598 193574 711590
rect 192954 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 193574 710598
rect 192954 710278 193574 710362
rect 192954 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 193574 710278
rect 189234 708678 189854 709670
rect 189234 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 189854 708678
rect 189234 708358 189854 708442
rect 189234 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 189854 708358
rect 185514 706758 186134 707750
rect 185514 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 186134 706758
rect 185514 706438 186134 706522
rect 185514 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 186134 706438
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 702000 182414 704282
rect 185514 702000 186134 706202
rect 189234 702000 189854 708122
rect 192954 702000 193574 710042
rect 210954 711558 211574 711590
rect 210954 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 211574 711558
rect 210954 711238 211574 711322
rect 210954 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 211574 711238
rect 207234 709638 207854 709670
rect 207234 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 207854 709638
rect 207234 709318 207854 709402
rect 207234 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 207854 709318
rect 203514 707718 204134 707750
rect 203514 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 204134 707718
rect 203514 707398 204134 707482
rect 203514 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 204134 707398
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 702000 200414 705242
rect 203514 702000 204134 707162
rect 207234 702000 207854 709082
rect 210954 702000 211574 711002
rect 228954 710598 229574 711590
rect 228954 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 229574 710598
rect 228954 710278 229574 710362
rect 228954 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 229574 710278
rect 225234 708678 225854 709670
rect 225234 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 225854 708678
rect 225234 708358 225854 708442
rect 225234 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 225854 708358
rect 221514 706758 222134 707750
rect 221514 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 222134 706758
rect 221514 706438 222134 706522
rect 221514 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 222134 706438
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 702000 218414 704282
rect 221514 702000 222134 706202
rect 225234 702000 225854 708122
rect 228954 702000 229574 710042
rect 246954 711558 247574 711590
rect 246954 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 247574 711558
rect 246954 711238 247574 711322
rect 246954 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 247574 711238
rect 243234 709638 243854 709670
rect 243234 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 243854 709638
rect 243234 709318 243854 709402
rect 243234 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 243854 709318
rect 239514 707718 240134 707750
rect 239514 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 240134 707718
rect 239514 707398 240134 707482
rect 239514 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 240134 707398
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 235794 702000 236414 705242
rect 239514 702000 240134 707162
rect 243234 702000 243854 709082
rect 246954 702000 247574 711002
rect 264954 710598 265574 711590
rect 264954 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 265574 710598
rect 264954 710278 265574 710362
rect 264954 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 265574 710278
rect 261234 708678 261854 709670
rect 261234 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 261854 708678
rect 261234 708358 261854 708442
rect 261234 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 261854 708358
rect 257514 706758 258134 707750
rect 257514 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 258134 706758
rect 257514 706438 258134 706522
rect 257514 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 258134 706438
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 702000 254414 704282
rect 257514 702000 258134 706202
rect 261234 702000 261854 708122
rect 264954 702000 265574 710042
rect 282954 711558 283574 711590
rect 282954 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 283574 711558
rect 282954 711238 283574 711322
rect 282954 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 283574 711238
rect 279234 709638 279854 709670
rect 279234 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 279854 709638
rect 279234 709318 279854 709402
rect 279234 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 279854 709318
rect 275514 707718 276134 707750
rect 275514 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 276134 707718
rect 275514 707398 276134 707482
rect 275514 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 276134 707398
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 271794 702000 272414 705242
rect 275514 702000 276134 707162
rect 279234 702000 279854 709082
rect 282954 702000 283574 711002
rect 300954 710598 301574 711590
rect 300954 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 301574 710598
rect 300954 710278 301574 710362
rect 300954 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 301574 710278
rect 297234 708678 297854 709670
rect 297234 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 297854 708678
rect 297234 708358 297854 708442
rect 297234 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 297854 708358
rect 293514 706758 294134 707750
rect 293514 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 294134 706758
rect 293514 706438 294134 706522
rect 293514 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 294134 706438
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 702000 290414 704282
rect 293514 702000 294134 706202
rect 297234 702000 297854 708122
rect 300954 702000 301574 710042
rect 318954 711558 319574 711590
rect 318954 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 319574 711558
rect 318954 711238 319574 711322
rect 318954 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 319574 711238
rect 315234 709638 315854 709670
rect 315234 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 315854 709638
rect 315234 709318 315854 709402
rect 315234 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 315854 709318
rect 311514 707718 312134 707750
rect 311514 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 312134 707718
rect 311514 707398 312134 707482
rect 311514 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 312134 707398
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 702000 308414 705242
rect 311514 702000 312134 707162
rect 315234 702000 315854 709082
rect 318954 702000 319574 711002
rect 336954 710598 337574 711590
rect 336954 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 337574 710598
rect 336954 710278 337574 710362
rect 336954 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 337574 710278
rect 333234 708678 333854 709670
rect 333234 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 333854 708678
rect 333234 708358 333854 708442
rect 333234 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 333854 708358
rect 329514 706758 330134 707750
rect 329514 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 330134 706758
rect 329514 706438 330134 706522
rect 329514 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 330134 706438
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 702000 326414 704282
rect 329514 702000 330134 706202
rect 333234 702000 333854 708122
rect 336954 702000 337574 710042
rect 354954 711558 355574 711590
rect 354954 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 355574 711558
rect 354954 711238 355574 711322
rect 354954 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 355574 711238
rect 351234 709638 351854 709670
rect 351234 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 351854 709638
rect 351234 709318 351854 709402
rect 351234 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 351854 709318
rect 347514 707718 348134 707750
rect 347514 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 348134 707718
rect 347514 707398 348134 707482
rect 347514 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 348134 707398
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 343794 702000 344414 705242
rect 347514 702000 348134 707162
rect 351234 702000 351854 709082
rect 354954 702000 355574 711002
rect 372954 710598 373574 711590
rect 372954 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 373574 710598
rect 372954 710278 373574 710362
rect 372954 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 373574 710278
rect 369234 708678 369854 709670
rect 369234 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 369854 708678
rect 369234 708358 369854 708442
rect 369234 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 369854 708358
rect 365514 706758 366134 707750
rect 365514 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 366134 706758
rect 365514 706438 366134 706522
rect 365514 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 366134 706438
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 702000 362414 704282
rect 365514 702000 366134 706202
rect 369234 702000 369854 708122
rect 372954 702000 373574 710042
rect 390954 711558 391574 711590
rect 390954 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 391574 711558
rect 390954 711238 391574 711322
rect 390954 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 391574 711238
rect 387234 709638 387854 709670
rect 387234 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 387854 709638
rect 387234 709318 387854 709402
rect 387234 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 387854 709318
rect 383514 707718 384134 707750
rect 383514 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 384134 707718
rect 383514 707398 384134 707482
rect 383514 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 384134 707398
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 379794 702000 380414 705242
rect 383514 702000 384134 707162
rect 387234 702000 387854 709082
rect 390954 702000 391574 711002
rect 408954 710598 409574 711590
rect 408954 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 409574 710598
rect 408954 710278 409574 710362
rect 408954 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 409574 710278
rect 405234 708678 405854 709670
rect 405234 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 405854 708678
rect 405234 708358 405854 708442
rect 405234 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 405854 708358
rect 401514 706758 402134 707750
rect 401514 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 402134 706758
rect 401514 706438 402134 706522
rect 401514 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 402134 706438
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 702000 398414 704282
rect 401514 702000 402134 706202
rect 405234 702000 405854 708122
rect 408954 702000 409574 710042
rect 426954 711558 427574 711590
rect 426954 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 427574 711558
rect 426954 711238 427574 711322
rect 426954 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 427574 711238
rect 423234 709638 423854 709670
rect 423234 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 423854 709638
rect 423234 709318 423854 709402
rect 423234 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 423854 709318
rect 419514 707718 420134 707750
rect 419514 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 420134 707718
rect 419514 707398 420134 707482
rect 419514 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 420134 707398
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 415794 702000 416414 705242
rect 419514 702000 420134 707162
rect 423234 702000 423854 709082
rect 426954 702000 427574 711002
rect 444954 710598 445574 711590
rect 444954 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 445574 710598
rect 444954 710278 445574 710362
rect 444954 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 445574 710278
rect 441234 708678 441854 709670
rect 441234 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 441854 708678
rect 441234 708358 441854 708442
rect 441234 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 441854 708358
rect 437514 706758 438134 707750
rect 437514 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 438134 706758
rect 437514 706438 438134 706522
rect 437514 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 438134 706438
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 702000 434414 704282
rect 437514 702000 438134 706202
rect 441234 702000 441854 708122
rect 444954 702000 445574 710042
rect 462954 711558 463574 711590
rect 462954 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 463574 711558
rect 462954 711238 463574 711322
rect 462954 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 463574 711238
rect 459234 709638 459854 709670
rect 459234 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 459854 709638
rect 459234 709318 459854 709402
rect 459234 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 459854 709318
rect 455514 707718 456134 707750
rect 455514 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 456134 707718
rect 455514 707398 456134 707482
rect 455514 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 456134 707398
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 702000 452414 705242
rect 455514 702000 456134 707162
rect 459234 702000 459854 709082
rect 462954 702000 463574 711002
rect 480954 710598 481574 711590
rect 480954 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 481574 710598
rect 480954 710278 481574 710362
rect 480954 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 481574 710278
rect 477234 708678 477854 709670
rect 477234 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 477854 708678
rect 477234 708358 477854 708442
rect 477234 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 477854 708358
rect 473514 706758 474134 707750
rect 473514 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 474134 706758
rect 473514 706438 474134 706522
rect 473514 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 474134 706438
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 702000 470414 704282
rect 473514 702000 474134 706202
rect 477234 702000 477854 708122
rect 480954 702000 481574 710042
rect 498954 711558 499574 711590
rect 498954 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 499574 711558
rect 498954 711238 499574 711322
rect 498954 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 499574 711238
rect 495234 709638 495854 709670
rect 495234 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 495854 709638
rect 495234 709318 495854 709402
rect 495234 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 495854 709318
rect 491514 707718 492134 707750
rect 491514 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 492134 707718
rect 491514 707398 492134 707482
rect 491514 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 492134 707398
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 487794 702000 488414 705242
rect 491514 702000 492134 707162
rect 495234 702000 495854 709082
rect 498954 702000 499574 711002
rect 516954 710598 517574 711590
rect 516954 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 517574 710598
rect 516954 710278 517574 710362
rect 516954 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 517574 710278
rect 513234 708678 513854 709670
rect 513234 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 513854 708678
rect 513234 708358 513854 708442
rect 513234 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 513854 708358
rect 509514 706758 510134 707750
rect 509514 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 510134 706758
rect 509514 706438 510134 706522
rect 509514 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 510134 706438
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 702000 506414 704282
rect 509514 702000 510134 706202
rect 513234 702000 513854 708122
rect 516954 702000 517574 710042
rect 534954 711558 535574 711590
rect 534954 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 535574 711558
rect 534954 711238 535574 711322
rect 534954 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 535574 711238
rect 531234 709638 531854 709670
rect 531234 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 531854 709638
rect 531234 709318 531854 709402
rect 531234 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 531854 709318
rect 527514 707718 528134 707750
rect 527514 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 528134 707718
rect 527514 707398 528134 707482
rect 527514 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 528134 707398
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 702000 524414 705242
rect 527514 702000 528134 707162
rect 531234 702000 531854 709082
rect 534954 702000 535574 711002
rect 552954 710598 553574 711590
rect 552954 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 553574 710598
rect 552954 710278 553574 710362
rect 552954 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 553574 710278
rect 549234 708678 549854 709670
rect 549234 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 549854 708678
rect 549234 708358 549854 708442
rect 549234 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 549854 708358
rect 545514 706758 546134 707750
rect 545514 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 546134 706758
rect 545514 706438 546134 706522
rect 545514 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 546134 706438
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 702000 542414 704282
rect 545514 702000 546134 706202
rect 549234 702000 549854 708122
rect 552954 702000 553574 710042
rect 570954 711558 571574 711590
rect 570954 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 571574 711558
rect 570954 711238 571574 711322
rect 570954 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 571574 711238
rect 567234 709638 567854 709670
rect 567234 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 567854 709638
rect 567234 709318 567854 709402
rect 567234 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 567854 709318
rect 563514 707718 564134 707750
rect 563514 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 564134 707718
rect 563514 707398 564134 707482
rect 563514 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 564134 707398
rect 559794 705798 560414 705830
rect 559794 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 560414 705798
rect 559794 705478 560414 705562
rect 559794 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 560414 705478
rect 559794 702000 560414 705242
rect 563514 702000 564134 707162
rect 13859 699412 13925 699413
rect 13859 699348 13860 699412
rect 13924 699348 13925 699412
rect 13859 699347 13925 699348
rect 21403 699412 21469 699413
rect 21403 699348 21404 699412
rect 21468 699348 21469 699412
rect 21403 699347 21469 699348
rect 69979 699412 70045 699413
rect 69979 699348 69980 699412
rect 70044 699348 70045 699412
rect 69979 699347 70045 699348
rect 82123 699412 82189 699413
rect 82123 699348 82124 699412
rect 82188 699348 82189 699412
rect 82123 699347 82189 699348
rect 418659 699412 418725 699413
rect 418659 699348 418660 699412
rect 418724 699348 418725 699412
rect 418659 699347 418725 699348
rect 423627 699412 423693 699413
rect 423627 699348 423628 699412
rect 423692 699348 423693 699412
rect 423627 699347 423693 699348
rect 433379 699412 433445 699413
rect 433379 699348 433380 699412
rect 433444 699348 433445 699412
rect 433379 699347 433445 699348
rect 448099 699412 448165 699413
rect 448099 699348 448100 699412
rect 448164 699348 448165 699412
rect 448099 699347 448165 699348
rect 465763 699412 465829 699413
rect 465763 699348 465764 699412
rect 465828 699348 465829 699412
rect 465763 699347 465829 699348
rect 477539 699412 477605 699413
rect 477539 699348 477540 699412
rect 477604 699348 477605 699412
rect 477539 699347 477605 699348
rect 539915 699412 539981 699413
rect 539915 699348 539916 699412
rect 539980 699348 539981 699412
rect 539915 699347 539981 699348
rect 13862 698325 13922 699347
rect 21406 698461 21466 699347
rect 69982 698733 70042 699347
rect 82126 698869 82186 699347
rect 82123 698868 82189 698869
rect 82123 698804 82124 698868
rect 82188 698804 82189 698868
rect 82123 698803 82189 698804
rect 69979 698732 70045 698733
rect 69979 698668 69980 698732
rect 70044 698668 70045 698732
rect 69979 698667 70045 698668
rect 21403 698460 21469 698461
rect 21403 698396 21404 698460
rect 21468 698396 21469 698460
rect 21403 698395 21469 698396
rect 13859 698324 13925 698325
rect 13859 698260 13860 698324
rect 13924 698260 13925 698324
rect 13859 698259 13925 698260
rect 418662 697781 418722 699347
rect 418843 699276 418909 699277
rect 418843 699212 418844 699276
rect 418908 699212 418909 699276
rect 418843 699211 418909 699212
rect 418846 697781 418906 699211
rect 423630 698189 423690 699347
rect 423627 698188 423693 698189
rect 423627 698124 423628 698188
rect 423692 698124 423693 698188
rect 423627 698123 423693 698124
rect 433382 698053 433442 699347
rect 433379 698052 433445 698053
rect 433379 697988 433380 698052
rect 433444 697988 433445 698052
rect 433379 697987 433445 697988
rect 448102 697917 448162 699347
rect 465766 699005 465826 699347
rect 465763 699004 465829 699005
rect 465763 698940 465764 699004
rect 465828 698940 465829 699004
rect 465763 698939 465829 698940
rect 448099 697916 448165 697917
rect 448099 697852 448100 697916
rect 448164 697852 448165 697916
rect 448099 697851 448165 697852
rect 418659 697780 418725 697781
rect 418659 697716 418660 697780
rect 418724 697716 418725 697780
rect 418659 697715 418725 697716
rect 418843 697780 418909 697781
rect 418843 697716 418844 697780
rect 418908 697716 418909 697780
rect 418843 697715 418909 697716
rect 477542 697645 477602 699347
rect 539918 698597 539978 699347
rect 539915 698596 539981 698597
rect 539915 698532 539916 698596
rect 539980 698532 539981 698596
rect 539915 698531 539981 698532
rect 477539 697644 477605 697645
rect 477539 697580 477540 697644
rect 477604 697580 477605 697644
rect 477539 697579 477605 697580
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect 8208 687454 8528 687486
rect 8208 687218 8250 687454
rect 8486 687218 8528 687454
rect 8208 687134 8528 687218
rect 8208 686898 8250 687134
rect 8486 686898 8528 687134
rect 8208 686866 8528 686898
rect 38928 687454 39248 687486
rect 38928 687218 38970 687454
rect 39206 687218 39248 687454
rect 38928 687134 39248 687218
rect 38928 686898 38970 687134
rect 39206 686898 39248 687134
rect 38928 686866 39248 686898
rect 69648 687454 69968 687486
rect 69648 687218 69690 687454
rect 69926 687218 69968 687454
rect 69648 687134 69968 687218
rect 69648 686898 69690 687134
rect 69926 686898 69968 687134
rect 69648 686866 69968 686898
rect 100368 687454 100688 687486
rect 100368 687218 100410 687454
rect 100646 687218 100688 687454
rect 100368 687134 100688 687218
rect 100368 686898 100410 687134
rect 100646 686898 100688 687134
rect 100368 686866 100688 686898
rect 131088 687454 131408 687486
rect 131088 687218 131130 687454
rect 131366 687218 131408 687454
rect 131088 687134 131408 687218
rect 131088 686898 131130 687134
rect 131366 686898 131408 687134
rect 131088 686866 131408 686898
rect 161808 687454 162128 687486
rect 161808 687218 161850 687454
rect 162086 687218 162128 687454
rect 161808 687134 162128 687218
rect 161808 686898 161850 687134
rect 162086 686898 162128 687134
rect 161808 686866 162128 686898
rect 192528 687454 192848 687486
rect 192528 687218 192570 687454
rect 192806 687218 192848 687454
rect 192528 687134 192848 687218
rect 192528 686898 192570 687134
rect 192806 686898 192848 687134
rect 192528 686866 192848 686898
rect 223248 687454 223568 687486
rect 223248 687218 223290 687454
rect 223526 687218 223568 687454
rect 223248 687134 223568 687218
rect 223248 686898 223290 687134
rect 223526 686898 223568 687134
rect 223248 686866 223568 686898
rect 253968 687454 254288 687486
rect 253968 687218 254010 687454
rect 254246 687218 254288 687454
rect 253968 687134 254288 687218
rect 253968 686898 254010 687134
rect 254246 686898 254288 687134
rect 253968 686866 254288 686898
rect 284688 687454 285008 687486
rect 284688 687218 284730 687454
rect 284966 687218 285008 687454
rect 284688 687134 285008 687218
rect 284688 686898 284730 687134
rect 284966 686898 285008 687134
rect 284688 686866 285008 686898
rect 315408 687454 315728 687486
rect 315408 687218 315450 687454
rect 315686 687218 315728 687454
rect 315408 687134 315728 687218
rect 315408 686898 315450 687134
rect 315686 686898 315728 687134
rect 315408 686866 315728 686898
rect 346128 687454 346448 687486
rect 346128 687218 346170 687454
rect 346406 687218 346448 687454
rect 346128 687134 346448 687218
rect 346128 686898 346170 687134
rect 346406 686898 346448 687134
rect 346128 686866 346448 686898
rect 376848 687454 377168 687486
rect 376848 687218 376890 687454
rect 377126 687218 377168 687454
rect 376848 687134 377168 687218
rect 376848 686898 376890 687134
rect 377126 686898 377168 687134
rect 376848 686866 377168 686898
rect 407568 687454 407888 687486
rect 407568 687218 407610 687454
rect 407846 687218 407888 687454
rect 407568 687134 407888 687218
rect 407568 686898 407610 687134
rect 407846 686898 407888 687134
rect 407568 686866 407888 686898
rect 438288 687454 438608 687486
rect 438288 687218 438330 687454
rect 438566 687218 438608 687454
rect 438288 687134 438608 687218
rect 438288 686898 438330 687134
rect 438566 686898 438608 687134
rect 438288 686866 438608 686898
rect 469008 687454 469328 687486
rect 469008 687218 469050 687454
rect 469286 687218 469328 687454
rect 469008 687134 469328 687218
rect 469008 686898 469050 687134
rect 469286 686898 469328 687134
rect 469008 686866 469328 686898
rect 499728 687454 500048 687486
rect 499728 687218 499770 687454
rect 500006 687218 500048 687454
rect 499728 687134 500048 687218
rect 499728 686898 499770 687134
rect 500006 686898 500048 687134
rect 499728 686866 500048 686898
rect 530448 687454 530768 687486
rect 530448 687218 530490 687454
rect 530726 687218 530768 687454
rect 530448 687134 530768 687218
rect 530448 686898 530490 687134
rect 530726 686898 530768 687134
rect 530448 686866 530768 686898
rect 561168 687454 561488 687486
rect 561168 687218 561210 687454
rect 561446 687218 561488 687454
rect 561168 687134 561488 687218
rect 561168 686898 561210 687134
rect 561446 686898 561488 687134
rect 561168 686866 561488 686898
rect 567234 676894 567854 709082
rect 567234 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 567854 676894
rect 567234 676574 567854 676658
rect 567234 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 567854 676574
rect 23568 669454 23888 669486
rect 23568 669218 23610 669454
rect 23846 669218 23888 669454
rect 23568 669134 23888 669218
rect 23568 668898 23610 669134
rect 23846 668898 23888 669134
rect 23568 668866 23888 668898
rect 54288 669454 54608 669486
rect 54288 669218 54330 669454
rect 54566 669218 54608 669454
rect 54288 669134 54608 669218
rect 54288 668898 54330 669134
rect 54566 668898 54608 669134
rect 54288 668866 54608 668898
rect 85008 669454 85328 669486
rect 85008 669218 85050 669454
rect 85286 669218 85328 669454
rect 85008 669134 85328 669218
rect 85008 668898 85050 669134
rect 85286 668898 85328 669134
rect 85008 668866 85328 668898
rect 115728 669454 116048 669486
rect 115728 669218 115770 669454
rect 116006 669218 116048 669454
rect 115728 669134 116048 669218
rect 115728 668898 115770 669134
rect 116006 668898 116048 669134
rect 115728 668866 116048 668898
rect 146448 669454 146768 669486
rect 146448 669218 146490 669454
rect 146726 669218 146768 669454
rect 146448 669134 146768 669218
rect 146448 668898 146490 669134
rect 146726 668898 146768 669134
rect 146448 668866 146768 668898
rect 177168 669454 177488 669486
rect 177168 669218 177210 669454
rect 177446 669218 177488 669454
rect 177168 669134 177488 669218
rect 177168 668898 177210 669134
rect 177446 668898 177488 669134
rect 177168 668866 177488 668898
rect 207888 669454 208208 669486
rect 207888 669218 207930 669454
rect 208166 669218 208208 669454
rect 207888 669134 208208 669218
rect 207888 668898 207930 669134
rect 208166 668898 208208 669134
rect 207888 668866 208208 668898
rect 238608 669454 238928 669486
rect 238608 669218 238650 669454
rect 238886 669218 238928 669454
rect 238608 669134 238928 669218
rect 238608 668898 238650 669134
rect 238886 668898 238928 669134
rect 238608 668866 238928 668898
rect 269328 669454 269648 669486
rect 269328 669218 269370 669454
rect 269606 669218 269648 669454
rect 269328 669134 269648 669218
rect 269328 668898 269370 669134
rect 269606 668898 269648 669134
rect 269328 668866 269648 668898
rect 300048 669454 300368 669486
rect 300048 669218 300090 669454
rect 300326 669218 300368 669454
rect 300048 669134 300368 669218
rect 300048 668898 300090 669134
rect 300326 668898 300368 669134
rect 300048 668866 300368 668898
rect 330768 669454 331088 669486
rect 330768 669218 330810 669454
rect 331046 669218 331088 669454
rect 330768 669134 331088 669218
rect 330768 668898 330810 669134
rect 331046 668898 331088 669134
rect 330768 668866 331088 668898
rect 361488 669454 361808 669486
rect 361488 669218 361530 669454
rect 361766 669218 361808 669454
rect 361488 669134 361808 669218
rect 361488 668898 361530 669134
rect 361766 668898 361808 669134
rect 361488 668866 361808 668898
rect 392208 669454 392528 669486
rect 392208 669218 392250 669454
rect 392486 669218 392528 669454
rect 392208 669134 392528 669218
rect 392208 668898 392250 669134
rect 392486 668898 392528 669134
rect 392208 668866 392528 668898
rect 422928 669454 423248 669486
rect 422928 669218 422970 669454
rect 423206 669218 423248 669454
rect 422928 669134 423248 669218
rect 422928 668898 422970 669134
rect 423206 668898 423248 669134
rect 422928 668866 423248 668898
rect 453648 669454 453968 669486
rect 453648 669218 453690 669454
rect 453926 669218 453968 669454
rect 453648 669134 453968 669218
rect 453648 668898 453690 669134
rect 453926 668898 453968 669134
rect 453648 668866 453968 668898
rect 484368 669454 484688 669486
rect 484368 669218 484410 669454
rect 484646 669218 484688 669454
rect 484368 669134 484688 669218
rect 484368 668898 484410 669134
rect 484646 668898 484688 669134
rect 484368 668866 484688 668898
rect 515088 669454 515408 669486
rect 515088 669218 515130 669454
rect 515366 669218 515408 669454
rect 515088 669134 515408 669218
rect 515088 668898 515130 669134
rect 515366 668898 515408 669134
rect 515088 668866 515408 668898
rect 545808 669454 546128 669486
rect 545808 669218 545850 669454
rect 546086 669218 546128 669454
rect 545808 669134 546128 669218
rect 545808 668898 545850 669134
rect 546086 668898 546128 669134
rect 545808 668866 546128 668898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect 8208 651454 8528 651486
rect 8208 651218 8250 651454
rect 8486 651218 8528 651454
rect 8208 651134 8528 651218
rect 8208 650898 8250 651134
rect 8486 650898 8528 651134
rect 8208 650866 8528 650898
rect 38928 651454 39248 651486
rect 38928 651218 38970 651454
rect 39206 651218 39248 651454
rect 38928 651134 39248 651218
rect 38928 650898 38970 651134
rect 39206 650898 39248 651134
rect 38928 650866 39248 650898
rect 69648 651454 69968 651486
rect 69648 651218 69690 651454
rect 69926 651218 69968 651454
rect 69648 651134 69968 651218
rect 69648 650898 69690 651134
rect 69926 650898 69968 651134
rect 69648 650866 69968 650898
rect 100368 651454 100688 651486
rect 100368 651218 100410 651454
rect 100646 651218 100688 651454
rect 100368 651134 100688 651218
rect 100368 650898 100410 651134
rect 100646 650898 100688 651134
rect 100368 650866 100688 650898
rect 131088 651454 131408 651486
rect 131088 651218 131130 651454
rect 131366 651218 131408 651454
rect 131088 651134 131408 651218
rect 131088 650898 131130 651134
rect 131366 650898 131408 651134
rect 131088 650866 131408 650898
rect 161808 651454 162128 651486
rect 161808 651218 161850 651454
rect 162086 651218 162128 651454
rect 161808 651134 162128 651218
rect 161808 650898 161850 651134
rect 162086 650898 162128 651134
rect 161808 650866 162128 650898
rect 192528 651454 192848 651486
rect 192528 651218 192570 651454
rect 192806 651218 192848 651454
rect 192528 651134 192848 651218
rect 192528 650898 192570 651134
rect 192806 650898 192848 651134
rect 192528 650866 192848 650898
rect 223248 651454 223568 651486
rect 223248 651218 223290 651454
rect 223526 651218 223568 651454
rect 223248 651134 223568 651218
rect 223248 650898 223290 651134
rect 223526 650898 223568 651134
rect 223248 650866 223568 650898
rect 253968 651454 254288 651486
rect 253968 651218 254010 651454
rect 254246 651218 254288 651454
rect 253968 651134 254288 651218
rect 253968 650898 254010 651134
rect 254246 650898 254288 651134
rect 253968 650866 254288 650898
rect 284688 651454 285008 651486
rect 284688 651218 284730 651454
rect 284966 651218 285008 651454
rect 284688 651134 285008 651218
rect 284688 650898 284730 651134
rect 284966 650898 285008 651134
rect 284688 650866 285008 650898
rect 315408 651454 315728 651486
rect 315408 651218 315450 651454
rect 315686 651218 315728 651454
rect 315408 651134 315728 651218
rect 315408 650898 315450 651134
rect 315686 650898 315728 651134
rect 315408 650866 315728 650898
rect 346128 651454 346448 651486
rect 346128 651218 346170 651454
rect 346406 651218 346448 651454
rect 346128 651134 346448 651218
rect 346128 650898 346170 651134
rect 346406 650898 346448 651134
rect 346128 650866 346448 650898
rect 376848 651454 377168 651486
rect 376848 651218 376890 651454
rect 377126 651218 377168 651454
rect 376848 651134 377168 651218
rect 376848 650898 376890 651134
rect 377126 650898 377168 651134
rect 376848 650866 377168 650898
rect 407568 651454 407888 651486
rect 407568 651218 407610 651454
rect 407846 651218 407888 651454
rect 407568 651134 407888 651218
rect 407568 650898 407610 651134
rect 407846 650898 407888 651134
rect 407568 650866 407888 650898
rect 438288 651454 438608 651486
rect 438288 651218 438330 651454
rect 438566 651218 438608 651454
rect 438288 651134 438608 651218
rect 438288 650898 438330 651134
rect 438566 650898 438608 651134
rect 438288 650866 438608 650898
rect 469008 651454 469328 651486
rect 469008 651218 469050 651454
rect 469286 651218 469328 651454
rect 469008 651134 469328 651218
rect 469008 650898 469050 651134
rect 469286 650898 469328 651134
rect 469008 650866 469328 650898
rect 499728 651454 500048 651486
rect 499728 651218 499770 651454
rect 500006 651218 500048 651454
rect 499728 651134 500048 651218
rect 499728 650898 499770 651134
rect 500006 650898 500048 651134
rect 499728 650866 500048 650898
rect 530448 651454 530768 651486
rect 530448 651218 530490 651454
rect 530726 651218 530768 651454
rect 530448 651134 530768 651218
rect 530448 650898 530490 651134
rect 530726 650898 530768 651134
rect 530448 650866 530768 650898
rect 561168 651454 561488 651486
rect 561168 651218 561210 651454
rect 561446 651218 561488 651454
rect 561168 651134 561488 651218
rect 561168 650898 561210 651134
rect 561446 650898 561488 651134
rect 561168 650866 561488 650898
rect 567234 640894 567854 676338
rect 567234 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 567854 640894
rect 567234 640574 567854 640658
rect 567234 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 567854 640574
rect 23568 633454 23888 633486
rect 23568 633218 23610 633454
rect 23846 633218 23888 633454
rect 23568 633134 23888 633218
rect 23568 632898 23610 633134
rect 23846 632898 23888 633134
rect 23568 632866 23888 632898
rect 54288 633454 54608 633486
rect 54288 633218 54330 633454
rect 54566 633218 54608 633454
rect 54288 633134 54608 633218
rect 54288 632898 54330 633134
rect 54566 632898 54608 633134
rect 54288 632866 54608 632898
rect 85008 633454 85328 633486
rect 85008 633218 85050 633454
rect 85286 633218 85328 633454
rect 85008 633134 85328 633218
rect 85008 632898 85050 633134
rect 85286 632898 85328 633134
rect 85008 632866 85328 632898
rect 115728 633454 116048 633486
rect 115728 633218 115770 633454
rect 116006 633218 116048 633454
rect 115728 633134 116048 633218
rect 115728 632898 115770 633134
rect 116006 632898 116048 633134
rect 115728 632866 116048 632898
rect 146448 633454 146768 633486
rect 146448 633218 146490 633454
rect 146726 633218 146768 633454
rect 146448 633134 146768 633218
rect 146448 632898 146490 633134
rect 146726 632898 146768 633134
rect 146448 632866 146768 632898
rect 177168 633454 177488 633486
rect 177168 633218 177210 633454
rect 177446 633218 177488 633454
rect 177168 633134 177488 633218
rect 177168 632898 177210 633134
rect 177446 632898 177488 633134
rect 177168 632866 177488 632898
rect 207888 633454 208208 633486
rect 207888 633218 207930 633454
rect 208166 633218 208208 633454
rect 207888 633134 208208 633218
rect 207888 632898 207930 633134
rect 208166 632898 208208 633134
rect 207888 632866 208208 632898
rect 238608 633454 238928 633486
rect 238608 633218 238650 633454
rect 238886 633218 238928 633454
rect 238608 633134 238928 633218
rect 238608 632898 238650 633134
rect 238886 632898 238928 633134
rect 238608 632866 238928 632898
rect 269328 633454 269648 633486
rect 269328 633218 269370 633454
rect 269606 633218 269648 633454
rect 269328 633134 269648 633218
rect 269328 632898 269370 633134
rect 269606 632898 269648 633134
rect 269328 632866 269648 632898
rect 300048 633454 300368 633486
rect 300048 633218 300090 633454
rect 300326 633218 300368 633454
rect 300048 633134 300368 633218
rect 300048 632898 300090 633134
rect 300326 632898 300368 633134
rect 300048 632866 300368 632898
rect 330768 633454 331088 633486
rect 330768 633218 330810 633454
rect 331046 633218 331088 633454
rect 330768 633134 331088 633218
rect 330768 632898 330810 633134
rect 331046 632898 331088 633134
rect 330768 632866 331088 632898
rect 361488 633454 361808 633486
rect 361488 633218 361530 633454
rect 361766 633218 361808 633454
rect 361488 633134 361808 633218
rect 361488 632898 361530 633134
rect 361766 632898 361808 633134
rect 361488 632866 361808 632898
rect 392208 633454 392528 633486
rect 392208 633218 392250 633454
rect 392486 633218 392528 633454
rect 392208 633134 392528 633218
rect 392208 632898 392250 633134
rect 392486 632898 392528 633134
rect 392208 632866 392528 632898
rect 422928 633454 423248 633486
rect 422928 633218 422970 633454
rect 423206 633218 423248 633454
rect 422928 633134 423248 633218
rect 422928 632898 422970 633134
rect 423206 632898 423248 633134
rect 422928 632866 423248 632898
rect 453648 633454 453968 633486
rect 453648 633218 453690 633454
rect 453926 633218 453968 633454
rect 453648 633134 453968 633218
rect 453648 632898 453690 633134
rect 453926 632898 453968 633134
rect 453648 632866 453968 632898
rect 484368 633454 484688 633486
rect 484368 633218 484410 633454
rect 484646 633218 484688 633454
rect 484368 633134 484688 633218
rect 484368 632898 484410 633134
rect 484646 632898 484688 633134
rect 484368 632866 484688 632898
rect 515088 633454 515408 633486
rect 515088 633218 515130 633454
rect 515366 633218 515408 633454
rect 515088 633134 515408 633218
rect 515088 632898 515130 633134
rect 515366 632898 515408 633134
rect 515088 632866 515408 632898
rect 545808 633454 546128 633486
rect 545808 633218 545850 633454
rect 546086 633218 546128 633454
rect 545808 633134 546128 633218
rect 545808 632898 545850 633134
rect 546086 632898 546128 633134
rect 545808 632866 546128 632898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect 8208 615454 8528 615486
rect 8208 615218 8250 615454
rect 8486 615218 8528 615454
rect 8208 615134 8528 615218
rect 8208 614898 8250 615134
rect 8486 614898 8528 615134
rect 8208 614866 8528 614898
rect 38928 615454 39248 615486
rect 38928 615218 38970 615454
rect 39206 615218 39248 615454
rect 38928 615134 39248 615218
rect 38928 614898 38970 615134
rect 39206 614898 39248 615134
rect 38928 614866 39248 614898
rect 69648 615454 69968 615486
rect 69648 615218 69690 615454
rect 69926 615218 69968 615454
rect 69648 615134 69968 615218
rect 69648 614898 69690 615134
rect 69926 614898 69968 615134
rect 69648 614866 69968 614898
rect 100368 615454 100688 615486
rect 100368 615218 100410 615454
rect 100646 615218 100688 615454
rect 100368 615134 100688 615218
rect 100368 614898 100410 615134
rect 100646 614898 100688 615134
rect 100368 614866 100688 614898
rect 131088 615454 131408 615486
rect 131088 615218 131130 615454
rect 131366 615218 131408 615454
rect 131088 615134 131408 615218
rect 131088 614898 131130 615134
rect 131366 614898 131408 615134
rect 131088 614866 131408 614898
rect 161808 615454 162128 615486
rect 161808 615218 161850 615454
rect 162086 615218 162128 615454
rect 161808 615134 162128 615218
rect 161808 614898 161850 615134
rect 162086 614898 162128 615134
rect 161808 614866 162128 614898
rect 192528 615454 192848 615486
rect 192528 615218 192570 615454
rect 192806 615218 192848 615454
rect 192528 615134 192848 615218
rect 192528 614898 192570 615134
rect 192806 614898 192848 615134
rect 192528 614866 192848 614898
rect 223248 615454 223568 615486
rect 223248 615218 223290 615454
rect 223526 615218 223568 615454
rect 223248 615134 223568 615218
rect 223248 614898 223290 615134
rect 223526 614898 223568 615134
rect 223248 614866 223568 614898
rect 253968 615454 254288 615486
rect 253968 615218 254010 615454
rect 254246 615218 254288 615454
rect 253968 615134 254288 615218
rect 253968 614898 254010 615134
rect 254246 614898 254288 615134
rect 253968 614866 254288 614898
rect 284688 615454 285008 615486
rect 284688 615218 284730 615454
rect 284966 615218 285008 615454
rect 284688 615134 285008 615218
rect 284688 614898 284730 615134
rect 284966 614898 285008 615134
rect 284688 614866 285008 614898
rect 315408 615454 315728 615486
rect 315408 615218 315450 615454
rect 315686 615218 315728 615454
rect 315408 615134 315728 615218
rect 315408 614898 315450 615134
rect 315686 614898 315728 615134
rect 315408 614866 315728 614898
rect 346128 615454 346448 615486
rect 346128 615218 346170 615454
rect 346406 615218 346448 615454
rect 346128 615134 346448 615218
rect 346128 614898 346170 615134
rect 346406 614898 346448 615134
rect 346128 614866 346448 614898
rect 376848 615454 377168 615486
rect 376848 615218 376890 615454
rect 377126 615218 377168 615454
rect 376848 615134 377168 615218
rect 376848 614898 376890 615134
rect 377126 614898 377168 615134
rect 376848 614866 377168 614898
rect 407568 615454 407888 615486
rect 407568 615218 407610 615454
rect 407846 615218 407888 615454
rect 407568 615134 407888 615218
rect 407568 614898 407610 615134
rect 407846 614898 407888 615134
rect 407568 614866 407888 614898
rect 438288 615454 438608 615486
rect 438288 615218 438330 615454
rect 438566 615218 438608 615454
rect 438288 615134 438608 615218
rect 438288 614898 438330 615134
rect 438566 614898 438608 615134
rect 438288 614866 438608 614898
rect 469008 615454 469328 615486
rect 469008 615218 469050 615454
rect 469286 615218 469328 615454
rect 469008 615134 469328 615218
rect 469008 614898 469050 615134
rect 469286 614898 469328 615134
rect 469008 614866 469328 614898
rect 499728 615454 500048 615486
rect 499728 615218 499770 615454
rect 500006 615218 500048 615454
rect 499728 615134 500048 615218
rect 499728 614898 499770 615134
rect 500006 614898 500048 615134
rect 499728 614866 500048 614898
rect 530448 615454 530768 615486
rect 530448 615218 530490 615454
rect 530726 615218 530768 615454
rect 530448 615134 530768 615218
rect 530448 614898 530490 615134
rect 530726 614898 530768 615134
rect 530448 614866 530768 614898
rect 561168 615454 561488 615486
rect 561168 615218 561210 615454
rect 561446 615218 561488 615454
rect 561168 615134 561488 615218
rect 561168 614898 561210 615134
rect 561446 614898 561488 615134
rect 561168 614866 561488 614898
rect 567234 604894 567854 640338
rect 567234 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 567854 604894
rect 567234 604574 567854 604658
rect 567234 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 567854 604574
rect 23568 597454 23888 597486
rect 23568 597218 23610 597454
rect 23846 597218 23888 597454
rect 23568 597134 23888 597218
rect 23568 596898 23610 597134
rect 23846 596898 23888 597134
rect 23568 596866 23888 596898
rect 54288 597454 54608 597486
rect 54288 597218 54330 597454
rect 54566 597218 54608 597454
rect 54288 597134 54608 597218
rect 54288 596898 54330 597134
rect 54566 596898 54608 597134
rect 54288 596866 54608 596898
rect 85008 597454 85328 597486
rect 85008 597218 85050 597454
rect 85286 597218 85328 597454
rect 85008 597134 85328 597218
rect 85008 596898 85050 597134
rect 85286 596898 85328 597134
rect 85008 596866 85328 596898
rect 115728 597454 116048 597486
rect 115728 597218 115770 597454
rect 116006 597218 116048 597454
rect 115728 597134 116048 597218
rect 115728 596898 115770 597134
rect 116006 596898 116048 597134
rect 115728 596866 116048 596898
rect 146448 597454 146768 597486
rect 146448 597218 146490 597454
rect 146726 597218 146768 597454
rect 146448 597134 146768 597218
rect 146448 596898 146490 597134
rect 146726 596898 146768 597134
rect 146448 596866 146768 596898
rect 177168 597454 177488 597486
rect 177168 597218 177210 597454
rect 177446 597218 177488 597454
rect 177168 597134 177488 597218
rect 177168 596898 177210 597134
rect 177446 596898 177488 597134
rect 177168 596866 177488 596898
rect 207888 597454 208208 597486
rect 207888 597218 207930 597454
rect 208166 597218 208208 597454
rect 207888 597134 208208 597218
rect 207888 596898 207930 597134
rect 208166 596898 208208 597134
rect 207888 596866 208208 596898
rect 238608 597454 238928 597486
rect 238608 597218 238650 597454
rect 238886 597218 238928 597454
rect 238608 597134 238928 597218
rect 238608 596898 238650 597134
rect 238886 596898 238928 597134
rect 238608 596866 238928 596898
rect 269328 597454 269648 597486
rect 269328 597218 269370 597454
rect 269606 597218 269648 597454
rect 269328 597134 269648 597218
rect 269328 596898 269370 597134
rect 269606 596898 269648 597134
rect 269328 596866 269648 596898
rect 300048 597454 300368 597486
rect 300048 597218 300090 597454
rect 300326 597218 300368 597454
rect 300048 597134 300368 597218
rect 300048 596898 300090 597134
rect 300326 596898 300368 597134
rect 300048 596866 300368 596898
rect 330768 597454 331088 597486
rect 330768 597218 330810 597454
rect 331046 597218 331088 597454
rect 330768 597134 331088 597218
rect 330768 596898 330810 597134
rect 331046 596898 331088 597134
rect 330768 596866 331088 596898
rect 361488 597454 361808 597486
rect 361488 597218 361530 597454
rect 361766 597218 361808 597454
rect 361488 597134 361808 597218
rect 361488 596898 361530 597134
rect 361766 596898 361808 597134
rect 361488 596866 361808 596898
rect 392208 597454 392528 597486
rect 392208 597218 392250 597454
rect 392486 597218 392528 597454
rect 392208 597134 392528 597218
rect 392208 596898 392250 597134
rect 392486 596898 392528 597134
rect 392208 596866 392528 596898
rect 422928 597454 423248 597486
rect 422928 597218 422970 597454
rect 423206 597218 423248 597454
rect 422928 597134 423248 597218
rect 422928 596898 422970 597134
rect 423206 596898 423248 597134
rect 422928 596866 423248 596898
rect 453648 597454 453968 597486
rect 453648 597218 453690 597454
rect 453926 597218 453968 597454
rect 453648 597134 453968 597218
rect 453648 596898 453690 597134
rect 453926 596898 453968 597134
rect 453648 596866 453968 596898
rect 484368 597454 484688 597486
rect 484368 597218 484410 597454
rect 484646 597218 484688 597454
rect 484368 597134 484688 597218
rect 484368 596898 484410 597134
rect 484646 596898 484688 597134
rect 484368 596866 484688 596898
rect 515088 597454 515408 597486
rect 515088 597218 515130 597454
rect 515366 597218 515408 597454
rect 515088 597134 515408 597218
rect 515088 596898 515130 597134
rect 515366 596898 515408 597134
rect 515088 596866 515408 596898
rect 545808 597454 546128 597486
rect 545808 597218 545850 597454
rect 546086 597218 546128 597454
rect 545808 597134 546128 597218
rect 545808 596898 545850 597134
rect 546086 596898 546128 597134
rect 545808 596866 546128 596898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect 8208 579454 8528 579486
rect 8208 579218 8250 579454
rect 8486 579218 8528 579454
rect 8208 579134 8528 579218
rect 8208 578898 8250 579134
rect 8486 578898 8528 579134
rect 8208 578866 8528 578898
rect 38928 579454 39248 579486
rect 38928 579218 38970 579454
rect 39206 579218 39248 579454
rect 38928 579134 39248 579218
rect 38928 578898 38970 579134
rect 39206 578898 39248 579134
rect 38928 578866 39248 578898
rect 69648 579454 69968 579486
rect 69648 579218 69690 579454
rect 69926 579218 69968 579454
rect 69648 579134 69968 579218
rect 69648 578898 69690 579134
rect 69926 578898 69968 579134
rect 69648 578866 69968 578898
rect 100368 579454 100688 579486
rect 100368 579218 100410 579454
rect 100646 579218 100688 579454
rect 100368 579134 100688 579218
rect 100368 578898 100410 579134
rect 100646 578898 100688 579134
rect 100368 578866 100688 578898
rect 131088 579454 131408 579486
rect 131088 579218 131130 579454
rect 131366 579218 131408 579454
rect 131088 579134 131408 579218
rect 131088 578898 131130 579134
rect 131366 578898 131408 579134
rect 131088 578866 131408 578898
rect 161808 579454 162128 579486
rect 161808 579218 161850 579454
rect 162086 579218 162128 579454
rect 161808 579134 162128 579218
rect 161808 578898 161850 579134
rect 162086 578898 162128 579134
rect 161808 578866 162128 578898
rect 192528 579454 192848 579486
rect 192528 579218 192570 579454
rect 192806 579218 192848 579454
rect 192528 579134 192848 579218
rect 192528 578898 192570 579134
rect 192806 578898 192848 579134
rect 192528 578866 192848 578898
rect 223248 579454 223568 579486
rect 223248 579218 223290 579454
rect 223526 579218 223568 579454
rect 223248 579134 223568 579218
rect 223248 578898 223290 579134
rect 223526 578898 223568 579134
rect 223248 578866 223568 578898
rect 253968 579454 254288 579486
rect 253968 579218 254010 579454
rect 254246 579218 254288 579454
rect 253968 579134 254288 579218
rect 253968 578898 254010 579134
rect 254246 578898 254288 579134
rect 253968 578866 254288 578898
rect 284688 579454 285008 579486
rect 284688 579218 284730 579454
rect 284966 579218 285008 579454
rect 284688 579134 285008 579218
rect 284688 578898 284730 579134
rect 284966 578898 285008 579134
rect 284688 578866 285008 578898
rect 315408 579454 315728 579486
rect 315408 579218 315450 579454
rect 315686 579218 315728 579454
rect 315408 579134 315728 579218
rect 315408 578898 315450 579134
rect 315686 578898 315728 579134
rect 315408 578866 315728 578898
rect 346128 579454 346448 579486
rect 346128 579218 346170 579454
rect 346406 579218 346448 579454
rect 346128 579134 346448 579218
rect 346128 578898 346170 579134
rect 346406 578898 346448 579134
rect 346128 578866 346448 578898
rect 376848 579454 377168 579486
rect 376848 579218 376890 579454
rect 377126 579218 377168 579454
rect 376848 579134 377168 579218
rect 376848 578898 376890 579134
rect 377126 578898 377168 579134
rect 376848 578866 377168 578898
rect 407568 579454 407888 579486
rect 407568 579218 407610 579454
rect 407846 579218 407888 579454
rect 407568 579134 407888 579218
rect 407568 578898 407610 579134
rect 407846 578898 407888 579134
rect 407568 578866 407888 578898
rect 438288 579454 438608 579486
rect 438288 579218 438330 579454
rect 438566 579218 438608 579454
rect 438288 579134 438608 579218
rect 438288 578898 438330 579134
rect 438566 578898 438608 579134
rect 438288 578866 438608 578898
rect 469008 579454 469328 579486
rect 469008 579218 469050 579454
rect 469286 579218 469328 579454
rect 469008 579134 469328 579218
rect 469008 578898 469050 579134
rect 469286 578898 469328 579134
rect 469008 578866 469328 578898
rect 499728 579454 500048 579486
rect 499728 579218 499770 579454
rect 500006 579218 500048 579454
rect 499728 579134 500048 579218
rect 499728 578898 499770 579134
rect 500006 578898 500048 579134
rect 499728 578866 500048 578898
rect 530448 579454 530768 579486
rect 530448 579218 530490 579454
rect 530726 579218 530768 579454
rect 530448 579134 530768 579218
rect 530448 578898 530490 579134
rect 530726 578898 530768 579134
rect 530448 578866 530768 578898
rect 561168 579454 561488 579486
rect 561168 579218 561210 579454
rect 561446 579218 561488 579454
rect 561168 579134 561488 579218
rect 561168 578898 561210 579134
rect 561446 578898 561488 579134
rect 561168 578866 561488 578898
rect 567234 568894 567854 604338
rect 567234 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 567854 568894
rect 567234 568574 567854 568658
rect 567234 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 567854 568574
rect 23568 561454 23888 561486
rect 23568 561218 23610 561454
rect 23846 561218 23888 561454
rect 23568 561134 23888 561218
rect 23568 560898 23610 561134
rect 23846 560898 23888 561134
rect 23568 560866 23888 560898
rect 54288 561454 54608 561486
rect 54288 561218 54330 561454
rect 54566 561218 54608 561454
rect 54288 561134 54608 561218
rect 54288 560898 54330 561134
rect 54566 560898 54608 561134
rect 54288 560866 54608 560898
rect 85008 561454 85328 561486
rect 85008 561218 85050 561454
rect 85286 561218 85328 561454
rect 85008 561134 85328 561218
rect 85008 560898 85050 561134
rect 85286 560898 85328 561134
rect 85008 560866 85328 560898
rect 115728 561454 116048 561486
rect 115728 561218 115770 561454
rect 116006 561218 116048 561454
rect 115728 561134 116048 561218
rect 115728 560898 115770 561134
rect 116006 560898 116048 561134
rect 115728 560866 116048 560898
rect 146448 561454 146768 561486
rect 146448 561218 146490 561454
rect 146726 561218 146768 561454
rect 146448 561134 146768 561218
rect 146448 560898 146490 561134
rect 146726 560898 146768 561134
rect 146448 560866 146768 560898
rect 177168 561454 177488 561486
rect 177168 561218 177210 561454
rect 177446 561218 177488 561454
rect 177168 561134 177488 561218
rect 177168 560898 177210 561134
rect 177446 560898 177488 561134
rect 177168 560866 177488 560898
rect 207888 561454 208208 561486
rect 207888 561218 207930 561454
rect 208166 561218 208208 561454
rect 207888 561134 208208 561218
rect 207888 560898 207930 561134
rect 208166 560898 208208 561134
rect 207888 560866 208208 560898
rect 238608 561454 238928 561486
rect 238608 561218 238650 561454
rect 238886 561218 238928 561454
rect 238608 561134 238928 561218
rect 238608 560898 238650 561134
rect 238886 560898 238928 561134
rect 238608 560866 238928 560898
rect 269328 561454 269648 561486
rect 269328 561218 269370 561454
rect 269606 561218 269648 561454
rect 269328 561134 269648 561218
rect 269328 560898 269370 561134
rect 269606 560898 269648 561134
rect 269328 560866 269648 560898
rect 300048 561454 300368 561486
rect 300048 561218 300090 561454
rect 300326 561218 300368 561454
rect 300048 561134 300368 561218
rect 300048 560898 300090 561134
rect 300326 560898 300368 561134
rect 300048 560866 300368 560898
rect 330768 561454 331088 561486
rect 330768 561218 330810 561454
rect 331046 561218 331088 561454
rect 330768 561134 331088 561218
rect 330768 560898 330810 561134
rect 331046 560898 331088 561134
rect 330768 560866 331088 560898
rect 361488 561454 361808 561486
rect 361488 561218 361530 561454
rect 361766 561218 361808 561454
rect 361488 561134 361808 561218
rect 361488 560898 361530 561134
rect 361766 560898 361808 561134
rect 361488 560866 361808 560898
rect 392208 561454 392528 561486
rect 392208 561218 392250 561454
rect 392486 561218 392528 561454
rect 392208 561134 392528 561218
rect 392208 560898 392250 561134
rect 392486 560898 392528 561134
rect 392208 560866 392528 560898
rect 422928 561454 423248 561486
rect 422928 561218 422970 561454
rect 423206 561218 423248 561454
rect 422928 561134 423248 561218
rect 422928 560898 422970 561134
rect 423206 560898 423248 561134
rect 422928 560866 423248 560898
rect 453648 561454 453968 561486
rect 453648 561218 453690 561454
rect 453926 561218 453968 561454
rect 453648 561134 453968 561218
rect 453648 560898 453690 561134
rect 453926 560898 453968 561134
rect 453648 560866 453968 560898
rect 484368 561454 484688 561486
rect 484368 561218 484410 561454
rect 484646 561218 484688 561454
rect 484368 561134 484688 561218
rect 484368 560898 484410 561134
rect 484646 560898 484688 561134
rect 484368 560866 484688 560898
rect 515088 561454 515408 561486
rect 515088 561218 515130 561454
rect 515366 561218 515408 561454
rect 515088 561134 515408 561218
rect 515088 560898 515130 561134
rect 515366 560898 515408 561134
rect 515088 560866 515408 560898
rect 545808 561454 546128 561486
rect 545808 561218 545850 561454
rect 546086 561218 546128 561454
rect 545808 561134 546128 561218
rect 545808 560898 545850 561134
rect 546086 560898 546128 561134
rect 545808 560866 546128 560898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect 8208 543454 8528 543486
rect 8208 543218 8250 543454
rect 8486 543218 8528 543454
rect 8208 543134 8528 543218
rect 8208 542898 8250 543134
rect 8486 542898 8528 543134
rect 8208 542866 8528 542898
rect 38928 543454 39248 543486
rect 38928 543218 38970 543454
rect 39206 543218 39248 543454
rect 38928 543134 39248 543218
rect 38928 542898 38970 543134
rect 39206 542898 39248 543134
rect 38928 542866 39248 542898
rect 69648 543454 69968 543486
rect 69648 543218 69690 543454
rect 69926 543218 69968 543454
rect 69648 543134 69968 543218
rect 69648 542898 69690 543134
rect 69926 542898 69968 543134
rect 69648 542866 69968 542898
rect 100368 543454 100688 543486
rect 100368 543218 100410 543454
rect 100646 543218 100688 543454
rect 100368 543134 100688 543218
rect 100368 542898 100410 543134
rect 100646 542898 100688 543134
rect 100368 542866 100688 542898
rect 131088 543454 131408 543486
rect 131088 543218 131130 543454
rect 131366 543218 131408 543454
rect 131088 543134 131408 543218
rect 131088 542898 131130 543134
rect 131366 542898 131408 543134
rect 131088 542866 131408 542898
rect 161808 543454 162128 543486
rect 161808 543218 161850 543454
rect 162086 543218 162128 543454
rect 161808 543134 162128 543218
rect 161808 542898 161850 543134
rect 162086 542898 162128 543134
rect 161808 542866 162128 542898
rect 192528 543454 192848 543486
rect 192528 543218 192570 543454
rect 192806 543218 192848 543454
rect 192528 543134 192848 543218
rect 192528 542898 192570 543134
rect 192806 542898 192848 543134
rect 192528 542866 192848 542898
rect 223248 543454 223568 543486
rect 223248 543218 223290 543454
rect 223526 543218 223568 543454
rect 223248 543134 223568 543218
rect 223248 542898 223290 543134
rect 223526 542898 223568 543134
rect 223248 542866 223568 542898
rect 253968 543454 254288 543486
rect 253968 543218 254010 543454
rect 254246 543218 254288 543454
rect 253968 543134 254288 543218
rect 253968 542898 254010 543134
rect 254246 542898 254288 543134
rect 253968 542866 254288 542898
rect 284688 543454 285008 543486
rect 284688 543218 284730 543454
rect 284966 543218 285008 543454
rect 284688 543134 285008 543218
rect 284688 542898 284730 543134
rect 284966 542898 285008 543134
rect 284688 542866 285008 542898
rect 315408 543454 315728 543486
rect 315408 543218 315450 543454
rect 315686 543218 315728 543454
rect 315408 543134 315728 543218
rect 315408 542898 315450 543134
rect 315686 542898 315728 543134
rect 315408 542866 315728 542898
rect 346128 543454 346448 543486
rect 346128 543218 346170 543454
rect 346406 543218 346448 543454
rect 346128 543134 346448 543218
rect 346128 542898 346170 543134
rect 346406 542898 346448 543134
rect 346128 542866 346448 542898
rect 376848 543454 377168 543486
rect 376848 543218 376890 543454
rect 377126 543218 377168 543454
rect 376848 543134 377168 543218
rect 376848 542898 376890 543134
rect 377126 542898 377168 543134
rect 376848 542866 377168 542898
rect 407568 543454 407888 543486
rect 407568 543218 407610 543454
rect 407846 543218 407888 543454
rect 407568 543134 407888 543218
rect 407568 542898 407610 543134
rect 407846 542898 407888 543134
rect 407568 542866 407888 542898
rect 438288 543454 438608 543486
rect 438288 543218 438330 543454
rect 438566 543218 438608 543454
rect 438288 543134 438608 543218
rect 438288 542898 438330 543134
rect 438566 542898 438608 543134
rect 438288 542866 438608 542898
rect 469008 543454 469328 543486
rect 469008 543218 469050 543454
rect 469286 543218 469328 543454
rect 469008 543134 469328 543218
rect 469008 542898 469050 543134
rect 469286 542898 469328 543134
rect 469008 542866 469328 542898
rect 499728 543454 500048 543486
rect 499728 543218 499770 543454
rect 500006 543218 500048 543454
rect 499728 543134 500048 543218
rect 499728 542898 499770 543134
rect 500006 542898 500048 543134
rect 499728 542866 500048 542898
rect 530448 543454 530768 543486
rect 530448 543218 530490 543454
rect 530726 543218 530768 543454
rect 530448 543134 530768 543218
rect 530448 542898 530490 543134
rect 530726 542898 530768 543134
rect 530448 542866 530768 542898
rect 561168 543454 561488 543486
rect 561168 543218 561210 543454
rect 561446 543218 561488 543454
rect 561168 543134 561488 543218
rect 561168 542898 561210 543134
rect 561446 542898 561488 543134
rect 561168 542866 561488 542898
rect 567234 532894 567854 568338
rect 567234 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 567854 532894
rect 567234 532574 567854 532658
rect 567234 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 567854 532574
rect 23568 525454 23888 525486
rect 23568 525218 23610 525454
rect 23846 525218 23888 525454
rect 23568 525134 23888 525218
rect 23568 524898 23610 525134
rect 23846 524898 23888 525134
rect 23568 524866 23888 524898
rect 54288 525454 54608 525486
rect 54288 525218 54330 525454
rect 54566 525218 54608 525454
rect 54288 525134 54608 525218
rect 54288 524898 54330 525134
rect 54566 524898 54608 525134
rect 54288 524866 54608 524898
rect 85008 525454 85328 525486
rect 85008 525218 85050 525454
rect 85286 525218 85328 525454
rect 85008 525134 85328 525218
rect 85008 524898 85050 525134
rect 85286 524898 85328 525134
rect 85008 524866 85328 524898
rect 115728 525454 116048 525486
rect 115728 525218 115770 525454
rect 116006 525218 116048 525454
rect 115728 525134 116048 525218
rect 115728 524898 115770 525134
rect 116006 524898 116048 525134
rect 115728 524866 116048 524898
rect 146448 525454 146768 525486
rect 146448 525218 146490 525454
rect 146726 525218 146768 525454
rect 146448 525134 146768 525218
rect 146448 524898 146490 525134
rect 146726 524898 146768 525134
rect 146448 524866 146768 524898
rect 177168 525454 177488 525486
rect 177168 525218 177210 525454
rect 177446 525218 177488 525454
rect 177168 525134 177488 525218
rect 177168 524898 177210 525134
rect 177446 524898 177488 525134
rect 177168 524866 177488 524898
rect 207888 525454 208208 525486
rect 207888 525218 207930 525454
rect 208166 525218 208208 525454
rect 207888 525134 208208 525218
rect 207888 524898 207930 525134
rect 208166 524898 208208 525134
rect 207888 524866 208208 524898
rect 238608 525454 238928 525486
rect 238608 525218 238650 525454
rect 238886 525218 238928 525454
rect 238608 525134 238928 525218
rect 238608 524898 238650 525134
rect 238886 524898 238928 525134
rect 238608 524866 238928 524898
rect 269328 525454 269648 525486
rect 269328 525218 269370 525454
rect 269606 525218 269648 525454
rect 269328 525134 269648 525218
rect 269328 524898 269370 525134
rect 269606 524898 269648 525134
rect 269328 524866 269648 524898
rect 300048 525454 300368 525486
rect 300048 525218 300090 525454
rect 300326 525218 300368 525454
rect 300048 525134 300368 525218
rect 300048 524898 300090 525134
rect 300326 524898 300368 525134
rect 300048 524866 300368 524898
rect 330768 525454 331088 525486
rect 330768 525218 330810 525454
rect 331046 525218 331088 525454
rect 330768 525134 331088 525218
rect 330768 524898 330810 525134
rect 331046 524898 331088 525134
rect 330768 524866 331088 524898
rect 361488 525454 361808 525486
rect 361488 525218 361530 525454
rect 361766 525218 361808 525454
rect 361488 525134 361808 525218
rect 361488 524898 361530 525134
rect 361766 524898 361808 525134
rect 361488 524866 361808 524898
rect 392208 525454 392528 525486
rect 392208 525218 392250 525454
rect 392486 525218 392528 525454
rect 392208 525134 392528 525218
rect 392208 524898 392250 525134
rect 392486 524898 392528 525134
rect 392208 524866 392528 524898
rect 422928 525454 423248 525486
rect 422928 525218 422970 525454
rect 423206 525218 423248 525454
rect 422928 525134 423248 525218
rect 422928 524898 422970 525134
rect 423206 524898 423248 525134
rect 422928 524866 423248 524898
rect 453648 525454 453968 525486
rect 453648 525218 453690 525454
rect 453926 525218 453968 525454
rect 453648 525134 453968 525218
rect 453648 524898 453690 525134
rect 453926 524898 453968 525134
rect 453648 524866 453968 524898
rect 484368 525454 484688 525486
rect 484368 525218 484410 525454
rect 484646 525218 484688 525454
rect 484368 525134 484688 525218
rect 484368 524898 484410 525134
rect 484646 524898 484688 525134
rect 484368 524866 484688 524898
rect 515088 525454 515408 525486
rect 515088 525218 515130 525454
rect 515366 525218 515408 525454
rect 515088 525134 515408 525218
rect 515088 524898 515130 525134
rect 515366 524898 515408 525134
rect 515088 524866 515408 524898
rect 545808 525454 546128 525486
rect 545808 525218 545850 525454
rect 546086 525218 546128 525454
rect 545808 525134 546128 525218
rect 545808 524898 545850 525134
rect 546086 524898 546128 525134
rect 545808 524866 546128 524898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect 8208 507454 8528 507486
rect 8208 507218 8250 507454
rect 8486 507218 8528 507454
rect 8208 507134 8528 507218
rect 8208 506898 8250 507134
rect 8486 506898 8528 507134
rect 8208 506866 8528 506898
rect 38928 507454 39248 507486
rect 38928 507218 38970 507454
rect 39206 507218 39248 507454
rect 38928 507134 39248 507218
rect 38928 506898 38970 507134
rect 39206 506898 39248 507134
rect 38928 506866 39248 506898
rect 69648 507454 69968 507486
rect 69648 507218 69690 507454
rect 69926 507218 69968 507454
rect 69648 507134 69968 507218
rect 69648 506898 69690 507134
rect 69926 506898 69968 507134
rect 69648 506866 69968 506898
rect 100368 507454 100688 507486
rect 100368 507218 100410 507454
rect 100646 507218 100688 507454
rect 100368 507134 100688 507218
rect 100368 506898 100410 507134
rect 100646 506898 100688 507134
rect 100368 506866 100688 506898
rect 131088 507454 131408 507486
rect 131088 507218 131130 507454
rect 131366 507218 131408 507454
rect 131088 507134 131408 507218
rect 131088 506898 131130 507134
rect 131366 506898 131408 507134
rect 131088 506866 131408 506898
rect 161808 507454 162128 507486
rect 161808 507218 161850 507454
rect 162086 507218 162128 507454
rect 161808 507134 162128 507218
rect 161808 506898 161850 507134
rect 162086 506898 162128 507134
rect 161808 506866 162128 506898
rect 192528 507454 192848 507486
rect 192528 507218 192570 507454
rect 192806 507218 192848 507454
rect 192528 507134 192848 507218
rect 192528 506898 192570 507134
rect 192806 506898 192848 507134
rect 192528 506866 192848 506898
rect 223248 507454 223568 507486
rect 223248 507218 223290 507454
rect 223526 507218 223568 507454
rect 223248 507134 223568 507218
rect 223248 506898 223290 507134
rect 223526 506898 223568 507134
rect 223248 506866 223568 506898
rect 253968 507454 254288 507486
rect 253968 507218 254010 507454
rect 254246 507218 254288 507454
rect 253968 507134 254288 507218
rect 253968 506898 254010 507134
rect 254246 506898 254288 507134
rect 253968 506866 254288 506898
rect 284688 507454 285008 507486
rect 284688 507218 284730 507454
rect 284966 507218 285008 507454
rect 284688 507134 285008 507218
rect 284688 506898 284730 507134
rect 284966 506898 285008 507134
rect 284688 506866 285008 506898
rect 315408 507454 315728 507486
rect 315408 507218 315450 507454
rect 315686 507218 315728 507454
rect 315408 507134 315728 507218
rect 315408 506898 315450 507134
rect 315686 506898 315728 507134
rect 315408 506866 315728 506898
rect 346128 507454 346448 507486
rect 346128 507218 346170 507454
rect 346406 507218 346448 507454
rect 346128 507134 346448 507218
rect 346128 506898 346170 507134
rect 346406 506898 346448 507134
rect 346128 506866 346448 506898
rect 376848 507454 377168 507486
rect 376848 507218 376890 507454
rect 377126 507218 377168 507454
rect 376848 507134 377168 507218
rect 376848 506898 376890 507134
rect 377126 506898 377168 507134
rect 376848 506866 377168 506898
rect 407568 507454 407888 507486
rect 407568 507218 407610 507454
rect 407846 507218 407888 507454
rect 407568 507134 407888 507218
rect 407568 506898 407610 507134
rect 407846 506898 407888 507134
rect 407568 506866 407888 506898
rect 438288 507454 438608 507486
rect 438288 507218 438330 507454
rect 438566 507218 438608 507454
rect 438288 507134 438608 507218
rect 438288 506898 438330 507134
rect 438566 506898 438608 507134
rect 438288 506866 438608 506898
rect 469008 507454 469328 507486
rect 469008 507218 469050 507454
rect 469286 507218 469328 507454
rect 469008 507134 469328 507218
rect 469008 506898 469050 507134
rect 469286 506898 469328 507134
rect 469008 506866 469328 506898
rect 499728 507454 500048 507486
rect 499728 507218 499770 507454
rect 500006 507218 500048 507454
rect 499728 507134 500048 507218
rect 499728 506898 499770 507134
rect 500006 506898 500048 507134
rect 499728 506866 500048 506898
rect 530448 507454 530768 507486
rect 530448 507218 530490 507454
rect 530726 507218 530768 507454
rect 530448 507134 530768 507218
rect 530448 506898 530490 507134
rect 530726 506898 530768 507134
rect 530448 506866 530768 506898
rect 561168 507454 561488 507486
rect 561168 507218 561210 507454
rect 561446 507218 561488 507454
rect 561168 507134 561488 507218
rect 561168 506898 561210 507134
rect 561446 506898 561488 507134
rect 561168 506866 561488 506898
rect 567234 496894 567854 532338
rect 567234 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 567854 496894
rect 567234 496574 567854 496658
rect 567234 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 567854 496574
rect 23568 489454 23888 489486
rect 23568 489218 23610 489454
rect 23846 489218 23888 489454
rect 23568 489134 23888 489218
rect 23568 488898 23610 489134
rect 23846 488898 23888 489134
rect 23568 488866 23888 488898
rect 54288 489454 54608 489486
rect 54288 489218 54330 489454
rect 54566 489218 54608 489454
rect 54288 489134 54608 489218
rect 54288 488898 54330 489134
rect 54566 488898 54608 489134
rect 54288 488866 54608 488898
rect 85008 489454 85328 489486
rect 85008 489218 85050 489454
rect 85286 489218 85328 489454
rect 85008 489134 85328 489218
rect 85008 488898 85050 489134
rect 85286 488898 85328 489134
rect 85008 488866 85328 488898
rect 115728 489454 116048 489486
rect 115728 489218 115770 489454
rect 116006 489218 116048 489454
rect 115728 489134 116048 489218
rect 115728 488898 115770 489134
rect 116006 488898 116048 489134
rect 115728 488866 116048 488898
rect 146448 489454 146768 489486
rect 146448 489218 146490 489454
rect 146726 489218 146768 489454
rect 146448 489134 146768 489218
rect 146448 488898 146490 489134
rect 146726 488898 146768 489134
rect 146448 488866 146768 488898
rect 177168 489454 177488 489486
rect 177168 489218 177210 489454
rect 177446 489218 177488 489454
rect 177168 489134 177488 489218
rect 177168 488898 177210 489134
rect 177446 488898 177488 489134
rect 177168 488866 177488 488898
rect 207888 489454 208208 489486
rect 207888 489218 207930 489454
rect 208166 489218 208208 489454
rect 207888 489134 208208 489218
rect 207888 488898 207930 489134
rect 208166 488898 208208 489134
rect 207888 488866 208208 488898
rect 238608 489454 238928 489486
rect 238608 489218 238650 489454
rect 238886 489218 238928 489454
rect 238608 489134 238928 489218
rect 238608 488898 238650 489134
rect 238886 488898 238928 489134
rect 238608 488866 238928 488898
rect 269328 489454 269648 489486
rect 269328 489218 269370 489454
rect 269606 489218 269648 489454
rect 269328 489134 269648 489218
rect 269328 488898 269370 489134
rect 269606 488898 269648 489134
rect 269328 488866 269648 488898
rect 300048 489454 300368 489486
rect 300048 489218 300090 489454
rect 300326 489218 300368 489454
rect 300048 489134 300368 489218
rect 300048 488898 300090 489134
rect 300326 488898 300368 489134
rect 300048 488866 300368 488898
rect 330768 489454 331088 489486
rect 330768 489218 330810 489454
rect 331046 489218 331088 489454
rect 330768 489134 331088 489218
rect 330768 488898 330810 489134
rect 331046 488898 331088 489134
rect 330768 488866 331088 488898
rect 361488 489454 361808 489486
rect 361488 489218 361530 489454
rect 361766 489218 361808 489454
rect 361488 489134 361808 489218
rect 361488 488898 361530 489134
rect 361766 488898 361808 489134
rect 361488 488866 361808 488898
rect 392208 489454 392528 489486
rect 392208 489218 392250 489454
rect 392486 489218 392528 489454
rect 392208 489134 392528 489218
rect 392208 488898 392250 489134
rect 392486 488898 392528 489134
rect 392208 488866 392528 488898
rect 422928 489454 423248 489486
rect 422928 489218 422970 489454
rect 423206 489218 423248 489454
rect 422928 489134 423248 489218
rect 422928 488898 422970 489134
rect 423206 488898 423248 489134
rect 422928 488866 423248 488898
rect 453648 489454 453968 489486
rect 453648 489218 453690 489454
rect 453926 489218 453968 489454
rect 453648 489134 453968 489218
rect 453648 488898 453690 489134
rect 453926 488898 453968 489134
rect 453648 488866 453968 488898
rect 484368 489454 484688 489486
rect 484368 489218 484410 489454
rect 484646 489218 484688 489454
rect 484368 489134 484688 489218
rect 484368 488898 484410 489134
rect 484646 488898 484688 489134
rect 484368 488866 484688 488898
rect 515088 489454 515408 489486
rect 515088 489218 515130 489454
rect 515366 489218 515408 489454
rect 515088 489134 515408 489218
rect 515088 488898 515130 489134
rect 515366 488898 515408 489134
rect 515088 488866 515408 488898
rect 545808 489454 546128 489486
rect 545808 489218 545850 489454
rect 546086 489218 546128 489454
rect 545808 489134 546128 489218
rect 545808 488898 545850 489134
rect 546086 488898 546128 489134
rect 545808 488866 546128 488898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect 8208 471454 8528 471486
rect 8208 471218 8250 471454
rect 8486 471218 8528 471454
rect 8208 471134 8528 471218
rect 8208 470898 8250 471134
rect 8486 470898 8528 471134
rect 8208 470866 8528 470898
rect 38928 471454 39248 471486
rect 38928 471218 38970 471454
rect 39206 471218 39248 471454
rect 38928 471134 39248 471218
rect 38928 470898 38970 471134
rect 39206 470898 39248 471134
rect 38928 470866 39248 470898
rect 69648 471454 69968 471486
rect 69648 471218 69690 471454
rect 69926 471218 69968 471454
rect 69648 471134 69968 471218
rect 69648 470898 69690 471134
rect 69926 470898 69968 471134
rect 69648 470866 69968 470898
rect 100368 471454 100688 471486
rect 100368 471218 100410 471454
rect 100646 471218 100688 471454
rect 100368 471134 100688 471218
rect 100368 470898 100410 471134
rect 100646 470898 100688 471134
rect 100368 470866 100688 470898
rect 131088 471454 131408 471486
rect 131088 471218 131130 471454
rect 131366 471218 131408 471454
rect 131088 471134 131408 471218
rect 131088 470898 131130 471134
rect 131366 470898 131408 471134
rect 131088 470866 131408 470898
rect 161808 471454 162128 471486
rect 161808 471218 161850 471454
rect 162086 471218 162128 471454
rect 161808 471134 162128 471218
rect 161808 470898 161850 471134
rect 162086 470898 162128 471134
rect 161808 470866 162128 470898
rect 192528 471454 192848 471486
rect 192528 471218 192570 471454
rect 192806 471218 192848 471454
rect 192528 471134 192848 471218
rect 192528 470898 192570 471134
rect 192806 470898 192848 471134
rect 192528 470866 192848 470898
rect 223248 471454 223568 471486
rect 223248 471218 223290 471454
rect 223526 471218 223568 471454
rect 223248 471134 223568 471218
rect 223248 470898 223290 471134
rect 223526 470898 223568 471134
rect 223248 470866 223568 470898
rect 253968 471454 254288 471486
rect 253968 471218 254010 471454
rect 254246 471218 254288 471454
rect 253968 471134 254288 471218
rect 253968 470898 254010 471134
rect 254246 470898 254288 471134
rect 253968 470866 254288 470898
rect 284688 471454 285008 471486
rect 284688 471218 284730 471454
rect 284966 471218 285008 471454
rect 284688 471134 285008 471218
rect 284688 470898 284730 471134
rect 284966 470898 285008 471134
rect 284688 470866 285008 470898
rect 315408 471454 315728 471486
rect 315408 471218 315450 471454
rect 315686 471218 315728 471454
rect 315408 471134 315728 471218
rect 315408 470898 315450 471134
rect 315686 470898 315728 471134
rect 315408 470866 315728 470898
rect 346128 471454 346448 471486
rect 346128 471218 346170 471454
rect 346406 471218 346448 471454
rect 346128 471134 346448 471218
rect 346128 470898 346170 471134
rect 346406 470898 346448 471134
rect 346128 470866 346448 470898
rect 376848 471454 377168 471486
rect 376848 471218 376890 471454
rect 377126 471218 377168 471454
rect 376848 471134 377168 471218
rect 376848 470898 376890 471134
rect 377126 470898 377168 471134
rect 376848 470866 377168 470898
rect 407568 471454 407888 471486
rect 407568 471218 407610 471454
rect 407846 471218 407888 471454
rect 407568 471134 407888 471218
rect 407568 470898 407610 471134
rect 407846 470898 407888 471134
rect 407568 470866 407888 470898
rect 438288 471454 438608 471486
rect 438288 471218 438330 471454
rect 438566 471218 438608 471454
rect 438288 471134 438608 471218
rect 438288 470898 438330 471134
rect 438566 470898 438608 471134
rect 438288 470866 438608 470898
rect 469008 471454 469328 471486
rect 469008 471218 469050 471454
rect 469286 471218 469328 471454
rect 469008 471134 469328 471218
rect 469008 470898 469050 471134
rect 469286 470898 469328 471134
rect 469008 470866 469328 470898
rect 499728 471454 500048 471486
rect 499728 471218 499770 471454
rect 500006 471218 500048 471454
rect 499728 471134 500048 471218
rect 499728 470898 499770 471134
rect 500006 470898 500048 471134
rect 499728 470866 500048 470898
rect 530448 471454 530768 471486
rect 530448 471218 530490 471454
rect 530726 471218 530768 471454
rect 530448 471134 530768 471218
rect 530448 470898 530490 471134
rect 530726 470898 530768 471134
rect 530448 470866 530768 470898
rect 561168 471454 561488 471486
rect 561168 471218 561210 471454
rect 561446 471218 561488 471454
rect 561168 471134 561488 471218
rect 561168 470898 561210 471134
rect 561446 470898 561488 471134
rect 561168 470866 561488 470898
rect 567234 460894 567854 496338
rect 567234 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 567854 460894
rect 567234 460574 567854 460658
rect 567234 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 567854 460574
rect 23568 453454 23888 453486
rect 23568 453218 23610 453454
rect 23846 453218 23888 453454
rect 23568 453134 23888 453218
rect 23568 452898 23610 453134
rect 23846 452898 23888 453134
rect 23568 452866 23888 452898
rect 54288 453454 54608 453486
rect 54288 453218 54330 453454
rect 54566 453218 54608 453454
rect 54288 453134 54608 453218
rect 54288 452898 54330 453134
rect 54566 452898 54608 453134
rect 54288 452866 54608 452898
rect 85008 453454 85328 453486
rect 85008 453218 85050 453454
rect 85286 453218 85328 453454
rect 85008 453134 85328 453218
rect 85008 452898 85050 453134
rect 85286 452898 85328 453134
rect 85008 452866 85328 452898
rect 115728 453454 116048 453486
rect 115728 453218 115770 453454
rect 116006 453218 116048 453454
rect 115728 453134 116048 453218
rect 115728 452898 115770 453134
rect 116006 452898 116048 453134
rect 115728 452866 116048 452898
rect 146448 453454 146768 453486
rect 146448 453218 146490 453454
rect 146726 453218 146768 453454
rect 146448 453134 146768 453218
rect 146448 452898 146490 453134
rect 146726 452898 146768 453134
rect 146448 452866 146768 452898
rect 177168 453454 177488 453486
rect 177168 453218 177210 453454
rect 177446 453218 177488 453454
rect 177168 453134 177488 453218
rect 177168 452898 177210 453134
rect 177446 452898 177488 453134
rect 177168 452866 177488 452898
rect 207888 453454 208208 453486
rect 207888 453218 207930 453454
rect 208166 453218 208208 453454
rect 207888 453134 208208 453218
rect 207888 452898 207930 453134
rect 208166 452898 208208 453134
rect 207888 452866 208208 452898
rect 238608 453454 238928 453486
rect 238608 453218 238650 453454
rect 238886 453218 238928 453454
rect 238608 453134 238928 453218
rect 238608 452898 238650 453134
rect 238886 452898 238928 453134
rect 238608 452866 238928 452898
rect 269328 453454 269648 453486
rect 269328 453218 269370 453454
rect 269606 453218 269648 453454
rect 269328 453134 269648 453218
rect 269328 452898 269370 453134
rect 269606 452898 269648 453134
rect 269328 452866 269648 452898
rect 300048 453454 300368 453486
rect 300048 453218 300090 453454
rect 300326 453218 300368 453454
rect 300048 453134 300368 453218
rect 300048 452898 300090 453134
rect 300326 452898 300368 453134
rect 300048 452866 300368 452898
rect 330768 453454 331088 453486
rect 330768 453218 330810 453454
rect 331046 453218 331088 453454
rect 330768 453134 331088 453218
rect 330768 452898 330810 453134
rect 331046 452898 331088 453134
rect 330768 452866 331088 452898
rect 361488 453454 361808 453486
rect 361488 453218 361530 453454
rect 361766 453218 361808 453454
rect 361488 453134 361808 453218
rect 361488 452898 361530 453134
rect 361766 452898 361808 453134
rect 361488 452866 361808 452898
rect 392208 453454 392528 453486
rect 392208 453218 392250 453454
rect 392486 453218 392528 453454
rect 392208 453134 392528 453218
rect 392208 452898 392250 453134
rect 392486 452898 392528 453134
rect 392208 452866 392528 452898
rect 422928 453454 423248 453486
rect 422928 453218 422970 453454
rect 423206 453218 423248 453454
rect 422928 453134 423248 453218
rect 422928 452898 422970 453134
rect 423206 452898 423248 453134
rect 422928 452866 423248 452898
rect 453648 453454 453968 453486
rect 453648 453218 453690 453454
rect 453926 453218 453968 453454
rect 453648 453134 453968 453218
rect 453648 452898 453690 453134
rect 453926 452898 453968 453134
rect 453648 452866 453968 452898
rect 484368 453454 484688 453486
rect 484368 453218 484410 453454
rect 484646 453218 484688 453454
rect 484368 453134 484688 453218
rect 484368 452898 484410 453134
rect 484646 452898 484688 453134
rect 484368 452866 484688 452898
rect 515088 453454 515408 453486
rect 515088 453218 515130 453454
rect 515366 453218 515408 453454
rect 515088 453134 515408 453218
rect 515088 452898 515130 453134
rect 515366 452898 515408 453134
rect 515088 452866 515408 452898
rect 545808 453454 546128 453486
rect 545808 453218 545850 453454
rect 546086 453218 546128 453454
rect 545808 453134 546128 453218
rect 545808 452898 545850 453134
rect 546086 452898 546128 453134
rect 545808 452866 546128 452898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect 8208 435454 8528 435486
rect 8208 435218 8250 435454
rect 8486 435218 8528 435454
rect 8208 435134 8528 435218
rect 8208 434898 8250 435134
rect 8486 434898 8528 435134
rect 8208 434866 8528 434898
rect 38928 435454 39248 435486
rect 38928 435218 38970 435454
rect 39206 435218 39248 435454
rect 38928 435134 39248 435218
rect 38928 434898 38970 435134
rect 39206 434898 39248 435134
rect 38928 434866 39248 434898
rect 69648 435454 69968 435486
rect 69648 435218 69690 435454
rect 69926 435218 69968 435454
rect 69648 435134 69968 435218
rect 69648 434898 69690 435134
rect 69926 434898 69968 435134
rect 69648 434866 69968 434898
rect 100368 435454 100688 435486
rect 100368 435218 100410 435454
rect 100646 435218 100688 435454
rect 100368 435134 100688 435218
rect 100368 434898 100410 435134
rect 100646 434898 100688 435134
rect 100368 434866 100688 434898
rect 131088 435454 131408 435486
rect 131088 435218 131130 435454
rect 131366 435218 131408 435454
rect 131088 435134 131408 435218
rect 131088 434898 131130 435134
rect 131366 434898 131408 435134
rect 131088 434866 131408 434898
rect 161808 435454 162128 435486
rect 161808 435218 161850 435454
rect 162086 435218 162128 435454
rect 161808 435134 162128 435218
rect 161808 434898 161850 435134
rect 162086 434898 162128 435134
rect 161808 434866 162128 434898
rect 192528 435454 192848 435486
rect 192528 435218 192570 435454
rect 192806 435218 192848 435454
rect 192528 435134 192848 435218
rect 192528 434898 192570 435134
rect 192806 434898 192848 435134
rect 192528 434866 192848 434898
rect 223248 435454 223568 435486
rect 223248 435218 223290 435454
rect 223526 435218 223568 435454
rect 223248 435134 223568 435218
rect 223248 434898 223290 435134
rect 223526 434898 223568 435134
rect 223248 434866 223568 434898
rect 253968 435454 254288 435486
rect 253968 435218 254010 435454
rect 254246 435218 254288 435454
rect 253968 435134 254288 435218
rect 253968 434898 254010 435134
rect 254246 434898 254288 435134
rect 253968 434866 254288 434898
rect 284688 435454 285008 435486
rect 284688 435218 284730 435454
rect 284966 435218 285008 435454
rect 284688 435134 285008 435218
rect 284688 434898 284730 435134
rect 284966 434898 285008 435134
rect 284688 434866 285008 434898
rect 315408 435454 315728 435486
rect 315408 435218 315450 435454
rect 315686 435218 315728 435454
rect 315408 435134 315728 435218
rect 315408 434898 315450 435134
rect 315686 434898 315728 435134
rect 315408 434866 315728 434898
rect 346128 435454 346448 435486
rect 346128 435218 346170 435454
rect 346406 435218 346448 435454
rect 346128 435134 346448 435218
rect 346128 434898 346170 435134
rect 346406 434898 346448 435134
rect 346128 434866 346448 434898
rect 376848 435454 377168 435486
rect 376848 435218 376890 435454
rect 377126 435218 377168 435454
rect 376848 435134 377168 435218
rect 376848 434898 376890 435134
rect 377126 434898 377168 435134
rect 376848 434866 377168 434898
rect 407568 435454 407888 435486
rect 407568 435218 407610 435454
rect 407846 435218 407888 435454
rect 407568 435134 407888 435218
rect 407568 434898 407610 435134
rect 407846 434898 407888 435134
rect 407568 434866 407888 434898
rect 438288 435454 438608 435486
rect 438288 435218 438330 435454
rect 438566 435218 438608 435454
rect 438288 435134 438608 435218
rect 438288 434898 438330 435134
rect 438566 434898 438608 435134
rect 438288 434866 438608 434898
rect 469008 435454 469328 435486
rect 469008 435218 469050 435454
rect 469286 435218 469328 435454
rect 469008 435134 469328 435218
rect 469008 434898 469050 435134
rect 469286 434898 469328 435134
rect 469008 434866 469328 434898
rect 499728 435454 500048 435486
rect 499728 435218 499770 435454
rect 500006 435218 500048 435454
rect 499728 435134 500048 435218
rect 499728 434898 499770 435134
rect 500006 434898 500048 435134
rect 499728 434866 500048 434898
rect 530448 435454 530768 435486
rect 530448 435218 530490 435454
rect 530726 435218 530768 435454
rect 530448 435134 530768 435218
rect 530448 434898 530490 435134
rect 530726 434898 530768 435134
rect 530448 434866 530768 434898
rect 561168 435454 561488 435486
rect 561168 435218 561210 435454
rect 561446 435218 561488 435454
rect 561168 435134 561488 435218
rect 561168 434898 561210 435134
rect 561446 434898 561488 435134
rect 561168 434866 561488 434898
rect 567234 424894 567854 460338
rect 567234 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 567854 424894
rect 567234 424574 567854 424658
rect 567234 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 567854 424574
rect 23568 417454 23888 417486
rect 23568 417218 23610 417454
rect 23846 417218 23888 417454
rect 23568 417134 23888 417218
rect 23568 416898 23610 417134
rect 23846 416898 23888 417134
rect 23568 416866 23888 416898
rect 54288 417454 54608 417486
rect 54288 417218 54330 417454
rect 54566 417218 54608 417454
rect 54288 417134 54608 417218
rect 54288 416898 54330 417134
rect 54566 416898 54608 417134
rect 54288 416866 54608 416898
rect 85008 417454 85328 417486
rect 85008 417218 85050 417454
rect 85286 417218 85328 417454
rect 85008 417134 85328 417218
rect 85008 416898 85050 417134
rect 85286 416898 85328 417134
rect 85008 416866 85328 416898
rect 115728 417454 116048 417486
rect 115728 417218 115770 417454
rect 116006 417218 116048 417454
rect 115728 417134 116048 417218
rect 115728 416898 115770 417134
rect 116006 416898 116048 417134
rect 115728 416866 116048 416898
rect 146448 417454 146768 417486
rect 146448 417218 146490 417454
rect 146726 417218 146768 417454
rect 146448 417134 146768 417218
rect 146448 416898 146490 417134
rect 146726 416898 146768 417134
rect 146448 416866 146768 416898
rect 177168 417454 177488 417486
rect 177168 417218 177210 417454
rect 177446 417218 177488 417454
rect 177168 417134 177488 417218
rect 177168 416898 177210 417134
rect 177446 416898 177488 417134
rect 177168 416866 177488 416898
rect 207888 417454 208208 417486
rect 207888 417218 207930 417454
rect 208166 417218 208208 417454
rect 207888 417134 208208 417218
rect 207888 416898 207930 417134
rect 208166 416898 208208 417134
rect 207888 416866 208208 416898
rect 238608 417454 238928 417486
rect 238608 417218 238650 417454
rect 238886 417218 238928 417454
rect 238608 417134 238928 417218
rect 238608 416898 238650 417134
rect 238886 416898 238928 417134
rect 238608 416866 238928 416898
rect 269328 417454 269648 417486
rect 269328 417218 269370 417454
rect 269606 417218 269648 417454
rect 269328 417134 269648 417218
rect 269328 416898 269370 417134
rect 269606 416898 269648 417134
rect 269328 416866 269648 416898
rect 300048 417454 300368 417486
rect 300048 417218 300090 417454
rect 300326 417218 300368 417454
rect 300048 417134 300368 417218
rect 300048 416898 300090 417134
rect 300326 416898 300368 417134
rect 300048 416866 300368 416898
rect 330768 417454 331088 417486
rect 330768 417218 330810 417454
rect 331046 417218 331088 417454
rect 330768 417134 331088 417218
rect 330768 416898 330810 417134
rect 331046 416898 331088 417134
rect 330768 416866 331088 416898
rect 361488 417454 361808 417486
rect 361488 417218 361530 417454
rect 361766 417218 361808 417454
rect 361488 417134 361808 417218
rect 361488 416898 361530 417134
rect 361766 416898 361808 417134
rect 361488 416866 361808 416898
rect 392208 417454 392528 417486
rect 392208 417218 392250 417454
rect 392486 417218 392528 417454
rect 392208 417134 392528 417218
rect 392208 416898 392250 417134
rect 392486 416898 392528 417134
rect 392208 416866 392528 416898
rect 422928 417454 423248 417486
rect 422928 417218 422970 417454
rect 423206 417218 423248 417454
rect 422928 417134 423248 417218
rect 422928 416898 422970 417134
rect 423206 416898 423248 417134
rect 422928 416866 423248 416898
rect 453648 417454 453968 417486
rect 453648 417218 453690 417454
rect 453926 417218 453968 417454
rect 453648 417134 453968 417218
rect 453648 416898 453690 417134
rect 453926 416898 453968 417134
rect 453648 416866 453968 416898
rect 484368 417454 484688 417486
rect 484368 417218 484410 417454
rect 484646 417218 484688 417454
rect 484368 417134 484688 417218
rect 484368 416898 484410 417134
rect 484646 416898 484688 417134
rect 484368 416866 484688 416898
rect 515088 417454 515408 417486
rect 515088 417218 515130 417454
rect 515366 417218 515408 417454
rect 515088 417134 515408 417218
rect 515088 416898 515130 417134
rect 515366 416898 515408 417134
rect 515088 416866 515408 416898
rect 545808 417454 546128 417486
rect 545808 417218 545850 417454
rect 546086 417218 546128 417454
rect 545808 417134 546128 417218
rect 545808 416898 545850 417134
rect 546086 416898 546128 417134
rect 545808 416866 546128 416898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect 8208 399454 8528 399486
rect 8208 399218 8250 399454
rect 8486 399218 8528 399454
rect 8208 399134 8528 399218
rect 8208 398898 8250 399134
rect 8486 398898 8528 399134
rect 8208 398866 8528 398898
rect 38928 399454 39248 399486
rect 38928 399218 38970 399454
rect 39206 399218 39248 399454
rect 38928 399134 39248 399218
rect 38928 398898 38970 399134
rect 39206 398898 39248 399134
rect 38928 398866 39248 398898
rect 69648 399454 69968 399486
rect 69648 399218 69690 399454
rect 69926 399218 69968 399454
rect 69648 399134 69968 399218
rect 69648 398898 69690 399134
rect 69926 398898 69968 399134
rect 69648 398866 69968 398898
rect 100368 399454 100688 399486
rect 100368 399218 100410 399454
rect 100646 399218 100688 399454
rect 100368 399134 100688 399218
rect 100368 398898 100410 399134
rect 100646 398898 100688 399134
rect 100368 398866 100688 398898
rect 131088 399454 131408 399486
rect 131088 399218 131130 399454
rect 131366 399218 131408 399454
rect 131088 399134 131408 399218
rect 131088 398898 131130 399134
rect 131366 398898 131408 399134
rect 131088 398866 131408 398898
rect 161808 399454 162128 399486
rect 161808 399218 161850 399454
rect 162086 399218 162128 399454
rect 161808 399134 162128 399218
rect 161808 398898 161850 399134
rect 162086 398898 162128 399134
rect 161808 398866 162128 398898
rect 192528 399454 192848 399486
rect 192528 399218 192570 399454
rect 192806 399218 192848 399454
rect 192528 399134 192848 399218
rect 192528 398898 192570 399134
rect 192806 398898 192848 399134
rect 192528 398866 192848 398898
rect 223248 399454 223568 399486
rect 223248 399218 223290 399454
rect 223526 399218 223568 399454
rect 223248 399134 223568 399218
rect 223248 398898 223290 399134
rect 223526 398898 223568 399134
rect 223248 398866 223568 398898
rect 253968 399454 254288 399486
rect 253968 399218 254010 399454
rect 254246 399218 254288 399454
rect 253968 399134 254288 399218
rect 253968 398898 254010 399134
rect 254246 398898 254288 399134
rect 253968 398866 254288 398898
rect 284688 399454 285008 399486
rect 284688 399218 284730 399454
rect 284966 399218 285008 399454
rect 284688 399134 285008 399218
rect 284688 398898 284730 399134
rect 284966 398898 285008 399134
rect 284688 398866 285008 398898
rect 315408 399454 315728 399486
rect 315408 399218 315450 399454
rect 315686 399218 315728 399454
rect 315408 399134 315728 399218
rect 315408 398898 315450 399134
rect 315686 398898 315728 399134
rect 315408 398866 315728 398898
rect 346128 399454 346448 399486
rect 346128 399218 346170 399454
rect 346406 399218 346448 399454
rect 346128 399134 346448 399218
rect 346128 398898 346170 399134
rect 346406 398898 346448 399134
rect 346128 398866 346448 398898
rect 376848 399454 377168 399486
rect 376848 399218 376890 399454
rect 377126 399218 377168 399454
rect 376848 399134 377168 399218
rect 376848 398898 376890 399134
rect 377126 398898 377168 399134
rect 376848 398866 377168 398898
rect 407568 399454 407888 399486
rect 407568 399218 407610 399454
rect 407846 399218 407888 399454
rect 407568 399134 407888 399218
rect 407568 398898 407610 399134
rect 407846 398898 407888 399134
rect 407568 398866 407888 398898
rect 438288 399454 438608 399486
rect 438288 399218 438330 399454
rect 438566 399218 438608 399454
rect 438288 399134 438608 399218
rect 438288 398898 438330 399134
rect 438566 398898 438608 399134
rect 438288 398866 438608 398898
rect 469008 399454 469328 399486
rect 469008 399218 469050 399454
rect 469286 399218 469328 399454
rect 469008 399134 469328 399218
rect 469008 398898 469050 399134
rect 469286 398898 469328 399134
rect 469008 398866 469328 398898
rect 499728 399454 500048 399486
rect 499728 399218 499770 399454
rect 500006 399218 500048 399454
rect 499728 399134 500048 399218
rect 499728 398898 499770 399134
rect 500006 398898 500048 399134
rect 499728 398866 500048 398898
rect 530448 399454 530768 399486
rect 530448 399218 530490 399454
rect 530726 399218 530768 399454
rect 530448 399134 530768 399218
rect 530448 398898 530490 399134
rect 530726 398898 530768 399134
rect 530448 398866 530768 398898
rect 561168 399454 561488 399486
rect 561168 399218 561210 399454
rect 561446 399218 561488 399454
rect 561168 399134 561488 399218
rect 561168 398898 561210 399134
rect 561446 398898 561488 399134
rect 561168 398866 561488 398898
rect 567234 388894 567854 424338
rect 567234 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 567854 388894
rect 567234 388574 567854 388658
rect 567234 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 567854 388574
rect 23568 381454 23888 381486
rect 23568 381218 23610 381454
rect 23846 381218 23888 381454
rect 23568 381134 23888 381218
rect 23568 380898 23610 381134
rect 23846 380898 23888 381134
rect 23568 380866 23888 380898
rect 54288 381454 54608 381486
rect 54288 381218 54330 381454
rect 54566 381218 54608 381454
rect 54288 381134 54608 381218
rect 54288 380898 54330 381134
rect 54566 380898 54608 381134
rect 54288 380866 54608 380898
rect 85008 381454 85328 381486
rect 85008 381218 85050 381454
rect 85286 381218 85328 381454
rect 85008 381134 85328 381218
rect 85008 380898 85050 381134
rect 85286 380898 85328 381134
rect 85008 380866 85328 380898
rect 115728 381454 116048 381486
rect 115728 381218 115770 381454
rect 116006 381218 116048 381454
rect 115728 381134 116048 381218
rect 115728 380898 115770 381134
rect 116006 380898 116048 381134
rect 115728 380866 116048 380898
rect 146448 381454 146768 381486
rect 146448 381218 146490 381454
rect 146726 381218 146768 381454
rect 146448 381134 146768 381218
rect 146448 380898 146490 381134
rect 146726 380898 146768 381134
rect 146448 380866 146768 380898
rect 177168 381454 177488 381486
rect 177168 381218 177210 381454
rect 177446 381218 177488 381454
rect 177168 381134 177488 381218
rect 177168 380898 177210 381134
rect 177446 380898 177488 381134
rect 177168 380866 177488 380898
rect 207888 381454 208208 381486
rect 207888 381218 207930 381454
rect 208166 381218 208208 381454
rect 207888 381134 208208 381218
rect 207888 380898 207930 381134
rect 208166 380898 208208 381134
rect 207888 380866 208208 380898
rect 238608 381454 238928 381486
rect 238608 381218 238650 381454
rect 238886 381218 238928 381454
rect 238608 381134 238928 381218
rect 238608 380898 238650 381134
rect 238886 380898 238928 381134
rect 238608 380866 238928 380898
rect 269328 381454 269648 381486
rect 269328 381218 269370 381454
rect 269606 381218 269648 381454
rect 269328 381134 269648 381218
rect 269328 380898 269370 381134
rect 269606 380898 269648 381134
rect 269328 380866 269648 380898
rect 300048 381454 300368 381486
rect 300048 381218 300090 381454
rect 300326 381218 300368 381454
rect 300048 381134 300368 381218
rect 300048 380898 300090 381134
rect 300326 380898 300368 381134
rect 300048 380866 300368 380898
rect 330768 381454 331088 381486
rect 330768 381218 330810 381454
rect 331046 381218 331088 381454
rect 330768 381134 331088 381218
rect 330768 380898 330810 381134
rect 331046 380898 331088 381134
rect 330768 380866 331088 380898
rect 361488 381454 361808 381486
rect 361488 381218 361530 381454
rect 361766 381218 361808 381454
rect 361488 381134 361808 381218
rect 361488 380898 361530 381134
rect 361766 380898 361808 381134
rect 361488 380866 361808 380898
rect 392208 381454 392528 381486
rect 392208 381218 392250 381454
rect 392486 381218 392528 381454
rect 392208 381134 392528 381218
rect 392208 380898 392250 381134
rect 392486 380898 392528 381134
rect 392208 380866 392528 380898
rect 422928 381454 423248 381486
rect 422928 381218 422970 381454
rect 423206 381218 423248 381454
rect 422928 381134 423248 381218
rect 422928 380898 422970 381134
rect 423206 380898 423248 381134
rect 422928 380866 423248 380898
rect 453648 381454 453968 381486
rect 453648 381218 453690 381454
rect 453926 381218 453968 381454
rect 453648 381134 453968 381218
rect 453648 380898 453690 381134
rect 453926 380898 453968 381134
rect 453648 380866 453968 380898
rect 484368 381454 484688 381486
rect 484368 381218 484410 381454
rect 484646 381218 484688 381454
rect 484368 381134 484688 381218
rect 484368 380898 484410 381134
rect 484646 380898 484688 381134
rect 484368 380866 484688 380898
rect 515088 381454 515408 381486
rect 515088 381218 515130 381454
rect 515366 381218 515408 381454
rect 515088 381134 515408 381218
rect 515088 380898 515130 381134
rect 515366 380898 515408 381134
rect 515088 380866 515408 380898
rect 545808 381454 546128 381486
rect 545808 381218 545850 381454
rect 546086 381218 546128 381454
rect 545808 381134 546128 381218
rect 545808 380898 545850 381134
rect 546086 380898 546128 381134
rect 545808 380866 546128 380898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect 8208 363454 8528 363486
rect 8208 363218 8250 363454
rect 8486 363218 8528 363454
rect 8208 363134 8528 363218
rect 8208 362898 8250 363134
rect 8486 362898 8528 363134
rect 8208 362866 8528 362898
rect 38928 363454 39248 363486
rect 38928 363218 38970 363454
rect 39206 363218 39248 363454
rect 38928 363134 39248 363218
rect 38928 362898 38970 363134
rect 39206 362898 39248 363134
rect 38928 362866 39248 362898
rect 69648 363454 69968 363486
rect 69648 363218 69690 363454
rect 69926 363218 69968 363454
rect 69648 363134 69968 363218
rect 69648 362898 69690 363134
rect 69926 362898 69968 363134
rect 69648 362866 69968 362898
rect 100368 363454 100688 363486
rect 100368 363218 100410 363454
rect 100646 363218 100688 363454
rect 100368 363134 100688 363218
rect 100368 362898 100410 363134
rect 100646 362898 100688 363134
rect 100368 362866 100688 362898
rect 131088 363454 131408 363486
rect 131088 363218 131130 363454
rect 131366 363218 131408 363454
rect 131088 363134 131408 363218
rect 131088 362898 131130 363134
rect 131366 362898 131408 363134
rect 131088 362866 131408 362898
rect 161808 363454 162128 363486
rect 161808 363218 161850 363454
rect 162086 363218 162128 363454
rect 161808 363134 162128 363218
rect 161808 362898 161850 363134
rect 162086 362898 162128 363134
rect 161808 362866 162128 362898
rect 192528 363454 192848 363486
rect 192528 363218 192570 363454
rect 192806 363218 192848 363454
rect 192528 363134 192848 363218
rect 192528 362898 192570 363134
rect 192806 362898 192848 363134
rect 192528 362866 192848 362898
rect 223248 363454 223568 363486
rect 223248 363218 223290 363454
rect 223526 363218 223568 363454
rect 223248 363134 223568 363218
rect 223248 362898 223290 363134
rect 223526 362898 223568 363134
rect 223248 362866 223568 362898
rect 253968 363454 254288 363486
rect 253968 363218 254010 363454
rect 254246 363218 254288 363454
rect 253968 363134 254288 363218
rect 253968 362898 254010 363134
rect 254246 362898 254288 363134
rect 253968 362866 254288 362898
rect 284688 363454 285008 363486
rect 284688 363218 284730 363454
rect 284966 363218 285008 363454
rect 284688 363134 285008 363218
rect 284688 362898 284730 363134
rect 284966 362898 285008 363134
rect 284688 362866 285008 362898
rect 315408 363454 315728 363486
rect 315408 363218 315450 363454
rect 315686 363218 315728 363454
rect 315408 363134 315728 363218
rect 315408 362898 315450 363134
rect 315686 362898 315728 363134
rect 315408 362866 315728 362898
rect 346128 363454 346448 363486
rect 346128 363218 346170 363454
rect 346406 363218 346448 363454
rect 346128 363134 346448 363218
rect 346128 362898 346170 363134
rect 346406 362898 346448 363134
rect 346128 362866 346448 362898
rect 376848 363454 377168 363486
rect 376848 363218 376890 363454
rect 377126 363218 377168 363454
rect 376848 363134 377168 363218
rect 376848 362898 376890 363134
rect 377126 362898 377168 363134
rect 376848 362866 377168 362898
rect 407568 363454 407888 363486
rect 407568 363218 407610 363454
rect 407846 363218 407888 363454
rect 407568 363134 407888 363218
rect 407568 362898 407610 363134
rect 407846 362898 407888 363134
rect 407568 362866 407888 362898
rect 438288 363454 438608 363486
rect 438288 363218 438330 363454
rect 438566 363218 438608 363454
rect 438288 363134 438608 363218
rect 438288 362898 438330 363134
rect 438566 362898 438608 363134
rect 438288 362866 438608 362898
rect 469008 363454 469328 363486
rect 469008 363218 469050 363454
rect 469286 363218 469328 363454
rect 469008 363134 469328 363218
rect 469008 362898 469050 363134
rect 469286 362898 469328 363134
rect 469008 362866 469328 362898
rect 499728 363454 500048 363486
rect 499728 363218 499770 363454
rect 500006 363218 500048 363454
rect 499728 363134 500048 363218
rect 499728 362898 499770 363134
rect 500006 362898 500048 363134
rect 499728 362866 500048 362898
rect 530448 363454 530768 363486
rect 530448 363218 530490 363454
rect 530726 363218 530768 363454
rect 530448 363134 530768 363218
rect 530448 362898 530490 363134
rect 530726 362898 530768 363134
rect 530448 362866 530768 362898
rect 561168 363454 561488 363486
rect 561168 363218 561210 363454
rect 561446 363218 561488 363454
rect 561168 363134 561488 363218
rect 561168 362898 561210 363134
rect 561446 362898 561488 363134
rect 561168 362866 561488 362898
rect 567234 352894 567854 388338
rect 567234 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 567854 352894
rect 567234 352574 567854 352658
rect 567234 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 567854 352574
rect 23568 345454 23888 345486
rect 23568 345218 23610 345454
rect 23846 345218 23888 345454
rect 23568 345134 23888 345218
rect 23568 344898 23610 345134
rect 23846 344898 23888 345134
rect 23568 344866 23888 344898
rect 54288 345454 54608 345486
rect 54288 345218 54330 345454
rect 54566 345218 54608 345454
rect 54288 345134 54608 345218
rect 54288 344898 54330 345134
rect 54566 344898 54608 345134
rect 54288 344866 54608 344898
rect 85008 345454 85328 345486
rect 85008 345218 85050 345454
rect 85286 345218 85328 345454
rect 85008 345134 85328 345218
rect 85008 344898 85050 345134
rect 85286 344898 85328 345134
rect 85008 344866 85328 344898
rect 115728 345454 116048 345486
rect 115728 345218 115770 345454
rect 116006 345218 116048 345454
rect 115728 345134 116048 345218
rect 115728 344898 115770 345134
rect 116006 344898 116048 345134
rect 115728 344866 116048 344898
rect 146448 345454 146768 345486
rect 146448 345218 146490 345454
rect 146726 345218 146768 345454
rect 146448 345134 146768 345218
rect 146448 344898 146490 345134
rect 146726 344898 146768 345134
rect 146448 344866 146768 344898
rect 177168 345454 177488 345486
rect 177168 345218 177210 345454
rect 177446 345218 177488 345454
rect 177168 345134 177488 345218
rect 177168 344898 177210 345134
rect 177446 344898 177488 345134
rect 177168 344866 177488 344898
rect 207888 345454 208208 345486
rect 207888 345218 207930 345454
rect 208166 345218 208208 345454
rect 207888 345134 208208 345218
rect 207888 344898 207930 345134
rect 208166 344898 208208 345134
rect 207888 344866 208208 344898
rect 238608 345454 238928 345486
rect 238608 345218 238650 345454
rect 238886 345218 238928 345454
rect 238608 345134 238928 345218
rect 238608 344898 238650 345134
rect 238886 344898 238928 345134
rect 238608 344866 238928 344898
rect 269328 345454 269648 345486
rect 269328 345218 269370 345454
rect 269606 345218 269648 345454
rect 269328 345134 269648 345218
rect 269328 344898 269370 345134
rect 269606 344898 269648 345134
rect 269328 344866 269648 344898
rect 300048 345454 300368 345486
rect 300048 345218 300090 345454
rect 300326 345218 300368 345454
rect 300048 345134 300368 345218
rect 300048 344898 300090 345134
rect 300326 344898 300368 345134
rect 300048 344866 300368 344898
rect 330768 345454 331088 345486
rect 330768 345218 330810 345454
rect 331046 345218 331088 345454
rect 330768 345134 331088 345218
rect 330768 344898 330810 345134
rect 331046 344898 331088 345134
rect 330768 344866 331088 344898
rect 361488 345454 361808 345486
rect 361488 345218 361530 345454
rect 361766 345218 361808 345454
rect 361488 345134 361808 345218
rect 361488 344898 361530 345134
rect 361766 344898 361808 345134
rect 361488 344866 361808 344898
rect 392208 345454 392528 345486
rect 392208 345218 392250 345454
rect 392486 345218 392528 345454
rect 392208 345134 392528 345218
rect 392208 344898 392250 345134
rect 392486 344898 392528 345134
rect 392208 344866 392528 344898
rect 422928 345454 423248 345486
rect 422928 345218 422970 345454
rect 423206 345218 423248 345454
rect 422928 345134 423248 345218
rect 422928 344898 422970 345134
rect 423206 344898 423248 345134
rect 422928 344866 423248 344898
rect 453648 345454 453968 345486
rect 453648 345218 453690 345454
rect 453926 345218 453968 345454
rect 453648 345134 453968 345218
rect 453648 344898 453690 345134
rect 453926 344898 453968 345134
rect 453648 344866 453968 344898
rect 484368 345454 484688 345486
rect 484368 345218 484410 345454
rect 484646 345218 484688 345454
rect 484368 345134 484688 345218
rect 484368 344898 484410 345134
rect 484646 344898 484688 345134
rect 484368 344866 484688 344898
rect 515088 345454 515408 345486
rect 515088 345218 515130 345454
rect 515366 345218 515408 345454
rect 515088 345134 515408 345218
rect 515088 344898 515130 345134
rect 515366 344898 515408 345134
rect 515088 344866 515408 344898
rect 545808 345454 546128 345486
rect 545808 345218 545850 345454
rect 546086 345218 546128 345454
rect 545808 345134 546128 345218
rect 545808 344898 545850 345134
rect 546086 344898 546128 345134
rect 545808 344866 546128 344898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect 8208 327454 8528 327486
rect 8208 327218 8250 327454
rect 8486 327218 8528 327454
rect 8208 327134 8528 327218
rect 8208 326898 8250 327134
rect 8486 326898 8528 327134
rect 8208 326866 8528 326898
rect 38928 327454 39248 327486
rect 38928 327218 38970 327454
rect 39206 327218 39248 327454
rect 38928 327134 39248 327218
rect 38928 326898 38970 327134
rect 39206 326898 39248 327134
rect 38928 326866 39248 326898
rect 69648 327454 69968 327486
rect 69648 327218 69690 327454
rect 69926 327218 69968 327454
rect 69648 327134 69968 327218
rect 69648 326898 69690 327134
rect 69926 326898 69968 327134
rect 69648 326866 69968 326898
rect 100368 327454 100688 327486
rect 100368 327218 100410 327454
rect 100646 327218 100688 327454
rect 100368 327134 100688 327218
rect 100368 326898 100410 327134
rect 100646 326898 100688 327134
rect 100368 326866 100688 326898
rect 131088 327454 131408 327486
rect 131088 327218 131130 327454
rect 131366 327218 131408 327454
rect 131088 327134 131408 327218
rect 131088 326898 131130 327134
rect 131366 326898 131408 327134
rect 131088 326866 131408 326898
rect 161808 327454 162128 327486
rect 161808 327218 161850 327454
rect 162086 327218 162128 327454
rect 161808 327134 162128 327218
rect 161808 326898 161850 327134
rect 162086 326898 162128 327134
rect 161808 326866 162128 326898
rect 192528 327454 192848 327486
rect 192528 327218 192570 327454
rect 192806 327218 192848 327454
rect 192528 327134 192848 327218
rect 192528 326898 192570 327134
rect 192806 326898 192848 327134
rect 192528 326866 192848 326898
rect 223248 327454 223568 327486
rect 223248 327218 223290 327454
rect 223526 327218 223568 327454
rect 223248 327134 223568 327218
rect 223248 326898 223290 327134
rect 223526 326898 223568 327134
rect 223248 326866 223568 326898
rect 253968 327454 254288 327486
rect 253968 327218 254010 327454
rect 254246 327218 254288 327454
rect 253968 327134 254288 327218
rect 253968 326898 254010 327134
rect 254246 326898 254288 327134
rect 253968 326866 254288 326898
rect 284688 327454 285008 327486
rect 284688 327218 284730 327454
rect 284966 327218 285008 327454
rect 284688 327134 285008 327218
rect 284688 326898 284730 327134
rect 284966 326898 285008 327134
rect 284688 326866 285008 326898
rect 315408 327454 315728 327486
rect 315408 327218 315450 327454
rect 315686 327218 315728 327454
rect 315408 327134 315728 327218
rect 315408 326898 315450 327134
rect 315686 326898 315728 327134
rect 315408 326866 315728 326898
rect 346128 327454 346448 327486
rect 346128 327218 346170 327454
rect 346406 327218 346448 327454
rect 346128 327134 346448 327218
rect 346128 326898 346170 327134
rect 346406 326898 346448 327134
rect 346128 326866 346448 326898
rect 376848 327454 377168 327486
rect 376848 327218 376890 327454
rect 377126 327218 377168 327454
rect 376848 327134 377168 327218
rect 376848 326898 376890 327134
rect 377126 326898 377168 327134
rect 376848 326866 377168 326898
rect 407568 327454 407888 327486
rect 407568 327218 407610 327454
rect 407846 327218 407888 327454
rect 407568 327134 407888 327218
rect 407568 326898 407610 327134
rect 407846 326898 407888 327134
rect 407568 326866 407888 326898
rect 438288 327454 438608 327486
rect 438288 327218 438330 327454
rect 438566 327218 438608 327454
rect 438288 327134 438608 327218
rect 438288 326898 438330 327134
rect 438566 326898 438608 327134
rect 438288 326866 438608 326898
rect 469008 327454 469328 327486
rect 469008 327218 469050 327454
rect 469286 327218 469328 327454
rect 469008 327134 469328 327218
rect 469008 326898 469050 327134
rect 469286 326898 469328 327134
rect 469008 326866 469328 326898
rect 499728 327454 500048 327486
rect 499728 327218 499770 327454
rect 500006 327218 500048 327454
rect 499728 327134 500048 327218
rect 499728 326898 499770 327134
rect 500006 326898 500048 327134
rect 499728 326866 500048 326898
rect 530448 327454 530768 327486
rect 530448 327218 530490 327454
rect 530726 327218 530768 327454
rect 530448 327134 530768 327218
rect 530448 326898 530490 327134
rect 530726 326898 530768 327134
rect 530448 326866 530768 326898
rect 561168 327454 561488 327486
rect 561168 327218 561210 327454
rect 561446 327218 561488 327454
rect 561168 327134 561488 327218
rect 561168 326898 561210 327134
rect 561446 326898 561488 327134
rect 561168 326866 561488 326898
rect 567234 316894 567854 352338
rect 567234 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 567854 316894
rect 567234 316574 567854 316658
rect 567234 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 567854 316574
rect 23568 309454 23888 309486
rect 23568 309218 23610 309454
rect 23846 309218 23888 309454
rect 23568 309134 23888 309218
rect 23568 308898 23610 309134
rect 23846 308898 23888 309134
rect 23568 308866 23888 308898
rect 54288 309454 54608 309486
rect 54288 309218 54330 309454
rect 54566 309218 54608 309454
rect 54288 309134 54608 309218
rect 54288 308898 54330 309134
rect 54566 308898 54608 309134
rect 54288 308866 54608 308898
rect 85008 309454 85328 309486
rect 85008 309218 85050 309454
rect 85286 309218 85328 309454
rect 85008 309134 85328 309218
rect 85008 308898 85050 309134
rect 85286 308898 85328 309134
rect 85008 308866 85328 308898
rect 115728 309454 116048 309486
rect 115728 309218 115770 309454
rect 116006 309218 116048 309454
rect 115728 309134 116048 309218
rect 115728 308898 115770 309134
rect 116006 308898 116048 309134
rect 115728 308866 116048 308898
rect 146448 309454 146768 309486
rect 146448 309218 146490 309454
rect 146726 309218 146768 309454
rect 146448 309134 146768 309218
rect 146448 308898 146490 309134
rect 146726 308898 146768 309134
rect 146448 308866 146768 308898
rect 177168 309454 177488 309486
rect 177168 309218 177210 309454
rect 177446 309218 177488 309454
rect 177168 309134 177488 309218
rect 177168 308898 177210 309134
rect 177446 308898 177488 309134
rect 177168 308866 177488 308898
rect 207888 309454 208208 309486
rect 207888 309218 207930 309454
rect 208166 309218 208208 309454
rect 207888 309134 208208 309218
rect 207888 308898 207930 309134
rect 208166 308898 208208 309134
rect 207888 308866 208208 308898
rect 238608 309454 238928 309486
rect 238608 309218 238650 309454
rect 238886 309218 238928 309454
rect 238608 309134 238928 309218
rect 238608 308898 238650 309134
rect 238886 308898 238928 309134
rect 238608 308866 238928 308898
rect 269328 309454 269648 309486
rect 269328 309218 269370 309454
rect 269606 309218 269648 309454
rect 269328 309134 269648 309218
rect 269328 308898 269370 309134
rect 269606 308898 269648 309134
rect 269328 308866 269648 308898
rect 300048 309454 300368 309486
rect 300048 309218 300090 309454
rect 300326 309218 300368 309454
rect 300048 309134 300368 309218
rect 300048 308898 300090 309134
rect 300326 308898 300368 309134
rect 300048 308866 300368 308898
rect 330768 309454 331088 309486
rect 330768 309218 330810 309454
rect 331046 309218 331088 309454
rect 330768 309134 331088 309218
rect 330768 308898 330810 309134
rect 331046 308898 331088 309134
rect 330768 308866 331088 308898
rect 361488 309454 361808 309486
rect 361488 309218 361530 309454
rect 361766 309218 361808 309454
rect 361488 309134 361808 309218
rect 361488 308898 361530 309134
rect 361766 308898 361808 309134
rect 361488 308866 361808 308898
rect 392208 309454 392528 309486
rect 392208 309218 392250 309454
rect 392486 309218 392528 309454
rect 392208 309134 392528 309218
rect 392208 308898 392250 309134
rect 392486 308898 392528 309134
rect 392208 308866 392528 308898
rect 422928 309454 423248 309486
rect 422928 309218 422970 309454
rect 423206 309218 423248 309454
rect 422928 309134 423248 309218
rect 422928 308898 422970 309134
rect 423206 308898 423248 309134
rect 422928 308866 423248 308898
rect 453648 309454 453968 309486
rect 453648 309218 453690 309454
rect 453926 309218 453968 309454
rect 453648 309134 453968 309218
rect 453648 308898 453690 309134
rect 453926 308898 453968 309134
rect 453648 308866 453968 308898
rect 484368 309454 484688 309486
rect 484368 309218 484410 309454
rect 484646 309218 484688 309454
rect 484368 309134 484688 309218
rect 484368 308898 484410 309134
rect 484646 308898 484688 309134
rect 484368 308866 484688 308898
rect 515088 309454 515408 309486
rect 515088 309218 515130 309454
rect 515366 309218 515408 309454
rect 515088 309134 515408 309218
rect 515088 308898 515130 309134
rect 515366 308898 515408 309134
rect 515088 308866 515408 308898
rect 545808 309454 546128 309486
rect 545808 309218 545850 309454
rect 546086 309218 546128 309454
rect 545808 309134 546128 309218
rect 545808 308898 545850 309134
rect 546086 308898 546128 309134
rect 545808 308866 546128 308898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect 8208 291454 8528 291486
rect 8208 291218 8250 291454
rect 8486 291218 8528 291454
rect 8208 291134 8528 291218
rect 8208 290898 8250 291134
rect 8486 290898 8528 291134
rect 8208 290866 8528 290898
rect 38928 291454 39248 291486
rect 38928 291218 38970 291454
rect 39206 291218 39248 291454
rect 38928 291134 39248 291218
rect 38928 290898 38970 291134
rect 39206 290898 39248 291134
rect 38928 290866 39248 290898
rect 69648 291454 69968 291486
rect 69648 291218 69690 291454
rect 69926 291218 69968 291454
rect 69648 291134 69968 291218
rect 69648 290898 69690 291134
rect 69926 290898 69968 291134
rect 69648 290866 69968 290898
rect 100368 291454 100688 291486
rect 100368 291218 100410 291454
rect 100646 291218 100688 291454
rect 100368 291134 100688 291218
rect 100368 290898 100410 291134
rect 100646 290898 100688 291134
rect 100368 290866 100688 290898
rect 131088 291454 131408 291486
rect 131088 291218 131130 291454
rect 131366 291218 131408 291454
rect 131088 291134 131408 291218
rect 131088 290898 131130 291134
rect 131366 290898 131408 291134
rect 131088 290866 131408 290898
rect 161808 291454 162128 291486
rect 161808 291218 161850 291454
rect 162086 291218 162128 291454
rect 161808 291134 162128 291218
rect 161808 290898 161850 291134
rect 162086 290898 162128 291134
rect 161808 290866 162128 290898
rect 192528 291454 192848 291486
rect 192528 291218 192570 291454
rect 192806 291218 192848 291454
rect 192528 291134 192848 291218
rect 192528 290898 192570 291134
rect 192806 290898 192848 291134
rect 192528 290866 192848 290898
rect 223248 291454 223568 291486
rect 223248 291218 223290 291454
rect 223526 291218 223568 291454
rect 223248 291134 223568 291218
rect 223248 290898 223290 291134
rect 223526 290898 223568 291134
rect 223248 290866 223568 290898
rect 253968 291454 254288 291486
rect 253968 291218 254010 291454
rect 254246 291218 254288 291454
rect 253968 291134 254288 291218
rect 253968 290898 254010 291134
rect 254246 290898 254288 291134
rect 253968 290866 254288 290898
rect 284688 291454 285008 291486
rect 284688 291218 284730 291454
rect 284966 291218 285008 291454
rect 284688 291134 285008 291218
rect 284688 290898 284730 291134
rect 284966 290898 285008 291134
rect 284688 290866 285008 290898
rect 315408 291454 315728 291486
rect 315408 291218 315450 291454
rect 315686 291218 315728 291454
rect 315408 291134 315728 291218
rect 315408 290898 315450 291134
rect 315686 290898 315728 291134
rect 315408 290866 315728 290898
rect 346128 291454 346448 291486
rect 346128 291218 346170 291454
rect 346406 291218 346448 291454
rect 346128 291134 346448 291218
rect 346128 290898 346170 291134
rect 346406 290898 346448 291134
rect 346128 290866 346448 290898
rect 376848 291454 377168 291486
rect 376848 291218 376890 291454
rect 377126 291218 377168 291454
rect 376848 291134 377168 291218
rect 376848 290898 376890 291134
rect 377126 290898 377168 291134
rect 376848 290866 377168 290898
rect 407568 291454 407888 291486
rect 407568 291218 407610 291454
rect 407846 291218 407888 291454
rect 407568 291134 407888 291218
rect 407568 290898 407610 291134
rect 407846 290898 407888 291134
rect 407568 290866 407888 290898
rect 438288 291454 438608 291486
rect 438288 291218 438330 291454
rect 438566 291218 438608 291454
rect 438288 291134 438608 291218
rect 438288 290898 438330 291134
rect 438566 290898 438608 291134
rect 438288 290866 438608 290898
rect 469008 291454 469328 291486
rect 469008 291218 469050 291454
rect 469286 291218 469328 291454
rect 469008 291134 469328 291218
rect 469008 290898 469050 291134
rect 469286 290898 469328 291134
rect 469008 290866 469328 290898
rect 499728 291454 500048 291486
rect 499728 291218 499770 291454
rect 500006 291218 500048 291454
rect 499728 291134 500048 291218
rect 499728 290898 499770 291134
rect 500006 290898 500048 291134
rect 499728 290866 500048 290898
rect 530448 291454 530768 291486
rect 530448 291218 530490 291454
rect 530726 291218 530768 291454
rect 530448 291134 530768 291218
rect 530448 290898 530490 291134
rect 530726 290898 530768 291134
rect 530448 290866 530768 290898
rect 561168 291454 561488 291486
rect 561168 291218 561210 291454
rect 561446 291218 561488 291454
rect 561168 291134 561488 291218
rect 561168 290898 561210 291134
rect 561446 290898 561488 291134
rect 561168 290866 561488 290898
rect 567234 280894 567854 316338
rect 567234 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 567854 280894
rect 567234 280574 567854 280658
rect 567234 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 567854 280574
rect 23568 273454 23888 273486
rect 23568 273218 23610 273454
rect 23846 273218 23888 273454
rect 23568 273134 23888 273218
rect 23568 272898 23610 273134
rect 23846 272898 23888 273134
rect 23568 272866 23888 272898
rect 54288 273454 54608 273486
rect 54288 273218 54330 273454
rect 54566 273218 54608 273454
rect 54288 273134 54608 273218
rect 54288 272898 54330 273134
rect 54566 272898 54608 273134
rect 54288 272866 54608 272898
rect 85008 273454 85328 273486
rect 85008 273218 85050 273454
rect 85286 273218 85328 273454
rect 85008 273134 85328 273218
rect 85008 272898 85050 273134
rect 85286 272898 85328 273134
rect 85008 272866 85328 272898
rect 115728 273454 116048 273486
rect 115728 273218 115770 273454
rect 116006 273218 116048 273454
rect 115728 273134 116048 273218
rect 115728 272898 115770 273134
rect 116006 272898 116048 273134
rect 115728 272866 116048 272898
rect 146448 273454 146768 273486
rect 146448 273218 146490 273454
rect 146726 273218 146768 273454
rect 146448 273134 146768 273218
rect 146448 272898 146490 273134
rect 146726 272898 146768 273134
rect 146448 272866 146768 272898
rect 177168 273454 177488 273486
rect 177168 273218 177210 273454
rect 177446 273218 177488 273454
rect 177168 273134 177488 273218
rect 177168 272898 177210 273134
rect 177446 272898 177488 273134
rect 177168 272866 177488 272898
rect 207888 273454 208208 273486
rect 207888 273218 207930 273454
rect 208166 273218 208208 273454
rect 207888 273134 208208 273218
rect 207888 272898 207930 273134
rect 208166 272898 208208 273134
rect 207888 272866 208208 272898
rect 238608 273454 238928 273486
rect 238608 273218 238650 273454
rect 238886 273218 238928 273454
rect 238608 273134 238928 273218
rect 238608 272898 238650 273134
rect 238886 272898 238928 273134
rect 238608 272866 238928 272898
rect 269328 273454 269648 273486
rect 269328 273218 269370 273454
rect 269606 273218 269648 273454
rect 269328 273134 269648 273218
rect 269328 272898 269370 273134
rect 269606 272898 269648 273134
rect 269328 272866 269648 272898
rect 300048 273454 300368 273486
rect 300048 273218 300090 273454
rect 300326 273218 300368 273454
rect 300048 273134 300368 273218
rect 300048 272898 300090 273134
rect 300326 272898 300368 273134
rect 300048 272866 300368 272898
rect 330768 273454 331088 273486
rect 330768 273218 330810 273454
rect 331046 273218 331088 273454
rect 330768 273134 331088 273218
rect 330768 272898 330810 273134
rect 331046 272898 331088 273134
rect 330768 272866 331088 272898
rect 361488 273454 361808 273486
rect 361488 273218 361530 273454
rect 361766 273218 361808 273454
rect 361488 273134 361808 273218
rect 361488 272898 361530 273134
rect 361766 272898 361808 273134
rect 361488 272866 361808 272898
rect 392208 273454 392528 273486
rect 392208 273218 392250 273454
rect 392486 273218 392528 273454
rect 392208 273134 392528 273218
rect 392208 272898 392250 273134
rect 392486 272898 392528 273134
rect 392208 272866 392528 272898
rect 422928 273454 423248 273486
rect 422928 273218 422970 273454
rect 423206 273218 423248 273454
rect 422928 273134 423248 273218
rect 422928 272898 422970 273134
rect 423206 272898 423248 273134
rect 422928 272866 423248 272898
rect 453648 273454 453968 273486
rect 453648 273218 453690 273454
rect 453926 273218 453968 273454
rect 453648 273134 453968 273218
rect 453648 272898 453690 273134
rect 453926 272898 453968 273134
rect 453648 272866 453968 272898
rect 484368 273454 484688 273486
rect 484368 273218 484410 273454
rect 484646 273218 484688 273454
rect 484368 273134 484688 273218
rect 484368 272898 484410 273134
rect 484646 272898 484688 273134
rect 484368 272866 484688 272898
rect 515088 273454 515408 273486
rect 515088 273218 515130 273454
rect 515366 273218 515408 273454
rect 515088 273134 515408 273218
rect 515088 272898 515130 273134
rect 515366 272898 515408 273134
rect 515088 272866 515408 272898
rect 545808 273454 546128 273486
rect 545808 273218 545850 273454
rect 546086 273218 546128 273454
rect 545808 273134 546128 273218
rect 545808 272898 545850 273134
rect 546086 272898 546128 273134
rect 545808 272866 546128 272898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect 8208 255454 8528 255486
rect 8208 255218 8250 255454
rect 8486 255218 8528 255454
rect 8208 255134 8528 255218
rect 8208 254898 8250 255134
rect 8486 254898 8528 255134
rect 8208 254866 8528 254898
rect 38928 255454 39248 255486
rect 38928 255218 38970 255454
rect 39206 255218 39248 255454
rect 38928 255134 39248 255218
rect 38928 254898 38970 255134
rect 39206 254898 39248 255134
rect 38928 254866 39248 254898
rect 69648 255454 69968 255486
rect 69648 255218 69690 255454
rect 69926 255218 69968 255454
rect 69648 255134 69968 255218
rect 69648 254898 69690 255134
rect 69926 254898 69968 255134
rect 69648 254866 69968 254898
rect 100368 255454 100688 255486
rect 100368 255218 100410 255454
rect 100646 255218 100688 255454
rect 100368 255134 100688 255218
rect 100368 254898 100410 255134
rect 100646 254898 100688 255134
rect 100368 254866 100688 254898
rect 131088 255454 131408 255486
rect 131088 255218 131130 255454
rect 131366 255218 131408 255454
rect 131088 255134 131408 255218
rect 131088 254898 131130 255134
rect 131366 254898 131408 255134
rect 131088 254866 131408 254898
rect 161808 255454 162128 255486
rect 161808 255218 161850 255454
rect 162086 255218 162128 255454
rect 161808 255134 162128 255218
rect 161808 254898 161850 255134
rect 162086 254898 162128 255134
rect 161808 254866 162128 254898
rect 192528 255454 192848 255486
rect 192528 255218 192570 255454
rect 192806 255218 192848 255454
rect 192528 255134 192848 255218
rect 192528 254898 192570 255134
rect 192806 254898 192848 255134
rect 192528 254866 192848 254898
rect 223248 255454 223568 255486
rect 223248 255218 223290 255454
rect 223526 255218 223568 255454
rect 223248 255134 223568 255218
rect 223248 254898 223290 255134
rect 223526 254898 223568 255134
rect 223248 254866 223568 254898
rect 253968 255454 254288 255486
rect 253968 255218 254010 255454
rect 254246 255218 254288 255454
rect 253968 255134 254288 255218
rect 253968 254898 254010 255134
rect 254246 254898 254288 255134
rect 253968 254866 254288 254898
rect 284688 255454 285008 255486
rect 284688 255218 284730 255454
rect 284966 255218 285008 255454
rect 284688 255134 285008 255218
rect 284688 254898 284730 255134
rect 284966 254898 285008 255134
rect 284688 254866 285008 254898
rect 315408 255454 315728 255486
rect 315408 255218 315450 255454
rect 315686 255218 315728 255454
rect 315408 255134 315728 255218
rect 315408 254898 315450 255134
rect 315686 254898 315728 255134
rect 315408 254866 315728 254898
rect 346128 255454 346448 255486
rect 346128 255218 346170 255454
rect 346406 255218 346448 255454
rect 346128 255134 346448 255218
rect 346128 254898 346170 255134
rect 346406 254898 346448 255134
rect 346128 254866 346448 254898
rect 376848 255454 377168 255486
rect 376848 255218 376890 255454
rect 377126 255218 377168 255454
rect 376848 255134 377168 255218
rect 376848 254898 376890 255134
rect 377126 254898 377168 255134
rect 376848 254866 377168 254898
rect 407568 255454 407888 255486
rect 407568 255218 407610 255454
rect 407846 255218 407888 255454
rect 407568 255134 407888 255218
rect 407568 254898 407610 255134
rect 407846 254898 407888 255134
rect 407568 254866 407888 254898
rect 438288 255454 438608 255486
rect 438288 255218 438330 255454
rect 438566 255218 438608 255454
rect 438288 255134 438608 255218
rect 438288 254898 438330 255134
rect 438566 254898 438608 255134
rect 438288 254866 438608 254898
rect 469008 255454 469328 255486
rect 469008 255218 469050 255454
rect 469286 255218 469328 255454
rect 469008 255134 469328 255218
rect 469008 254898 469050 255134
rect 469286 254898 469328 255134
rect 469008 254866 469328 254898
rect 499728 255454 500048 255486
rect 499728 255218 499770 255454
rect 500006 255218 500048 255454
rect 499728 255134 500048 255218
rect 499728 254898 499770 255134
rect 500006 254898 500048 255134
rect 499728 254866 500048 254898
rect 530448 255454 530768 255486
rect 530448 255218 530490 255454
rect 530726 255218 530768 255454
rect 530448 255134 530768 255218
rect 530448 254898 530490 255134
rect 530726 254898 530768 255134
rect 530448 254866 530768 254898
rect 561168 255454 561488 255486
rect 561168 255218 561210 255454
rect 561446 255218 561488 255454
rect 561168 255134 561488 255218
rect 561168 254898 561210 255134
rect 561446 254898 561488 255134
rect 561168 254866 561488 254898
rect 567234 244894 567854 280338
rect 567234 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 567854 244894
rect 567234 244574 567854 244658
rect 567234 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 567854 244574
rect 23568 237454 23888 237486
rect 23568 237218 23610 237454
rect 23846 237218 23888 237454
rect 23568 237134 23888 237218
rect 23568 236898 23610 237134
rect 23846 236898 23888 237134
rect 23568 236866 23888 236898
rect 54288 237454 54608 237486
rect 54288 237218 54330 237454
rect 54566 237218 54608 237454
rect 54288 237134 54608 237218
rect 54288 236898 54330 237134
rect 54566 236898 54608 237134
rect 54288 236866 54608 236898
rect 85008 237454 85328 237486
rect 85008 237218 85050 237454
rect 85286 237218 85328 237454
rect 85008 237134 85328 237218
rect 85008 236898 85050 237134
rect 85286 236898 85328 237134
rect 85008 236866 85328 236898
rect 115728 237454 116048 237486
rect 115728 237218 115770 237454
rect 116006 237218 116048 237454
rect 115728 237134 116048 237218
rect 115728 236898 115770 237134
rect 116006 236898 116048 237134
rect 115728 236866 116048 236898
rect 146448 237454 146768 237486
rect 146448 237218 146490 237454
rect 146726 237218 146768 237454
rect 146448 237134 146768 237218
rect 146448 236898 146490 237134
rect 146726 236898 146768 237134
rect 146448 236866 146768 236898
rect 177168 237454 177488 237486
rect 177168 237218 177210 237454
rect 177446 237218 177488 237454
rect 177168 237134 177488 237218
rect 177168 236898 177210 237134
rect 177446 236898 177488 237134
rect 177168 236866 177488 236898
rect 207888 237454 208208 237486
rect 207888 237218 207930 237454
rect 208166 237218 208208 237454
rect 207888 237134 208208 237218
rect 207888 236898 207930 237134
rect 208166 236898 208208 237134
rect 207888 236866 208208 236898
rect 238608 237454 238928 237486
rect 238608 237218 238650 237454
rect 238886 237218 238928 237454
rect 238608 237134 238928 237218
rect 238608 236898 238650 237134
rect 238886 236898 238928 237134
rect 238608 236866 238928 236898
rect 269328 237454 269648 237486
rect 269328 237218 269370 237454
rect 269606 237218 269648 237454
rect 269328 237134 269648 237218
rect 269328 236898 269370 237134
rect 269606 236898 269648 237134
rect 269328 236866 269648 236898
rect 300048 237454 300368 237486
rect 300048 237218 300090 237454
rect 300326 237218 300368 237454
rect 300048 237134 300368 237218
rect 300048 236898 300090 237134
rect 300326 236898 300368 237134
rect 300048 236866 300368 236898
rect 330768 237454 331088 237486
rect 330768 237218 330810 237454
rect 331046 237218 331088 237454
rect 330768 237134 331088 237218
rect 330768 236898 330810 237134
rect 331046 236898 331088 237134
rect 330768 236866 331088 236898
rect 361488 237454 361808 237486
rect 361488 237218 361530 237454
rect 361766 237218 361808 237454
rect 361488 237134 361808 237218
rect 361488 236898 361530 237134
rect 361766 236898 361808 237134
rect 361488 236866 361808 236898
rect 392208 237454 392528 237486
rect 392208 237218 392250 237454
rect 392486 237218 392528 237454
rect 392208 237134 392528 237218
rect 392208 236898 392250 237134
rect 392486 236898 392528 237134
rect 392208 236866 392528 236898
rect 422928 237454 423248 237486
rect 422928 237218 422970 237454
rect 423206 237218 423248 237454
rect 422928 237134 423248 237218
rect 422928 236898 422970 237134
rect 423206 236898 423248 237134
rect 422928 236866 423248 236898
rect 453648 237454 453968 237486
rect 453648 237218 453690 237454
rect 453926 237218 453968 237454
rect 453648 237134 453968 237218
rect 453648 236898 453690 237134
rect 453926 236898 453968 237134
rect 453648 236866 453968 236898
rect 484368 237454 484688 237486
rect 484368 237218 484410 237454
rect 484646 237218 484688 237454
rect 484368 237134 484688 237218
rect 484368 236898 484410 237134
rect 484646 236898 484688 237134
rect 484368 236866 484688 236898
rect 515088 237454 515408 237486
rect 515088 237218 515130 237454
rect 515366 237218 515408 237454
rect 515088 237134 515408 237218
rect 515088 236898 515130 237134
rect 515366 236898 515408 237134
rect 515088 236866 515408 236898
rect 545808 237454 546128 237486
rect 545808 237218 545850 237454
rect 546086 237218 546128 237454
rect 545808 237134 546128 237218
rect 545808 236898 545850 237134
rect 546086 236898 546128 237134
rect 545808 236866 546128 236898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect 8208 219454 8528 219486
rect 8208 219218 8250 219454
rect 8486 219218 8528 219454
rect 8208 219134 8528 219218
rect 8208 218898 8250 219134
rect 8486 218898 8528 219134
rect 8208 218866 8528 218898
rect 38928 219454 39248 219486
rect 38928 219218 38970 219454
rect 39206 219218 39248 219454
rect 38928 219134 39248 219218
rect 38928 218898 38970 219134
rect 39206 218898 39248 219134
rect 38928 218866 39248 218898
rect 69648 219454 69968 219486
rect 69648 219218 69690 219454
rect 69926 219218 69968 219454
rect 69648 219134 69968 219218
rect 69648 218898 69690 219134
rect 69926 218898 69968 219134
rect 69648 218866 69968 218898
rect 100368 219454 100688 219486
rect 100368 219218 100410 219454
rect 100646 219218 100688 219454
rect 100368 219134 100688 219218
rect 100368 218898 100410 219134
rect 100646 218898 100688 219134
rect 100368 218866 100688 218898
rect 131088 219454 131408 219486
rect 131088 219218 131130 219454
rect 131366 219218 131408 219454
rect 131088 219134 131408 219218
rect 131088 218898 131130 219134
rect 131366 218898 131408 219134
rect 131088 218866 131408 218898
rect 161808 219454 162128 219486
rect 161808 219218 161850 219454
rect 162086 219218 162128 219454
rect 161808 219134 162128 219218
rect 161808 218898 161850 219134
rect 162086 218898 162128 219134
rect 161808 218866 162128 218898
rect 192528 219454 192848 219486
rect 192528 219218 192570 219454
rect 192806 219218 192848 219454
rect 192528 219134 192848 219218
rect 192528 218898 192570 219134
rect 192806 218898 192848 219134
rect 192528 218866 192848 218898
rect 223248 219454 223568 219486
rect 223248 219218 223290 219454
rect 223526 219218 223568 219454
rect 223248 219134 223568 219218
rect 223248 218898 223290 219134
rect 223526 218898 223568 219134
rect 223248 218866 223568 218898
rect 253968 219454 254288 219486
rect 253968 219218 254010 219454
rect 254246 219218 254288 219454
rect 253968 219134 254288 219218
rect 253968 218898 254010 219134
rect 254246 218898 254288 219134
rect 253968 218866 254288 218898
rect 284688 219454 285008 219486
rect 284688 219218 284730 219454
rect 284966 219218 285008 219454
rect 284688 219134 285008 219218
rect 284688 218898 284730 219134
rect 284966 218898 285008 219134
rect 284688 218866 285008 218898
rect 315408 219454 315728 219486
rect 315408 219218 315450 219454
rect 315686 219218 315728 219454
rect 315408 219134 315728 219218
rect 315408 218898 315450 219134
rect 315686 218898 315728 219134
rect 315408 218866 315728 218898
rect 346128 219454 346448 219486
rect 346128 219218 346170 219454
rect 346406 219218 346448 219454
rect 346128 219134 346448 219218
rect 346128 218898 346170 219134
rect 346406 218898 346448 219134
rect 346128 218866 346448 218898
rect 376848 219454 377168 219486
rect 376848 219218 376890 219454
rect 377126 219218 377168 219454
rect 376848 219134 377168 219218
rect 376848 218898 376890 219134
rect 377126 218898 377168 219134
rect 376848 218866 377168 218898
rect 407568 219454 407888 219486
rect 407568 219218 407610 219454
rect 407846 219218 407888 219454
rect 407568 219134 407888 219218
rect 407568 218898 407610 219134
rect 407846 218898 407888 219134
rect 407568 218866 407888 218898
rect 438288 219454 438608 219486
rect 438288 219218 438330 219454
rect 438566 219218 438608 219454
rect 438288 219134 438608 219218
rect 438288 218898 438330 219134
rect 438566 218898 438608 219134
rect 438288 218866 438608 218898
rect 469008 219454 469328 219486
rect 469008 219218 469050 219454
rect 469286 219218 469328 219454
rect 469008 219134 469328 219218
rect 469008 218898 469050 219134
rect 469286 218898 469328 219134
rect 469008 218866 469328 218898
rect 499728 219454 500048 219486
rect 499728 219218 499770 219454
rect 500006 219218 500048 219454
rect 499728 219134 500048 219218
rect 499728 218898 499770 219134
rect 500006 218898 500048 219134
rect 499728 218866 500048 218898
rect 530448 219454 530768 219486
rect 530448 219218 530490 219454
rect 530726 219218 530768 219454
rect 530448 219134 530768 219218
rect 530448 218898 530490 219134
rect 530726 218898 530768 219134
rect 530448 218866 530768 218898
rect 561168 219454 561488 219486
rect 561168 219218 561210 219454
rect 561446 219218 561488 219454
rect 561168 219134 561488 219218
rect 561168 218898 561210 219134
rect 561446 218898 561488 219134
rect 561168 218866 561488 218898
rect 567234 208894 567854 244338
rect 567234 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 567854 208894
rect 567234 208574 567854 208658
rect 567234 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 567854 208574
rect 23568 201454 23888 201486
rect 23568 201218 23610 201454
rect 23846 201218 23888 201454
rect 23568 201134 23888 201218
rect 23568 200898 23610 201134
rect 23846 200898 23888 201134
rect 23568 200866 23888 200898
rect 54288 201454 54608 201486
rect 54288 201218 54330 201454
rect 54566 201218 54608 201454
rect 54288 201134 54608 201218
rect 54288 200898 54330 201134
rect 54566 200898 54608 201134
rect 54288 200866 54608 200898
rect 85008 201454 85328 201486
rect 85008 201218 85050 201454
rect 85286 201218 85328 201454
rect 85008 201134 85328 201218
rect 85008 200898 85050 201134
rect 85286 200898 85328 201134
rect 85008 200866 85328 200898
rect 115728 201454 116048 201486
rect 115728 201218 115770 201454
rect 116006 201218 116048 201454
rect 115728 201134 116048 201218
rect 115728 200898 115770 201134
rect 116006 200898 116048 201134
rect 115728 200866 116048 200898
rect 146448 201454 146768 201486
rect 146448 201218 146490 201454
rect 146726 201218 146768 201454
rect 146448 201134 146768 201218
rect 146448 200898 146490 201134
rect 146726 200898 146768 201134
rect 146448 200866 146768 200898
rect 177168 201454 177488 201486
rect 177168 201218 177210 201454
rect 177446 201218 177488 201454
rect 177168 201134 177488 201218
rect 177168 200898 177210 201134
rect 177446 200898 177488 201134
rect 177168 200866 177488 200898
rect 207888 201454 208208 201486
rect 207888 201218 207930 201454
rect 208166 201218 208208 201454
rect 207888 201134 208208 201218
rect 207888 200898 207930 201134
rect 208166 200898 208208 201134
rect 207888 200866 208208 200898
rect 238608 201454 238928 201486
rect 238608 201218 238650 201454
rect 238886 201218 238928 201454
rect 238608 201134 238928 201218
rect 238608 200898 238650 201134
rect 238886 200898 238928 201134
rect 238608 200866 238928 200898
rect 269328 201454 269648 201486
rect 269328 201218 269370 201454
rect 269606 201218 269648 201454
rect 269328 201134 269648 201218
rect 269328 200898 269370 201134
rect 269606 200898 269648 201134
rect 269328 200866 269648 200898
rect 300048 201454 300368 201486
rect 300048 201218 300090 201454
rect 300326 201218 300368 201454
rect 300048 201134 300368 201218
rect 300048 200898 300090 201134
rect 300326 200898 300368 201134
rect 300048 200866 300368 200898
rect 330768 201454 331088 201486
rect 330768 201218 330810 201454
rect 331046 201218 331088 201454
rect 330768 201134 331088 201218
rect 330768 200898 330810 201134
rect 331046 200898 331088 201134
rect 330768 200866 331088 200898
rect 361488 201454 361808 201486
rect 361488 201218 361530 201454
rect 361766 201218 361808 201454
rect 361488 201134 361808 201218
rect 361488 200898 361530 201134
rect 361766 200898 361808 201134
rect 361488 200866 361808 200898
rect 392208 201454 392528 201486
rect 392208 201218 392250 201454
rect 392486 201218 392528 201454
rect 392208 201134 392528 201218
rect 392208 200898 392250 201134
rect 392486 200898 392528 201134
rect 392208 200866 392528 200898
rect 422928 201454 423248 201486
rect 422928 201218 422970 201454
rect 423206 201218 423248 201454
rect 422928 201134 423248 201218
rect 422928 200898 422970 201134
rect 423206 200898 423248 201134
rect 422928 200866 423248 200898
rect 453648 201454 453968 201486
rect 453648 201218 453690 201454
rect 453926 201218 453968 201454
rect 453648 201134 453968 201218
rect 453648 200898 453690 201134
rect 453926 200898 453968 201134
rect 453648 200866 453968 200898
rect 484368 201454 484688 201486
rect 484368 201218 484410 201454
rect 484646 201218 484688 201454
rect 484368 201134 484688 201218
rect 484368 200898 484410 201134
rect 484646 200898 484688 201134
rect 484368 200866 484688 200898
rect 515088 201454 515408 201486
rect 515088 201218 515130 201454
rect 515366 201218 515408 201454
rect 515088 201134 515408 201218
rect 515088 200898 515130 201134
rect 515366 200898 515408 201134
rect 515088 200866 515408 200898
rect 545808 201454 546128 201486
rect 545808 201218 545850 201454
rect 546086 201218 546128 201454
rect 545808 201134 546128 201218
rect 545808 200898 545850 201134
rect 546086 200898 546128 201134
rect 545808 200866 546128 200898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect 8208 183454 8528 183486
rect 8208 183218 8250 183454
rect 8486 183218 8528 183454
rect 8208 183134 8528 183218
rect 8208 182898 8250 183134
rect 8486 182898 8528 183134
rect 8208 182866 8528 182898
rect 38928 183454 39248 183486
rect 38928 183218 38970 183454
rect 39206 183218 39248 183454
rect 38928 183134 39248 183218
rect 38928 182898 38970 183134
rect 39206 182898 39248 183134
rect 38928 182866 39248 182898
rect 69648 183454 69968 183486
rect 69648 183218 69690 183454
rect 69926 183218 69968 183454
rect 69648 183134 69968 183218
rect 69648 182898 69690 183134
rect 69926 182898 69968 183134
rect 69648 182866 69968 182898
rect 100368 183454 100688 183486
rect 100368 183218 100410 183454
rect 100646 183218 100688 183454
rect 100368 183134 100688 183218
rect 100368 182898 100410 183134
rect 100646 182898 100688 183134
rect 100368 182866 100688 182898
rect 131088 183454 131408 183486
rect 131088 183218 131130 183454
rect 131366 183218 131408 183454
rect 131088 183134 131408 183218
rect 131088 182898 131130 183134
rect 131366 182898 131408 183134
rect 131088 182866 131408 182898
rect 161808 183454 162128 183486
rect 161808 183218 161850 183454
rect 162086 183218 162128 183454
rect 161808 183134 162128 183218
rect 161808 182898 161850 183134
rect 162086 182898 162128 183134
rect 161808 182866 162128 182898
rect 192528 183454 192848 183486
rect 192528 183218 192570 183454
rect 192806 183218 192848 183454
rect 192528 183134 192848 183218
rect 192528 182898 192570 183134
rect 192806 182898 192848 183134
rect 192528 182866 192848 182898
rect 223248 183454 223568 183486
rect 223248 183218 223290 183454
rect 223526 183218 223568 183454
rect 223248 183134 223568 183218
rect 223248 182898 223290 183134
rect 223526 182898 223568 183134
rect 223248 182866 223568 182898
rect 253968 183454 254288 183486
rect 253968 183218 254010 183454
rect 254246 183218 254288 183454
rect 253968 183134 254288 183218
rect 253968 182898 254010 183134
rect 254246 182898 254288 183134
rect 253968 182866 254288 182898
rect 284688 183454 285008 183486
rect 284688 183218 284730 183454
rect 284966 183218 285008 183454
rect 284688 183134 285008 183218
rect 284688 182898 284730 183134
rect 284966 182898 285008 183134
rect 284688 182866 285008 182898
rect 315408 183454 315728 183486
rect 315408 183218 315450 183454
rect 315686 183218 315728 183454
rect 315408 183134 315728 183218
rect 315408 182898 315450 183134
rect 315686 182898 315728 183134
rect 315408 182866 315728 182898
rect 346128 183454 346448 183486
rect 346128 183218 346170 183454
rect 346406 183218 346448 183454
rect 346128 183134 346448 183218
rect 346128 182898 346170 183134
rect 346406 182898 346448 183134
rect 346128 182866 346448 182898
rect 376848 183454 377168 183486
rect 376848 183218 376890 183454
rect 377126 183218 377168 183454
rect 376848 183134 377168 183218
rect 376848 182898 376890 183134
rect 377126 182898 377168 183134
rect 376848 182866 377168 182898
rect 407568 183454 407888 183486
rect 407568 183218 407610 183454
rect 407846 183218 407888 183454
rect 407568 183134 407888 183218
rect 407568 182898 407610 183134
rect 407846 182898 407888 183134
rect 407568 182866 407888 182898
rect 438288 183454 438608 183486
rect 438288 183218 438330 183454
rect 438566 183218 438608 183454
rect 438288 183134 438608 183218
rect 438288 182898 438330 183134
rect 438566 182898 438608 183134
rect 438288 182866 438608 182898
rect 469008 183454 469328 183486
rect 469008 183218 469050 183454
rect 469286 183218 469328 183454
rect 469008 183134 469328 183218
rect 469008 182898 469050 183134
rect 469286 182898 469328 183134
rect 469008 182866 469328 182898
rect 499728 183454 500048 183486
rect 499728 183218 499770 183454
rect 500006 183218 500048 183454
rect 499728 183134 500048 183218
rect 499728 182898 499770 183134
rect 500006 182898 500048 183134
rect 499728 182866 500048 182898
rect 530448 183454 530768 183486
rect 530448 183218 530490 183454
rect 530726 183218 530768 183454
rect 530448 183134 530768 183218
rect 530448 182898 530490 183134
rect 530726 182898 530768 183134
rect 530448 182866 530768 182898
rect 561168 183454 561488 183486
rect 561168 183218 561210 183454
rect 561446 183218 561488 183454
rect 561168 183134 561488 183218
rect 561168 182898 561210 183134
rect 561446 182898 561488 183134
rect 561168 182866 561488 182898
rect 567234 172894 567854 208338
rect 567234 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 567854 172894
rect 567234 172574 567854 172658
rect 567234 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 567854 172574
rect 23568 165454 23888 165486
rect 23568 165218 23610 165454
rect 23846 165218 23888 165454
rect 23568 165134 23888 165218
rect 23568 164898 23610 165134
rect 23846 164898 23888 165134
rect 23568 164866 23888 164898
rect 54288 165454 54608 165486
rect 54288 165218 54330 165454
rect 54566 165218 54608 165454
rect 54288 165134 54608 165218
rect 54288 164898 54330 165134
rect 54566 164898 54608 165134
rect 54288 164866 54608 164898
rect 85008 165454 85328 165486
rect 85008 165218 85050 165454
rect 85286 165218 85328 165454
rect 85008 165134 85328 165218
rect 85008 164898 85050 165134
rect 85286 164898 85328 165134
rect 85008 164866 85328 164898
rect 115728 165454 116048 165486
rect 115728 165218 115770 165454
rect 116006 165218 116048 165454
rect 115728 165134 116048 165218
rect 115728 164898 115770 165134
rect 116006 164898 116048 165134
rect 115728 164866 116048 164898
rect 146448 165454 146768 165486
rect 146448 165218 146490 165454
rect 146726 165218 146768 165454
rect 146448 165134 146768 165218
rect 146448 164898 146490 165134
rect 146726 164898 146768 165134
rect 146448 164866 146768 164898
rect 177168 165454 177488 165486
rect 177168 165218 177210 165454
rect 177446 165218 177488 165454
rect 177168 165134 177488 165218
rect 177168 164898 177210 165134
rect 177446 164898 177488 165134
rect 177168 164866 177488 164898
rect 207888 165454 208208 165486
rect 207888 165218 207930 165454
rect 208166 165218 208208 165454
rect 207888 165134 208208 165218
rect 207888 164898 207930 165134
rect 208166 164898 208208 165134
rect 207888 164866 208208 164898
rect 238608 165454 238928 165486
rect 238608 165218 238650 165454
rect 238886 165218 238928 165454
rect 238608 165134 238928 165218
rect 238608 164898 238650 165134
rect 238886 164898 238928 165134
rect 238608 164866 238928 164898
rect 269328 165454 269648 165486
rect 269328 165218 269370 165454
rect 269606 165218 269648 165454
rect 269328 165134 269648 165218
rect 269328 164898 269370 165134
rect 269606 164898 269648 165134
rect 269328 164866 269648 164898
rect 300048 165454 300368 165486
rect 300048 165218 300090 165454
rect 300326 165218 300368 165454
rect 300048 165134 300368 165218
rect 300048 164898 300090 165134
rect 300326 164898 300368 165134
rect 300048 164866 300368 164898
rect 330768 165454 331088 165486
rect 330768 165218 330810 165454
rect 331046 165218 331088 165454
rect 330768 165134 331088 165218
rect 330768 164898 330810 165134
rect 331046 164898 331088 165134
rect 330768 164866 331088 164898
rect 361488 165454 361808 165486
rect 361488 165218 361530 165454
rect 361766 165218 361808 165454
rect 361488 165134 361808 165218
rect 361488 164898 361530 165134
rect 361766 164898 361808 165134
rect 361488 164866 361808 164898
rect 392208 165454 392528 165486
rect 392208 165218 392250 165454
rect 392486 165218 392528 165454
rect 392208 165134 392528 165218
rect 392208 164898 392250 165134
rect 392486 164898 392528 165134
rect 392208 164866 392528 164898
rect 422928 165454 423248 165486
rect 422928 165218 422970 165454
rect 423206 165218 423248 165454
rect 422928 165134 423248 165218
rect 422928 164898 422970 165134
rect 423206 164898 423248 165134
rect 422928 164866 423248 164898
rect 453648 165454 453968 165486
rect 453648 165218 453690 165454
rect 453926 165218 453968 165454
rect 453648 165134 453968 165218
rect 453648 164898 453690 165134
rect 453926 164898 453968 165134
rect 453648 164866 453968 164898
rect 484368 165454 484688 165486
rect 484368 165218 484410 165454
rect 484646 165218 484688 165454
rect 484368 165134 484688 165218
rect 484368 164898 484410 165134
rect 484646 164898 484688 165134
rect 484368 164866 484688 164898
rect 515088 165454 515408 165486
rect 515088 165218 515130 165454
rect 515366 165218 515408 165454
rect 515088 165134 515408 165218
rect 515088 164898 515130 165134
rect 515366 164898 515408 165134
rect 515088 164866 515408 164898
rect 545808 165454 546128 165486
rect 545808 165218 545850 165454
rect 546086 165218 546128 165454
rect 545808 165134 546128 165218
rect 545808 164898 545850 165134
rect 546086 164898 546128 165134
rect 545808 164866 546128 164898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect 8208 147454 8528 147486
rect 8208 147218 8250 147454
rect 8486 147218 8528 147454
rect 8208 147134 8528 147218
rect 8208 146898 8250 147134
rect 8486 146898 8528 147134
rect 8208 146866 8528 146898
rect 38928 147454 39248 147486
rect 38928 147218 38970 147454
rect 39206 147218 39248 147454
rect 38928 147134 39248 147218
rect 38928 146898 38970 147134
rect 39206 146898 39248 147134
rect 38928 146866 39248 146898
rect 69648 147454 69968 147486
rect 69648 147218 69690 147454
rect 69926 147218 69968 147454
rect 69648 147134 69968 147218
rect 69648 146898 69690 147134
rect 69926 146898 69968 147134
rect 69648 146866 69968 146898
rect 100368 147454 100688 147486
rect 100368 147218 100410 147454
rect 100646 147218 100688 147454
rect 100368 147134 100688 147218
rect 100368 146898 100410 147134
rect 100646 146898 100688 147134
rect 100368 146866 100688 146898
rect 131088 147454 131408 147486
rect 131088 147218 131130 147454
rect 131366 147218 131408 147454
rect 131088 147134 131408 147218
rect 131088 146898 131130 147134
rect 131366 146898 131408 147134
rect 131088 146866 131408 146898
rect 161808 147454 162128 147486
rect 161808 147218 161850 147454
rect 162086 147218 162128 147454
rect 161808 147134 162128 147218
rect 161808 146898 161850 147134
rect 162086 146898 162128 147134
rect 161808 146866 162128 146898
rect 192528 147454 192848 147486
rect 192528 147218 192570 147454
rect 192806 147218 192848 147454
rect 192528 147134 192848 147218
rect 192528 146898 192570 147134
rect 192806 146898 192848 147134
rect 192528 146866 192848 146898
rect 223248 147454 223568 147486
rect 223248 147218 223290 147454
rect 223526 147218 223568 147454
rect 223248 147134 223568 147218
rect 223248 146898 223290 147134
rect 223526 146898 223568 147134
rect 223248 146866 223568 146898
rect 253968 147454 254288 147486
rect 253968 147218 254010 147454
rect 254246 147218 254288 147454
rect 253968 147134 254288 147218
rect 253968 146898 254010 147134
rect 254246 146898 254288 147134
rect 253968 146866 254288 146898
rect 284688 147454 285008 147486
rect 284688 147218 284730 147454
rect 284966 147218 285008 147454
rect 284688 147134 285008 147218
rect 284688 146898 284730 147134
rect 284966 146898 285008 147134
rect 284688 146866 285008 146898
rect 315408 147454 315728 147486
rect 315408 147218 315450 147454
rect 315686 147218 315728 147454
rect 315408 147134 315728 147218
rect 315408 146898 315450 147134
rect 315686 146898 315728 147134
rect 315408 146866 315728 146898
rect 346128 147454 346448 147486
rect 346128 147218 346170 147454
rect 346406 147218 346448 147454
rect 346128 147134 346448 147218
rect 346128 146898 346170 147134
rect 346406 146898 346448 147134
rect 346128 146866 346448 146898
rect 376848 147454 377168 147486
rect 376848 147218 376890 147454
rect 377126 147218 377168 147454
rect 376848 147134 377168 147218
rect 376848 146898 376890 147134
rect 377126 146898 377168 147134
rect 376848 146866 377168 146898
rect 407568 147454 407888 147486
rect 407568 147218 407610 147454
rect 407846 147218 407888 147454
rect 407568 147134 407888 147218
rect 407568 146898 407610 147134
rect 407846 146898 407888 147134
rect 407568 146866 407888 146898
rect 438288 147454 438608 147486
rect 438288 147218 438330 147454
rect 438566 147218 438608 147454
rect 438288 147134 438608 147218
rect 438288 146898 438330 147134
rect 438566 146898 438608 147134
rect 438288 146866 438608 146898
rect 469008 147454 469328 147486
rect 469008 147218 469050 147454
rect 469286 147218 469328 147454
rect 469008 147134 469328 147218
rect 469008 146898 469050 147134
rect 469286 146898 469328 147134
rect 469008 146866 469328 146898
rect 499728 147454 500048 147486
rect 499728 147218 499770 147454
rect 500006 147218 500048 147454
rect 499728 147134 500048 147218
rect 499728 146898 499770 147134
rect 500006 146898 500048 147134
rect 499728 146866 500048 146898
rect 530448 147454 530768 147486
rect 530448 147218 530490 147454
rect 530726 147218 530768 147454
rect 530448 147134 530768 147218
rect 530448 146898 530490 147134
rect 530726 146898 530768 147134
rect 530448 146866 530768 146898
rect 561168 147454 561488 147486
rect 561168 147218 561210 147454
rect 561446 147218 561488 147454
rect 561168 147134 561488 147218
rect 561168 146898 561210 147134
rect 561446 146898 561488 147134
rect 561168 146866 561488 146898
rect 567234 136894 567854 172338
rect 567234 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 567854 136894
rect 567234 136574 567854 136658
rect 567234 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 567854 136574
rect 23568 129454 23888 129486
rect 23568 129218 23610 129454
rect 23846 129218 23888 129454
rect 23568 129134 23888 129218
rect 23568 128898 23610 129134
rect 23846 128898 23888 129134
rect 23568 128866 23888 128898
rect 54288 129454 54608 129486
rect 54288 129218 54330 129454
rect 54566 129218 54608 129454
rect 54288 129134 54608 129218
rect 54288 128898 54330 129134
rect 54566 128898 54608 129134
rect 54288 128866 54608 128898
rect 85008 129454 85328 129486
rect 85008 129218 85050 129454
rect 85286 129218 85328 129454
rect 85008 129134 85328 129218
rect 85008 128898 85050 129134
rect 85286 128898 85328 129134
rect 85008 128866 85328 128898
rect 115728 129454 116048 129486
rect 115728 129218 115770 129454
rect 116006 129218 116048 129454
rect 115728 129134 116048 129218
rect 115728 128898 115770 129134
rect 116006 128898 116048 129134
rect 115728 128866 116048 128898
rect 146448 129454 146768 129486
rect 146448 129218 146490 129454
rect 146726 129218 146768 129454
rect 146448 129134 146768 129218
rect 146448 128898 146490 129134
rect 146726 128898 146768 129134
rect 146448 128866 146768 128898
rect 177168 129454 177488 129486
rect 177168 129218 177210 129454
rect 177446 129218 177488 129454
rect 177168 129134 177488 129218
rect 177168 128898 177210 129134
rect 177446 128898 177488 129134
rect 177168 128866 177488 128898
rect 207888 129454 208208 129486
rect 207888 129218 207930 129454
rect 208166 129218 208208 129454
rect 207888 129134 208208 129218
rect 207888 128898 207930 129134
rect 208166 128898 208208 129134
rect 207888 128866 208208 128898
rect 238608 129454 238928 129486
rect 238608 129218 238650 129454
rect 238886 129218 238928 129454
rect 238608 129134 238928 129218
rect 238608 128898 238650 129134
rect 238886 128898 238928 129134
rect 238608 128866 238928 128898
rect 269328 129454 269648 129486
rect 269328 129218 269370 129454
rect 269606 129218 269648 129454
rect 269328 129134 269648 129218
rect 269328 128898 269370 129134
rect 269606 128898 269648 129134
rect 269328 128866 269648 128898
rect 300048 129454 300368 129486
rect 300048 129218 300090 129454
rect 300326 129218 300368 129454
rect 300048 129134 300368 129218
rect 300048 128898 300090 129134
rect 300326 128898 300368 129134
rect 300048 128866 300368 128898
rect 330768 129454 331088 129486
rect 330768 129218 330810 129454
rect 331046 129218 331088 129454
rect 330768 129134 331088 129218
rect 330768 128898 330810 129134
rect 331046 128898 331088 129134
rect 330768 128866 331088 128898
rect 361488 129454 361808 129486
rect 361488 129218 361530 129454
rect 361766 129218 361808 129454
rect 361488 129134 361808 129218
rect 361488 128898 361530 129134
rect 361766 128898 361808 129134
rect 361488 128866 361808 128898
rect 392208 129454 392528 129486
rect 392208 129218 392250 129454
rect 392486 129218 392528 129454
rect 392208 129134 392528 129218
rect 392208 128898 392250 129134
rect 392486 128898 392528 129134
rect 392208 128866 392528 128898
rect 422928 129454 423248 129486
rect 422928 129218 422970 129454
rect 423206 129218 423248 129454
rect 422928 129134 423248 129218
rect 422928 128898 422970 129134
rect 423206 128898 423248 129134
rect 422928 128866 423248 128898
rect 453648 129454 453968 129486
rect 453648 129218 453690 129454
rect 453926 129218 453968 129454
rect 453648 129134 453968 129218
rect 453648 128898 453690 129134
rect 453926 128898 453968 129134
rect 453648 128866 453968 128898
rect 484368 129454 484688 129486
rect 484368 129218 484410 129454
rect 484646 129218 484688 129454
rect 484368 129134 484688 129218
rect 484368 128898 484410 129134
rect 484646 128898 484688 129134
rect 484368 128866 484688 128898
rect 515088 129454 515408 129486
rect 515088 129218 515130 129454
rect 515366 129218 515408 129454
rect 515088 129134 515408 129218
rect 515088 128898 515130 129134
rect 515366 128898 515408 129134
rect 515088 128866 515408 128898
rect 545808 129454 546128 129486
rect 545808 129218 545850 129454
rect 546086 129218 546128 129454
rect 545808 129134 546128 129218
rect 545808 128898 545850 129134
rect 546086 128898 546128 129134
rect 545808 128866 546128 128898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect 8208 111454 8528 111486
rect 8208 111218 8250 111454
rect 8486 111218 8528 111454
rect 8208 111134 8528 111218
rect 8208 110898 8250 111134
rect 8486 110898 8528 111134
rect 8208 110866 8528 110898
rect 38928 111454 39248 111486
rect 38928 111218 38970 111454
rect 39206 111218 39248 111454
rect 38928 111134 39248 111218
rect 38928 110898 38970 111134
rect 39206 110898 39248 111134
rect 38928 110866 39248 110898
rect 69648 111454 69968 111486
rect 69648 111218 69690 111454
rect 69926 111218 69968 111454
rect 69648 111134 69968 111218
rect 69648 110898 69690 111134
rect 69926 110898 69968 111134
rect 69648 110866 69968 110898
rect 100368 111454 100688 111486
rect 100368 111218 100410 111454
rect 100646 111218 100688 111454
rect 100368 111134 100688 111218
rect 100368 110898 100410 111134
rect 100646 110898 100688 111134
rect 100368 110866 100688 110898
rect 131088 111454 131408 111486
rect 131088 111218 131130 111454
rect 131366 111218 131408 111454
rect 131088 111134 131408 111218
rect 131088 110898 131130 111134
rect 131366 110898 131408 111134
rect 131088 110866 131408 110898
rect 161808 111454 162128 111486
rect 161808 111218 161850 111454
rect 162086 111218 162128 111454
rect 161808 111134 162128 111218
rect 161808 110898 161850 111134
rect 162086 110898 162128 111134
rect 161808 110866 162128 110898
rect 192528 111454 192848 111486
rect 192528 111218 192570 111454
rect 192806 111218 192848 111454
rect 192528 111134 192848 111218
rect 192528 110898 192570 111134
rect 192806 110898 192848 111134
rect 192528 110866 192848 110898
rect 223248 111454 223568 111486
rect 223248 111218 223290 111454
rect 223526 111218 223568 111454
rect 223248 111134 223568 111218
rect 223248 110898 223290 111134
rect 223526 110898 223568 111134
rect 223248 110866 223568 110898
rect 253968 111454 254288 111486
rect 253968 111218 254010 111454
rect 254246 111218 254288 111454
rect 253968 111134 254288 111218
rect 253968 110898 254010 111134
rect 254246 110898 254288 111134
rect 253968 110866 254288 110898
rect 284688 111454 285008 111486
rect 284688 111218 284730 111454
rect 284966 111218 285008 111454
rect 284688 111134 285008 111218
rect 284688 110898 284730 111134
rect 284966 110898 285008 111134
rect 284688 110866 285008 110898
rect 315408 111454 315728 111486
rect 315408 111218 315450 111454
rect 315686 111218 315728 111454
rect 315408 111134 315728 111218
rect 315408 110898 315450 111134
rect 315686 110898 315728 111134
rect 315408 110866 315728 110898
rect 346128 111454 346448 111486
rect 346128 111218 346170 111454
rect 346406 111218 346448 111454
rect 346128 111134 346448 111218
rect 346128 110898 346170 111134
rect 346406 110898 346448 111134
rect 346128 110866 346448 110898
rect 376848 111454 377168 111486
rect 376848 111218 376890 111454
rect 377126 111218 377168 111454
rect 376848 111134 377168 111218
rect 376848 110898 376890 111134
rect 377126 110898 377168 111134
rect 376848 110866 377168 110898
rect 407568 111454 407888 111486
rect 407568 111218 407610 111454
rect 407846 111218 407888 111454
rect 407568 111134 407888 111218
rect 407568 110898 407610 111134
rect 407846 110898 407888 111134
rect 407568 110866 407888 110898
rect 438288 111454 438608 111486
rect 438288 111218 438330 111454
rect 438566 111218 438608 111454
rect 438288 111134 438608 111218
rect 438288 110898 438330 111134
rect 438566 110898 438608 111134
rect 438288 110866 438608 110898
rect 469008 111454 469328 111486
rect 469008 111218 469050 111454
rect 469286 111218 469328 111454
rect 469008 111134 469328 111218
rect 469008 110898 469050 111134
rect 469286 110898 469328 111134
rect 469008 110866 469328 110898
rect 499728 111454 500048 111486
rect 499728 111218 499770 111454
rect 500006 111218 500048 111454
rect 499728 111134 500048 111218
rect 499728 110898 499770 111134
rect 500006 110898 500048 111134
rect 499728 110866 500048 110898
rect 530448 111454 530768 111486
rect 530448 111218 530490 111454
rect 530726 111218 530768 111454
rect 530448 111134 530768 111218
rect 530448 110898 530490 111134
rect 530726 110898 530768 111134
rect 530448 110866 530768 110898
rect 561168 111454 561488 111486
rect 561168 111218 561210 111454
rect 561446 111218 561488 111454
rect 561168 111134 561488 111218
rect 561168 110898 561210 111134
rect 561446 110898 561488 111134
rect 561168 110866 561488 110898
rect 567234 100894 567854 136338
rect 567234 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 567854 100894
rect 567234 100574 567854 100658
rect 567234 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 567854 100574
rect 23568 93454 23888 93486
rect 23568 93218 23610 93454
rect 23846 93218 23888 93454
rect 23568 93134 23888 93218
rect 23568 92898 23610 93134
rect 23846 92898 23888 93134
rect 23568 92866 23888 92898
rect 54288 93454 54608 93486
rect 54288 93218 54330 93454
rect 54566 93218 54608 93454
rect 54288 93134 54608 93218
rect 54288 92898 54330 93134
rect 54566 92898 54608 93134
rect 54288 92866 54608 92898
rect 85008 93454 85328 93486
rect 85008 93218 85050 93454
rect 85286 93218 85328 93454
rect 85008 93134 85328 93218
rect 85008 92898 85050 93134
rect 85286 92898 85328 93134
rect 85008 92866 85328 92898
rect 115728 93454 116048 93486
rect 115728 93218 115770 93454
rect 116006 93218 116048 93454
rect 115728 93134 116048 93218
rect 115728 92898 115770 93134
rect 116006 92898 116048 93134
rect 115728 92866 116048 92898
rect 146448 93454 146768 93486
rect 146448 93218 146490 93454
rect 146726 93218 146768 93454
rect 146448 93134 146768 93218
rect 146448 92898 146490 93134
rect 146726 92898 146768 93134
rect 146448 92866 146768 92898
rect 177168 93454 177488 93486
rect 177168 93218 177210 93454
rect 177446 93218 177488 93454
rect 177168 93134 177488 93218
rect 177168 92898 177210 93134
rect 177446 92898 177488 93134
rect 177168 92866 177488 92898
rect 207888 93454 208208 93486
rect 207888 93218 207930 93454
rect 208166 93218 208208 93454
rect 207888 93134 208208 93218
rect 207888 92898 207930 93134
rect 208166 92898 208208 93134
rect 207888 92866 208208 92898
rect 238608 93454 238928 93486
rect 238608 93218 238650 93454
rect 238886 93218 238928 93454
rect 238608 93134 238928 93218
rect 238608 92898 238650 93134
rect 238886 92898 238928 93134
rect 238608 92866 238928 92898
rect 269328 93454 269648 93486
rect 269328 93218 269370 93454
rect 269606 93218 269648 93454
rect 269328 93134 269648 93218
rect 269328 92898 269370 93134
rect 269606 92898 269648 93134
rect 269328 92866 269648 92898
rect 300048 93454 300368 93486
rect 300048 93218 300090 93454
rect 300326 93218 300368 93454
rect 300048 93134 300368 93218
rect 300048 92898 300090 93134
rect 300326 92898 300368 93134
rect 300048 92866 300368 92898
rect 330768 93454 331088 93486
rect 330768 93218 330810 93454
rect 331046 93218 331088 93454
rect 330768 93134 331088 93218
rect 330768 92898 330810 93134
rect 331046 92898 331088 93134
rect 330768 92866 331088 92898
rect 361488 93454 361808 93486
rect 361488 93218 361530 93454
rect 361766 93218 361808 93454
rect 361488 93134 361808 93218
rect 361488 92898 361530 93134
rect 361766 92898 361808 93134
rect 361488 92866 361808 92898
rect 392208 93454 392528 93486
rect 392208 93218 392250 93454
rect 392486 93218 392528 93454
rect 392208 93134 392528 93218
rect 392208 92898 392250 93134
rect 392486 92898 392528 93134
rect 392208 92866 392528 92898
rect 422928 93454 423248 93486
rect 422928 93218 422970 93454
rect 423206 93218 423248 93454
rect 422928 93134 423248 93218
rect 422928 92898 422970 93134
rect 423206 92898 423248 93134
rect 422928 92866 423248 92898
rect 453648 93454 453968 93486
rect 453648 93218 453690 93454
rect 453926 93218 453968 93454
rect 453648 93134 453968 93218
rect 453648 92898 453690 93134
rect 453926 92898 453968 93134
rect 453648 92866 453968 92898
rect 484368 93454 484688 93486
rect 484368 93218 484410 93454
rect 484646 93218 484688 93454
rect 484368 93134 484688 93218
rect 484368 92898 484410 93134
rect 484646 92898 484688 93134
rect 484368 92866 484688 92898
rect 515088 93454 515408 93486
rect 515088 93218 515130 93454
rect 515366 93218 515408 93454
rect 515088 93134 515408 93218
rect 515088 92898 515130 93134
rect 515366 92898 515408 93134
rect 515088 92866 515408 92898
rect 545808 93454 546128 93486
rect 545808 93218 545850 93454
rect 546086 93218 546128 93454
rect 545808 93134 546128 93218
rect 545808 92898 545850 93134
rect 546086 92898 546128 93134
rect 545808 92866 546128 92898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect 8208 75454 8528 75486
rect 8208 75218 8250 75454
rect 8486 75218 8528 75454
rect 8208 75134 8528 75218
rect 8208 74898 8250 75134
rect 8486 74898 8528 75134
rect 8208 74866 8528 74898
rect 38928 75454 39248 75486
rect 38928 75218 38970 75454
rect 39206 75218 39248 75454
rect 38928 75134 39248 75218
rect 38928 74898 38970 75134
rect 39206 74898 39248 75134
rect 38928 74866 39248 74898
rect 69648 75454 69968 75486
rect 69648 75218 69690 75454
rect 69926 75218 69968 75454
rect 69648 75134 69968 75218
rect 69648 74898 69690 75134
rect 69926 74898 69968 75134
rect 69648 74866 69968 74898
rect 100368 75454 100688 75486
rect 100368 75218 100410 75454
rect 100646 75218 100688 75454
rect 100368 75134 100688 75218
rect 100368 74898 100410 75134
rect 100646 74898 100688 75134
rect 100368 74866 100688 74898
rect 131088 75454 131408 75486
rect 131088 75218 131130 75454
rect 131366 75218 131408 75454
rect 131088 75134 131408 75218
rect 131088 74898 131130 75134
rect 131366 74898 131408 75134
rect 131088 74866 131408 74898
rect 161808 75454 162128 75486
rect 161808 75218 161850 75454
rect 162086 75218 162128 75454
rect 161808 75134 162128 75218
rect 161808 74898 161850 75134
rect 162086 74898 162128 75134
rect 161808 74866 162128 74898
rect 192528 75454 192848 75486
rect 192528 75218 192570 75454
rect 192806 75218 192848 75454
rect 192528 75134 192848 75218
rect 192528 74898 192570 75134
rect 192806 74898 192848 75134
rect 192528 74866 192848 74898
rect 223248 75454 223568 75486
rect 223248 75218 223290 75454
rect 223526 75218 223568 75454
rect 223248 75134 223568 75218
rect 223248 74898 223290 75134
rect 223526 74898 223568 75134
rect 223248 74866 223568 74898
rect 253968 75454 254288 75486
rect 253968 75218 254010 75454
rect 254246 75218 254288 75454
rect 253968 75134 254288 75218
rect 253968 74898 254010 75134
rect 254246 74898 254288 75134
rect 253968 74866 254288 74898
rect 284688 75454 285008 75486
rect 284688 75218 284730 75454
rect 284966 75218 285008 75454
rect 284688 75134 285008 75218
rect 284688 74898 284730 75134
rect 284966 74898 285008 75134
rect 284688 74866 285008 74898
rect 315408 75454 315728 75486
rect 315408 75218 315450 75454
rect 315686 75218 315728 75454
rect 315408 75134 315728 75218
rect 315408 74898 315450 75134
rect 315686 74898 315728 75134
rect 315408 74866 315728 74898
rect 346128 75454 346448 75486
rect 346128 75218 346170 75454
rect 346406 75218 346448 75454
rect 346128 75134 346448 75218
rect 346128 74898 346170 75134
rect 346406 74898 346448 75134
rect 346128 74866 346448 74898
rect 376848 75454 377168 75486
rect 376848 75218 376890 75454
rect 377126 75218 377168 75454
rect 376848 75134 377168 75218
rect 376848 74898 376890 75134
rect 377126 74898 377168 75134
rect 376848 74866 377168 74898
rect 407568 75454 407888 75486
rect 407568 75218 407610 75454
rect 407846 75218 407888 75454
rect 407568 75134 407888 75218
rect 407568 74898 407610 75134
rect 407846 74898 407888 75134
rect 407568 74866 407888 74898
rect 438288 75454 438608 75486
rect 438288 75218 438330 75454
rect 438566 75218 438608 75454
rect 438288 75134 438608 75218
rect 438288 74898 438330 75134
rect 438566 74898 438608 75134
rect 438288 74866 438608 74898
rect 469008 75454 469328 75486
rect 469008 75218 469050 75454
rect 469286 75218 469328 75454
rect 469008 75134 469328 75218
rect 469008 74898 469050 75134
rect 469286 74898 469328 75134
rect 469008 74866 469328 74898
rect 499728 75454 500048 75486
rect 499728 75218 499770 75454
rect 500006 75218 500048 75454
rect 499728 75134 500048 75218
rect 499728 74898 499770 75134
rect 500006 74898 500048 75134
rect 499728 74866 500048 74898
rect 530448 75454 530768 75486
rect 530448 75218 530490 75454
rect 530726 75218 530768 75454
rect 530448 75134 530768 75218
rect 530448 74898 530490 75134
rect 530726 74898 530768 75134
rect 530448 74866 530768 74898
rect 561168 75454 561488 75486
rect 561168 75218 561210 75454
rect 561446 75218 561488 75454
rect 561168 75134 561488 75218
rect 561168 74898 561210 75134
rect 561446 74898 561488 75134
rect 561168 74866 561488 74898
rect 567234 64894 567854 100338
rect 567234 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 567854 64894
rect 567234 64574 567854 64658
rect 567234 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 567854 64574
rect 23568 57454 23888 57486
rect 23568 57218 23610 57454
rect 23846 57218 23888 57454
rect 23568 57134 23888 57218
rect 23568 56898 23610 57134
rect 23846 56898 23888 57134
rect 23568 56866 23888 56898
rect 54288 57454 54608 57486
rect 54288 57218 54330 57454
rect 54566 57218 54608 57454
rect 54288 57134 54608 57218
rect 54288 56898 54330 57134
rect 54566 56898 54608 57134
rect 54288 56866 54608 56898
rect 85008 57454 85328 57486
rect 85008 57218 85050 57454
rect 85286 57218 85328 57454
rect 85008 57134 85328 57218
rect 85008 56898 85050 57134
rect 85286 56898 85328 57134
rect 85008 56866 85328 56898
rect 115728 57454 116048 57486
rect 115728 57218 115770 57454
rect 116006 57218 116048 57454
rect 115728 57134 116048 57218
rect 115728 56898 115770 57134
rect 116006 56898 116048 57134
rect 115728 56866 116048 56898
rect 146448 57454 146768 57486
rect 146448 57218 146490 57454
rect 146726 57218 146768 57454
rect 146448 57134 146768 57218
rect 146448 56898 146490 57134
rect 146726 56898 146768 57134
rect 146448 56866 146768 56898
rect 177168 57454 177488 57486
rect 177168 57218 177210 57454
rect 177446 57218 177488 57454
rect 177168 57134 177488 57218
rect 177168 56898 177210 57134
rect 177446 56898 177488 57134
rect 177168 56866 177488 56898
rect 207888 57454 208208 57486
rect 207888 57218 207930 57454
rect 208166 57218 208208 57454
rect 207888 57134 208208 57218
rect 207888 56898 207930 57134
rect 208166 56898 208208 57134
rect 207888 56866 208208 56898
rect 238608 57454 238928 57486
rect 238608 57218 238650 57454
rect 238886 57218 238928 57454
rect 238608 57134 238928 57218
rect 238608 56898 238650 57134
rect 238886 56898 238928 57134
rect 238608 56866 238928 56898
rect 269328 57454 269648 57486
rect 269328 57218 269370 57454
rect 269606 57218 269648 57454
rect 269328 57134 269648 57218
rect 269328 56898 269370 57134
rect 269606 56898 269648 57134
rect 269328 56866 269648 56898
rect 300048 57454 300368 57486
rect 300048 57218 300090 57454
rect 300326 57218 300368 57454
rect 300048 57134 300368 57218
rect 300048 56898 300090 57134
rect 300326 56898 300368 57134
rect 300048 56866 300368 56898
rect 330768 57454 331088 57486
rect 330768 57218 330810 57454
rect 331046 57218 331088 57454
rect 330768 57134 331088 57218
rect 330768 56898 330810 57134
rect 331046 56898 331088 57134
rect 330768 56866 331088 56898
rect 361488 57454 361808 57486
rect 361488 57218 361530 57454
rect 361766 57218 361808 57454
rect 361488 57134 361808 57218
rect 361488 56898 361530 57134
rect 361766 56898 361808 57134
rect 361488 56866 361808 56898
rect 392208 57454 392528 57486
rect 392208 57218 392250 57454
rect 392486 57218 392528 57454
rect 392208 57134 392528 57218
rect 392208 56898 392250 57134
rect 392486 56898 392528 57134
rect 392208 56866 392528 56898
rect 422928 57454 423248 57486
rect 422928 57218 422970 57454
rect 423206 57218 423248 57454
rect 422928 57134 423248 57218
rect 422928 56898 422970 57134
rect 423206 56898 423248 57134
rect 422928 56866 423248 56898
rect 453648 57454 453968 57486
rect 453648 57218 453690 57454
rect 453926 57218 453968 57454
rect 453648 57134 453968 57218
rect 453648 56898 453690 57134
rect 453926 56898 453968 57134
rect 453648 56866 453968 56898
rect 484368 57454 484688 57486
rect 484368 57218 484410 57454
rect 484646 57218 484688 57454
rect 484368 57134 484688 57218
rect 484368 56898 484410 57134
rect 484646 56898 484688 57134
rect 484368 56866 484688 56898
rect 515088 57454 515408 57486
rect 515088 57218 515130 57454
rect 515366 57218 515408 57454
rect 515088 57134 515408 57218
rect 515088 56898 515130 57134
rect 515366 56898 515408 57134
rect 515088 56866 515408 56898
rect 545808 57454 546128 57486
rect 545808 57218 545850 57454
rect 546086 57218 546128 57454
rect 545808 57134 546128 57218
rect 545808 56898 545850 57134
rect 546086 56898 546128 57134
rect 545808 56866 546128 56898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect 8208 39454 8528 39486
rect 8208 39218 8250 39454
rect 8486 39218 8528 39454
rect 8208 39134 8528 39218
rect 8208 38898 8250 39134
rect 8486 38898 8528 39134
rect 8208 38866 8528 38898
rect 38928 39454 39248 39486
rect 38928 39218 38970 39454
rect 39206 39218 39248 39454
rect 38928 39134 39248 39218
rect 38928 38898 38970 39134
rect 39206 38898 39248 39134
rect 38928 38866 39248 38898
rect 69648 39454 69968 39486
rect 69648 39218 69690 39454
rect 69926 39218 69968 39454
rect 69648 39134 69968 39218
rect 69648 38898 69690 39134
rect 69926 38898 69968 39134
rect 69648 38866 69968 38898
rect 100368 39454 100688 39486
rect 100368 39218 100410 39454
rect 100646 39218 100688 39454
rect 100368 39134 100688 39218
rect 100368 38898 100410 39134
rect 100646 38898 100688 39134
rect 100368 38866 100688 38898
rect 131088 39454 131408 39486
rect 131088 39218 131130 39454
rect 131366 39218 131408 39454
rect 131088 39134 131408 39218
rect 131088 38898 131130 39134
rect 131366 38898 131408 39134
rect 131088 38866 131408 38898
rect 161808 39454 162128 39486
rect 161808 39218 161850 39454
rect 162086 39218 162128 39454
rect 161808 39134 162128 39218
rect 161808 38898 161850 39134
rect 162086 38898 162128 39134
rect 161808 38866 162128 38898
rect 192528 39454 192848 39486
rect 192528 39218 192570 39454
rect 192806 39218 192848 39454
rect 192528 39134 192848 39218
rect 192528 38898 192570 39134
rect 192806 38898 192848 39134
rect 192528 38866 192848 38898
rect 223248 39454 223568 39486
rect 223248 39218 223290 39454
rect 223526 39218 223568 39454
rect 223248 39134 223568 39218
rect 223248 38898 223290 39134
rect 223526 38898 223568 39134
rect 223248 38866 223568 38898
rect 253968 39454 254288 39486
rect 253968 39218 254010 39454
rect 254246 39218 254288 39454
rect 253968 39134 254288 39218
rect 253968 38898 254010 39134
rect 254246 38898 254288 39134
rect 253968 38866 254288 38898
rect 284688 39454 285008 39486
rect 284688 39218 284730 39454
rect 284966 39218 285008 39454
rect 284688 39134 285008 39218
rect 284688 38898 284730 39134
rect 284966 38898 285008 39134
rect 284688 38866 285008 38898
rect 315408 39454 315728 39486
rect 315408 39218 315450 39454
rect 315686 39218 315728 39454
rect 315408 39134 315728 39218
rect 315408 38898 315450 39134
rect 315686 38898 315728 39134
rect 315408 38866 315728 38898
rect 346128 39454 346448 39486
rect 346128 39218 346170 39454
rect 346406 39218 346448 39454
rect 346128 39134 346448 39218
rect 346128 38898 346170 39134
rect 346406 38898 346448 39134
rect 346128 38866 346448 38898
rect 376848 39454 377168 39486
rect 376848 39218 376890 39454
rect 377126 39218 377168 39454
rect 376848 39134 377168 39218
rect 376848 38898 376890 39134
rect 377126 38898 377168 39134
rect 376848 38866 377168 38898
rect 407568 39454 407888 39486
rect 407568 39218 407610 39454
rect 407846 39218 407888 39454
rect 407568 39134 407888 39218
rect 407568 38898 407610 39134
rect 407846 38898 407888 39134
rect 407568 38866 407888 38898
rect 438288 39454 438608 39486
rect 438288 39218 438330 39454
rect 438566 39218 438608 39454
rect 438288 39134 438608 39218
rect 438288 38898 438330 39134
rect 438566 38898 438608 39134
rect 438288 38866 438608 38898
rect 469008 39454 469328 39486
rect 469008 39218 469050 39454
rect 469286 39218 469328 39454
rect 469008 39134 469328 39218
rect 469008 38898 469050 39134
rect 469286 38898 469328 39134
rect 469008 38866 469328 38898
rect 499728 39454 500048 39486
rect 499728 39218 499770 39454
rect 500006 39218 500048 39454
rect 499728 39134 500048 39218
rect 499728 38898 499770 39134
rect 500006 38898 500048 39134
rect 499728 38866 500048 38898
rect 530448 39454 530768 39486
rect 530448 39218 530490 39454
rect 530726 39218 530768 39454
rect 530448 39134 530768 39218
rect 530448 38898 530490 39134
rect 530726 38898 530768 39134
rect 530448 38866 530768 38898
rect 561168 39454 561488 39486
rect 561168 39218 561210 39454
rect 561446 39218 561488 39454
rect 561168 39134 561488 39218
rect 561168 38898 561210 39134
rect 561446 38898 561488 39134
rect 561168 38866 561488 38898
rect 567234 28894 567854 64338
rect 567234 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 567854 28894
rect 567234 28574 567854 28658
rect 567234 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 567854 28574
rect 23568 21454 23888 21486
rect 23568 21218 23610 21454
rect 23846 21218 23888 21454
rect 23568 21134 23888 21218
rect 23568 20898 23610 21134
rect 23846 20898 23888 21134
rect 23568 20866 23888 20898
rect 54288 21454 54608 21486
rect 54288 21218 54330 21454
rect 54566 21218 54608 21454
rect 54288 21134 54608 21218
rect 54288 20898 54330 21134
rect 54566 20898 54608 21134
rect 54288 20866 54608 20898
rect 85008 21454 85328 21486
rect 85008 21218 85050 21454
rect 85286 21218 85328 21454
rect 85008 21134 85328 21218
rect 85008 20898 85050 21134
rect 85286 20898 85328 21134
rect 85008 20866 85328 20898
rect 115728 21454 116048 21486
rect 115728 21218 115770 21454
rect 116006 21218 116048 21454
rect 115728 21134 116048 21218
rect 115728 20898 115770 21134
rect 116006 20898 116048 21134
rect 115728 20866 116048 20898
rect 146448 21454 146768 21486
rect 146448 21218 146490 21454
rect 146726 21218 146768 21454
rect 146448 21134 146768 21218
rect 146448 20898 146490 21134
rect 146726 20898 146768 21134
rect 146448 20866 146768 20898
rect 177168 21454 177488 21486
rect 177168 21218 177210 21454
rect 177446 21218 177488 21454
rect 177168 21134 177488 21218
rect 177168 20898 177210 21134
rect 177446 20898 177488 21134
rect 177168 20866 177488 20898
rect 207888 21454 208208 21486
rect 207888 21218 207930 21454
rect 208166 21218 208208 21454
rect 207888 21134 208208 21218
rect 207888 20898 207930 21134
rect 208166 20898 208208 21134
rect 207888 20866 208208 20898
rect 238608 21454 238928 21486
rect 238608 21218 238650 21454
rect 238886 21218 238928 21454
rect 238608 21134 238928 21218
rect 238608 20898 238650 21134
rect 238886 20898 238928 21134
rect 238608 20866 238928 20898
rect 269328 21454 269648 21486
rect 269328 21218 269370 21454
rect 269606 21218 269648 21454
rect 269328 21134 269648 21218
rect 269328 20898 269370 21134
rect 269606 20898 269648 21134
rect 269328 20866 269648 20898
rect 300048 21454 300368 21486
rect 300048 21218 300090 21454
rect 300326 21218 300368 21454
rect 300048 21134 300368 21218
rect 300048 20898 300090 21134
rect 300326 20898 300368 21134
rect 300048 20866 300368 20898
rect 330768 21454 331088 21486
rect 330768 21218 330810 21454
rect 331046 21218 331088 21454
rect 330768 21134 331088 21218
rect 330768 20898 330810 21134
rect 331046 20898 331088 21134
rect 330768 20866 331088 20898
rect 361488 21454 361808 21486
rect 361488 21218 361530 21454
rect 361766 21218 361808 21454
rect 361488 21134 361808 21218
rect 361488 20898 361530 21134
rect 361766 20898 361808 21134
rect 361488 20866 361808 20898
rect 392208 21454 392528 21486
rect 392208 21218 392250 21454
rect 392486 21218 392528 21454
rect 392208 21134 392528 21218
rect 392208 20898 392250 21134
rect 392486 20898 392528 21134
rect 392208 20866 392528 20898
rect 422928 21454 423248 21486
rect 422928 21218 422970 21454
rect 423206 21218 423248 21454
rect 422928 21134 423248 21218
rect 422928 20898 422970 21134
rect 423206 20898 423248 21134
rect 422928 20866 423248 20898
rect 453648 21454 453968 21486
rect 453648 21218 453690 21454
rect 453926 21218 453968 21454
rect 453648 21134 453968 21218
rect 453648 20898 453690 21134
rect 453926 20898 453968 21134
rect 453648 20866 453968 20898
rect 484368 21454 484688 21486
rect 484368 21218 484410 21454
rect 484646 21218 484688 21454
rect 484368 21134 484688 21218
rect 484368 20898 484410 21134
rect 484646 20898 484688 21134
rect 484368 20866 484688 20898
rect 515088 21454 515408 21486
rect 515088 21218 515130 21454
rect 515366 21218 515408 21454
rect 515088 21134 515408 21218
rect 515088 20898 515130 21134
rect 515366 20898 515408 21134
rect 515088 20866 515408 20898
rect 545808 21454 546128 21486
rect 545808 21218 545850 21454
rect 546086 21218 546128 21454
rect 545808 21134 546128 21218
rect 545808 20898 545850 21134
rect 546086 20898 546128 21134
rect 545808 20866 546128 20898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect 8208 3454 8528 3486
rect 8208 3218 8250 3454
rect 8486 3218 8528 3454
rect 8208 3134 8528 3218
rect 8208 2898 8250 3134
rect 8486 2898 8528 3134
rect 8208 2866 8528 2898
rect 38928 3454 39248 3486
rect 38928 3218 38970 3454
rect 39206 3218 39248 3454
rect 38928 3134 39248 3218
rect 38928 2898 38970 3134
rect 39206 2898 39248 3134
rect 38928 2866 39248 2898
rect 69648 3454 69968 3486
rect 69648 3218 69690 3454
rect 69926 3218 69968 3454
rect 69648 3134 69968 3218
rect 69648 2898 69690 3134
rect 69926 2898 69968 3134
rect 69648 2866 69968 2898
rect 100368 3454 100688 3486
rect 100368 3218 100410 3454
rect 100646 3218 100688 3454
rect 100368 3134 100688 3218
rect 100368 2898 100410 3134
rect 100646 2898 100688 3134
rect 100368 2866 100688 2898
rect 131088 3454 131408 3486
rect 131088 3218 131130 3454
rect 131366 3218 131408 3454
rect 131088 3134 131408 3218
rect 131088 2898 131130 3134
rect 131366 2898 131408 3134
rect 131088 2866 131408 2898
rect 161808 3454 162128 3486
rect 161808 3218 161850 3454
rect 162086 3218 162128 3454
rect 161808 3134 162128 3218
rect 161808 2898 161850 3134
rect 162086 2898 162128 3134
rect 161808 2866 162128 2898
rect 192528 3454 192848 3486
rect 192528 3218 192570 3454
rect 192806 3218 192848 3454
rect 192528 3134 192848 3218
rect 192528 2898 192570 3134
rect 192806 2898 192848 3134
rect 192528 2866 192848 2898
rect 223248 3454 223568 3486
rect 223248 3218 223290 3454
rect 223526 3218 223568 3454
rect 223248 3134 223568 3218
rect 223248 2898 223290 3134
rect 223526 2898 223568 3134
rect 223248 2866 223568 2898
rect 253968 3454 254288 3486
rect 253968 3218 254010 3454
rect 254246 3218 254288 3454
rect 253968 3134 254288 3218
rect 253968 2898 254010 3134
rect 254246 2898 254288 3134
rect 253968 2866 254288 2898
rect 284688 3454 285008 3486
rect 284688 3218 284730 3454
rect 284966 3218 285008 3454
rect 284688 3134 285008 3218
rect 284688 2898 284730 3134
rect 284966 2898 285008 3134
rect 284688 2866 285008 2898
rect 315408 3454 315728 3486
rect 315408 3218 315450 3454
rect 315686 3218 315728 3454
rect 315408 3134 315728 3218
rect 315408 2898 315450 3134
rect 315686 2898 315728 3134
rect 315408 2866 315728 2898
rect 346128 3454 346448 3486
rect 346128 3218 346170 3454
rect 346406 3218 346448 3454
rect 346128 3134 346448 3218
rect 346128 2898 346170 3134
rect 346406 2898 346448 3134
rect 346128 2866 346448 2898
rect 376848 3454 377168 3486
rect 376848 3218 376890 3454
rect 377126 3218 377168 3454
rect 376848 3134 377168 3218
rect 376848 2898 376890 3134
rect 377126 2898 377168 3134
rect 376848 2866 377168 2898
rect 407568 3454 407888 3486
rect 407568 3218 407610 3454
rect 407846 3218 407888 3454
rect 407568 3134 407888 3218
rect 407568 2898 407610 3134
rect 407846 2898 407888 3134
rect 407568 2866 407888 2898
rect 438288 3454 438608 3486
rect 438288 3218 438330 3454
rect 438566 3218 438608 3454
rect 438288 3134 438608 3218
rect 438288 2898 438330 3134
rect 438566 2898 438608 3134
rect 438288 2866 438608 2898
rect 469008 3454 469328 3486
rect 469008 3218 469050 3454
rect 469286 3218 469328 3454
rect 469008 3134 469328 3218
rect 469008 2898 469050 3134
rect 469286 2898 469328 3134
rect 469008 2866 469328 2898
rect 499728 3454 500048 3486
rect 499728 3218 499770 3454
rect 500006 3218 500048 3454
rect 499728 3134 500048 3218
rect 499728 2898 499770 3134
rect 500006 2898 500048 3134
rect 499728 2866 500048 2898
rect 530448 3454 530768 3486
rect 530448 3218 530490 3454
rect 530726 3218 530768 3454
rect 530448 3134 530768 3218
rect 530448 2898 530490 3134
rect 530726 2898 530768 3134
rect 530448 2866 530768 2898
rect 561168 3454 561488 3486
rect 561168 3218 561210 3454
rect 561446 3218 561488 3454
rect 561168 3134 561488 3218
rect 561168 2898 561210 3134
rect 561446 2898 561488 3134
rect 561168 2866 561488 2898
rect 551323 916 551389 917
rect 551323 852 551324 916
rect 551388 852 551389 916
rect 551323 851 551389 852
rect 551326 645 551386 851
rect 551323 644 551389 645
rect 551323 580 551324 644
rect 551388 580 551389 644
rect 551323 579 551389 580
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 -2000
rect 5514 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 6134 -2266
rect 5514 -2586 6134 -2502
rect 5514 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 6134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 -2000
rect 9234 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 9854 -4186
rect 9234 -4506 9854 -4422
rect 9234 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 9854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 -2000
rect 23514 -3226 24134 -2000
rect 23514 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 24134 -3226
rect 23514 -3546 24134 -3462
rect 23514 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 24134 -3546
rect 23514 -3814 24134 -3782
rect 27234 -5146 27854 -2000
rect 27234 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 27854 -5146
rect 27234 -5466 27854 -5382
rect 27234 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 27854 -5466
rect 27234 -5734 27854 -5702
rect 12954 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 13574 -6106
rect 12954 -6426 13574 -6342
rect 12954 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 13574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 -2000
rect 41514 -2266 42134 -2000
rect 41514 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 42134 -2266
rect 41514 -2586 42134 -2502
rect 41514 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 42134 -2586
rect 41514 -3814 42134 -2822
rect 45234 -4186 45854 -2000
rect 45234 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 45854 -4186
rect 45234 -4506 45854 -4422
rect 45234 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 45854 -4506
rect 45234 -5734 45854 -4742
rect 30954 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 31574 -7066
rect 30954 -7386 31574 -7302
rect 30954 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 31574 -7386
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 -2000
rect 59514 -3226 60134 -2000
rect 59514 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 60134 -3226
rect 59514 -3546 60134 -3462
rect 59514 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 60134 -3546
rect 59514 -3814 60134 -3782
rect 63234 -5146 63854 -2000
rect 63234 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 63854 -5146
rect 63234 -5466 63854 -5382
rect 63234 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 63854 -5466
rect 63234 -5734 63854 -5702
rect 48954 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 49574 -6106
rect 48954 -6426 49574 -6342
rect 48954 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 49574 -6426
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 -2000
rect 77514 -2266 78134 -2000
rect 77514 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 78134 -2266
rect 77514 -2586 78134 -2502
rect 77514 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 78134 -2586
rect 77514 -3814 78134 -2822
rect 81234 -4186 81854 -2000
rect 81234 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 81854 -4186
rect 81234 -4506 81854 -4422
rect 81234 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 81854 -4506
rect 81234 -5734 81854 -4742
rect 66954 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 67574 -7066
rect 66954 -7386 67574 -7302
rect 66954 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 67574 -7386
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 -2000
rect 95514 -3226 96134 -2000
rect 95514 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 96134 -3226
rect 95514 -3546 96134 -3462
rect 95514 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 96134 -3546
rect 95514 -3814 96134 -3782
rect 99234 -5146 99854 -2000
rect 99234 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 99854 -5146
rect 99234 -5466 99854 -5382
rect 99234 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 99854 -5466
rect 99234 -5734 99854 -5702
rect 84954 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 85574 -6106
rect 84954 -6426 85574 -6342
rect 84954 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 85574 -6426
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 -2000
rect 113514 -2266 114134 -2000
rect 113514 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 114134 -2266
rect 113514 -2586 114134 -2502
rect 113514 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 114134 -2586
rect 113514 -3814 114134 -2822
rect 117234 -4186 117854 -2000
rect 117234 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 117854 -4186
rect 117234 -4506 117854 -4422
rect 117234 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 117854 -4506
rect 117234 -5734 117854 -4742
rect 102954 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 103574 -7066
rect 102954 -7386 103574 -7302
rect 102954 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 103574 -7386
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 -2000
rect 131514 -3226 132134 -2000
rect 131514 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 132134 -3226
rect 131514 -3546 132134 -3462
rect 131514 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 132134 -3546
rect 131514 -3814 132134 -3782
rect 135234 -5146 135854 -2000
rect 135234 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 135854 -5146
rect 135234 -5466 135854 -5382
rect 135234 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 135854 -5466
rect 135234 -5734 135854 -5702
rect 120954 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 121574 -6106
rect 120954 -6426 121574 -6342
rect 120954 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 121574 -6426
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 -2000
rect 149514 -2266 150134 -2000
rect 149514 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 150134 -2266
rect 149514 -2586 150134 -2502
rect 149514 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 150134 -2586
rect 149514 -3814 150134 -2822
rect 153234 -4186 153854 -2000
rect 153234 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 153854 -4186
rect 153234 -4506 153854 -4422
rect 153234 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 153854 -4506
rect 153234 -5734 153854 -4742
rect 138954 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 139574 -7066
rect 138954 -7386 139574 -7302
rect 138954 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 139574 -7386
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 -2000
rect 167514 -3226 168134 -2000
rect 167514 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 168134 -3226
rect 167514 -3546 168134 -3462
rect 167514 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 168134 -3546
rect 167514 -3814 168134 -3782
rect 171234 -5146 171854 -2000
rect 171234 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 171854 -5146
rect 171234 -5466 171854 -5382
rect 171234 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 171854 -5466
rect 171234 -5734 171854 -5702
rect 156954 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 157574 -6106
rect 156954 -6426 157574 -6342
rect 156954 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 157574 -6426
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 -2000
rect 185514 -2266 186134 -2000
rect 185514 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 186134 -2266
rect 185514 -2586 186134 -2502
rect 185514 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 186134 -2586
rect 185514 -3814 186134 -2822
rect 189234 -4186 189854 -2000
rect 189234 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 189854 -4186
rect 189234 -4506 189854 -4422
rect 189234 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 189854 -4506
rect 189234 -5734 189854 -4742
rect 174954 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 175574 -7066
rect 174954 -7386 175574 -7302
rect 174954 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 175574 -7386
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 -2000
rect 203514 -3226 204134 -2000
rect 203514 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 204134 -3226
rect 203514 -3546 204134 -3462
rect 203514 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 204134 -3546
rect 203514 -3814 204134 -3782
rect 207234 -5146 207854 -2000
rect 207234 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 207854 -5146
rect 207234 -5466 207854 -5382
rect 207234 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 207854 -5466
rect 207234 -5734 207854 -5702
rect 192954 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 193574 -6106
rect 192954 -6426 193574 -6342
rect 192954 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 193574 -6426
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 -2000
rect 221514 -2266 222134 -2000
rect 221514 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 222134 -2266
rect 221514 -2586 222134 -2502
rect 221514 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 222134 -2586
rect 221514 -3814 222134 -2822
rect 225234 -4186 225854 -2000
rect 225234 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 225854 -4186
rect 225234 -4506 225854 -4422
rect 225234 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 225854 -4506
rect 225234 -5734 225854 -4742
rect 210954 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 211574 -7066
rect 210954 -7386 211574 -7302
rect 210954 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 211574 -7386
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 -2000
rect 239514 -3226 240134 -2000
rect 239514 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 240134 -3226
rect 239514 -3546 240134 -3462
rect 239514 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 240134 -3546
rect 239514 -3814 240134 -3782
rect 243234 -5146 243854 -2000
rect 243234 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 243854 -5146
rect 243234 -5466 243854 -5382
rect 243234 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 243854 -5466
rect 243234 -5734 243854 -5702
rect 228954 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 229574 -6106
rect 228954 -6426 229574 -6342
rect 228954 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 229574 -6426
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 -2000
rect 257514 -2266 258134 -2000
rect 257514 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 258134 -2266
rect 257514 -2586 258134 -2502
rect 257514 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 258134 -2586
rect 257514 -3814 258134 -2822
rect 261234 -4186 261854 -2000
rect 261234 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 261854 -4186
rect 261234 -4506 261854 -4422
rect 261234 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 261854 -4506
rect 261234 -5734 261854 -4742
rect 246954 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 247574 -7066
rect 246954 -7386 247574 -7302
rect 246954 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 247574 -7386
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 -2000
rect 275514 -3226 276134 -2000
rect 275514 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 276134 -3226
rect 275514 -3546 276134 -3462
rect 275514 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 276134 -3546
rect 275514 -3814 276134 -3782
rect 279234 -5146 279854 -2000
rect 279234 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 279854 -5146
rect 279234 -5466 279854 -5382
rect 279234 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 279854 -5466
rect 279234 -5734 279854 -5702
rect 264954 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 265574 -6106
rect 264954 -6426 265574 -6342
rect 264954 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 265574 -6426
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 -2000
rect 293514 -2266 294134 -2000
rect 293514 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 294134 -2266
rect 293514 -2586 294134 -2502
rect 293514 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 294134 -2586
rect 293514 -3814 294134 -2822
rect 297234 -4186 297854 -2000
rect 297234 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 297854 -4186
rect 297234 -4506 297854 -4422
rect 297234 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 297854 -4506
rect 297234 -5734 297854 -4742
rect 282954 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 283574 -7066
rect 282954 -7386 283574 -7302
rect 282954 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 283574 -7386
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 -2000
rect 311514 -3226 312134 -2000
rect 311514 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 312134 -3226
rect 311514 -3546 312134 -3462
rect 311514 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 312134 -3546
rect 311514 -3814 312134 -3782
rect 315234 -5146 315854 -2000
rect 315234 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 315854 -5146
rect 315234 -5466 315854 -5382
rect 315234 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 315854 -5466
rect 315234 -5734 315854 -5702
rect 300954 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 301574 -6106
rect 300954 -6426 301574 -6342
rect 300954 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 301574 -6426
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 -2000
rect 329514 -2266 330134 -2000
rect 329514 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 330134 -2266
rect 329514 -2586 330134 -2502
rect 329514 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 330134 -2586
rect 329514 -3814 330134 -2822
rect 333234 -4186 333854 -2000
rect 333234 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 333854 -4186
rect 333234 -4506 333854 -4422
rect 333234 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 333854 -4506
rect 333234 -5734 333854 -4742
rect 318954 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 319574 -7066
rect 318954 -7386 319574 -7302
rect 318954 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 319574 -7386
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 -2000
rect 347514 -3226 348134 -2000
rect 347514 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 348134 -3226
rect 347514 -3546 348134 -3462
rect 347514 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 348134 -3546
rect 347514 -3814 348134 -3782
rect 351234 -5146 351854 -2000
rect 351234 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 351854 -5146
rect 351234 -5466 351854 -5382
rect 351234 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 351854 -5466
rect 351234 -5734 351854 -5702
rect 336954 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 337574 -6106
rect 336954 -6426 337574 -6342
rect 336954 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 337574 -6426
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 -2000
rect 365514 -2266 366134 -2000
rect 365514 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 366134 -2266
rect 365514 -2586 366134 -2502
rect 365514 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 366134 -2586
rect 365514 -3814 366134 -2822
rect 369234 -4186 369854 -2000
rect 369234 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 369854 -4186
rect 369234 -4506 369854 -4422
rect 369234 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 369854 -4506
rect 369234 -5734 369854 -4742
rect 354954 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 355574 -7066
rect 354954 -7386 355574 -7302
rect 354954 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 355574 -7386
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 -2000
rect 383514 -3226 384134 -2000
rect 383514 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 384134 -3226
rect 383514 -3546 384134 -3462
rect 383514 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 384134 -3546
rect 383514 -3814 384134 -3782
rect 387234 -5146 387854 -2000
rect 387234 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 387854 -5146
rect 387234 -5466 387854 -5382
rect 387234 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 387854 -5466
rect 387234 -5734 387854 -5702
rect 372954 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 373574 -6106
rect 372954 -6426 373574 -6342
rect 372954 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 373574 -6426
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 -2000
rect 401514 -2266 402134 -2000
rect 401514 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 402134 -2266
rect 401514 -2586 402134 -2502
rect 401514 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 402134 -2586
rect 401514 -3814 402134 -2822
rect 405234 -4186 405854 -2000
rect 405234 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 405854 -4186
rect 405234 -4506 405854 -4422
rect 405234 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 405854 -4506
rect 405234 -5734 405854 -4742
rect 390954 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 391574 -7066
rect 390954 -7386 391574 -7302
rect 390954 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 391574 -7386
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 -2000
rect 419514 -3226 420134 -2000
rect 419514 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 420134 -3226
rect 419514 -3546 420134 -3462
rect 419514 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 420134 -3546
rect 419514 -3814 420134 -3782
rect 423234 -5146 423854 -2000
rect 423234 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 423854 -5146
rect 423234 -5466 423854 -5382
rect 423234 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 423854 -5466
rect 423234 -5734 423854 -5702
rect 408954 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 409574 -6106
rect 408954 -6426 409574 -6342
rect 408954 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 409574 -6426
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 -2000
rect 437514 -2266 438134 -2000
rect 437514 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 438134 -2266
rect 437514 -2586 438134 -2502
rect 437514 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 438134 -2586
rect 437514 -3814 438134 -2822
rect 441234 -4186 441854 -2000
rect 441234 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 441854 -4186
rect 441234 -4506 441854 -4422
rect 441234 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 441854 -4506
rect 441234 -5734 441854 -4742
rect 426954 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 427574 -7066
rect 426954 -7386 427574 -7302
rect 426954 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 427574 -7386
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 -2000
rect 455514 -3226 456134 -2000
rect 455514 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 456134 -3226
rect 455514 -3546 456134 -3462
rect 455514 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 456134 -3546
rect 455514 -3814 456134 -3782
rect 459234 -5146 459854 -2000
rect 459234 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 459854 -5146
rect 459234 -5466 459854 -5382
rect 459234 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 459854 -5466
rect 459234 -5734 459854 -5702
rect 444954 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 445574 -6106
rect 444954 -6426 445574 -6342
rect 444954 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 445574 -6426
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 -2000
rect 473514 -2266 474134 -2000
rect 473514 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 474134 -2266
rect 473514 -2586 474134 -2502
rect 473514 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 474134 -2586
rect 473514 -3814 474134 -2822
rect 477234 -4186 477854 -2000
rect 477234 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 477854 -4186
rect 477234 -4506 477854 -4422
rect 477234 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 477854 -4506
rect 477234 -5734 477854 -4742
rect 462954 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 463574 -7066
rect 462954 -7386 463574 -7302
rect 462954 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 463574 -7386
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 -2000
rect 491514 -3226 492134 -2000
rect 491514 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 492134 -3226
rect 491514 -3546 492134 -3462
rect 491514 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 492134 -3546
rect 491514 -3814 492134 -3782
rect 495234 -5146 495854 -2000
rect 495234 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 495854 -5146
rect 495234 -5466 495854 -5382
rect 495234 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 495854 -5466
rect 495234 -5734 495854 -5702
rect 480954 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 481574 -6106
rect 480954 -6426 481574 -6342
rect 480954 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 481574 -6426
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 -2000
rect 509514 -2266 510134 -2000
rect 509514 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 510134 -2266
rect 509514 -2586 510134 -2502
rect 509514 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 510134 -2586
rect 509514 -3814 510134 -2822
rect 513234 -4186 513854 -2000
rect 513234 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 513854 -4186
rect 513234 -4506 513854 -4422
rect 513234 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 513854 -4506
rect 513234 -5734 513854 -4742
rect 498954 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 499574 -7066
rect 498954 -7386 499574 -7302
rect 498954 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 499574 -7386
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 -2000
rect 527514 -3226 528134 -2000
rect 527514 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 528134 -3226
rect 527514 -3546 528134 -3462
rect 527514 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 528134 -3546
rect 527514 -3814 528134 -3782
rect 531234 -5146 531854 -2000
rect 531234 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 531854 -5146
rect 531234 -5466 531854 -5382
rect 531234 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 531854 -5466
rect 531234 -5734 531854 -5702
rect 516954 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 517574 -6106
rect 516954 -6426 517574 -6342
rect 516954 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 517574 -6426
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 -2000
rect 545514 -2266 546134 -2000
rect 545514 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 546134 -2266
rect 545514 -2586 546134 -2502
rect 545514 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 546134 -2586
rect 545514 -3814 546134 -2822
rect 549234 -4186 549854 -2000
rect 549234 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 549854 -4186
rect 549234 -4506 549854 -4422
rect 549234 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 549854 -4506
rect 549234 -5734 549854 -4742
rect 534954 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 535574 -7066
rect 534954 -7386 535574 -7302
rect 534954 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 535574 -7386
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 -2000
rect 563514 -3226 564134 -2000
rect 563514 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 564134 -3226
rect 563514 -3546 564134 -3462
rect 563514 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 564134 -3546
rect 563514 -3814 564134 -3782
rect 567234 -5146 567854 28338
rect 567234 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 567854 -5146
rect 567234 -5466 567854 -5382
rect 567234 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 567854 -5466
rect 567234 -5734 567854 -5702
rect 570954 680614 571574 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 581514 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 582134 706758
rect 581514 706438 582134 706522
rect 581514 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 582134 706438
rect 570954 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 571574 680614
rect 570954 680294 571574 680378
rect 570954 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 571574 680294
rect 570954 644614 571574 680058
rect 570954 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 571574 644614
rect 570954 644294 571574 644378
rect 570954 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 571574 644294
rect 570954 608614 571574 644058
rect 570954 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 571574 608614
rect 570954 608294 571574 608378
rect 570954 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 571574 608294
rect 570954 572614 571574 608058
rect 570954 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 571574 572614
rect 570954 572294 571574 572378
rect 570954 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 571574 572294
rect 570954 536614 571574 572058
rect 570954 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 571574 536614
rect 570954 536294 571574 536378
rect 570954 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 571574 536294
rect 570954 500614 571574 536058
rect 570954 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 571574 500614
rect 570954 500294 571574 500378
rect 570954 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 571574 500294
rect 570954 464614 571574 500058
rect 570954 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 571574 464614
rect 570954 464294 571574 464378
rect 570954 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 571574 464294
rect 570954 428614 571574 464058
rect 570954 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 571574 428614
rect 570954 428294 571574 428378
rect 570954 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 571574 428294
rect 570954 392614 571574 428058
rect 570954 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 571574 392614
rect 570954 392294 571574 392378
rect 570954 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 571574 392294
rect 570954 356614 571574 392058
rect 570954 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 571574 356614
rect 570954 356294 571574 356378
rect 570954 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 571574 356294
rect 570954 320614 571574 356058
rect 570954 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 571574 320614
rect 570954 320294 571574 320378
rect 570954 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 571574 320294
rect 570954 284614 571574 320058
rect 570954 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 571574 284614
rect 570954 284294 571574 284378
rect 570954 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 571574 284294
rect 570954 248614 571574 284058
rect 570954 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 571574 248614
rect 570954 248294 571574 248378
rect 570954 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 571574 248294
rect 570954 212614 571574 248058
rect 570954 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 571574 212614
rect 570954 212294 571574 212378
rect 570954 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 571574 212294
rect 570954 176614 571574 212058
rect 570954 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 571574 176614
rect 570954 176294 571574 176378
rect 570954 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 571574 176294
rect 570954 140614 571574 176058
rect 570954 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 571574 140614
rect 570954 140294 571574 140378
rect 570954 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 571574 140294
rect 570954 104614 571574 140058
rect 570954 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 571574 104614
rect 570954 104294 571574 104378
rect 570954 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 571574 104294
rect 570954 68614 571574 104058
rect 570954 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 571574 68614
rect 570954 68294 571574 68378
rect 570954 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 571574 68294
rect 570954 32614 571574 68058
rect 570954 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 571574 32614
rect 570954 32294 571574 32378
rect 570954 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 571574 32294
rect 552954 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 553574 -6106
rect 552954 -6426 553574 -6342
rect 552954 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 553574 -6426
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 32058
rect 577794 704838 578414 705830
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 581514 691174 582134 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -2266 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 587850 691174
rect 587230 690854 587850 690938
rect 587230 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 587850 690854
rect 587230 655174 587850 690618
rect 587230 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 587850 655174
rect 587230 654854 587850 654938
rect 587230 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 587850 654854
rect 587230 619174 587850 654618
rect 587230 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 587850 619174
rect 587230 618854 587850 618938
rect 587230 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 587850 618854
rect 587230 583174 587850 618618
rect 587230 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 587850 583174
rect 587230 582854 587850 582938
rect 587230 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 587850 582854
rect 587230 547174 587850 582618
rect 587230 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 587850 547174
rect 587230 546854 587850 546938
rect 587230 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 587850 546854
rect 587230 511174 587850 546618
rect 587230 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 587850 511174
rect 587230 510854 587850 510938
rect 587230 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 587850 510854
rect 587230 475174 587850 510618
rect 587230 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 587850 475174
rect 587230 474854 587850 474938
rect 587230 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 587850 474854
rect 587230 439174 587850 474618
rect 587230 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 587850 439174
rect 587230 438854 587850 438938
rect 587230 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 587850 438854
rect 587230 403174 587850 438618
rect 587230 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 587850 403174
rect 587230 402854 587850 402938
rect 587230 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 587850 402854
rect 587230 367174 587850 402618
rect 587230 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 587850 367174
rect 587230 366854 587850 366938
rect 587230 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 587850 366854
rect 587230 331174 587850 366618
rect 587230 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 587850 331174
rect 587230 330854 587850 330938
rect 587230 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 587850 330854
rect 587230 295174 587850 330618
rect 587230 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 587850 295174
rect 587230 294854 587850 294938
rect 587230 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 587850 294854
rect 587230 259174 587850 294618
rect 587230 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 587850 259174
rect 587230 258854 587850 258938
rect 587230 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 587850 258854
rect 587230 223174 587850 258618
rect 587230 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 587850 223174
rect 587230 222854 587850 222938
rect 587230 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 587850 222854
rect 587230 187174 587850 222618
rect 587230 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 587850 187174
rect 587230 186854 587850 186938
rect 587230 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 587850 186854
rect 587230 151174 587850 186618
rect 587230 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 587850 151174
rect 587230 150854 587850 150938
rect 587230 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 587850 150854
rect 587230 115174 587850 150618
rect 587230 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 587850 115174
rect 587230 114854 587850 114938
rect 587230 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 587850 114854
rect 587230 79174 587850 114618
rect 587230 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 587850 79174
rect 587230 78854 587850 78938
rect 587230 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 587850 78854
rect 587230 43174 587850 78618
rect 587230 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 587850 43174
rect 587230 42854 587850 42938
rect 587230 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 587850 42854
rect 587230 7174 587850 42618
rect 587230 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 587850 7174
rect 587230 6854 587850 6938
rect 587230 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 587850 6854
rect 581514 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 582134 -2266
rect 581514 -2586 582134 -2502
rect 581514 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 582134 -2586
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect 588190 672854 588810 672938
rect 588190 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect 588190 637174 588810 672618
rect 588190 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect 588190 636854 588810 636938
rect 588190 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect 588190 601174 588810 636618
rect 588190 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect 588190 600854 588810 600938
rect 588190 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect 588190 565174 588810 600618
rect 588190 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect 588190 564854 588810 564938
rect 588190 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect 588190 529174 588810 564618
rect 588190 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect 588190 528854 588810 528938
rect 588190 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect 588190 493174 588810 528618
rect 588190 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect 588190 492854 588810 492938
rect 588190 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect 588190 457174 588810 492618
rect 588190 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect 588190 456854 588810 456938
rect 588190 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect 588190 421174 588810 456618
rect 588190 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 588190 420854 588810 420938
rect 588190 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 588190 385174 588810 420618
rect 588190 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 588190 384854 588810 384938
rect 588190 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 588190 349174 588810 384618
rect 588190 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 588190 348854 588810 348938
rect 588190 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 588190 313174 588810 348618
rect 588190 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 588190 312854 588810 312938
rect 588190 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 588190 277174 588810 312618
rect 588190 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 588190 276854 588810 276938
rect 588190 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 588190 241174 588810 276618
rect 588190 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 588190 240854 588810 240938
rect 588190 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 588190 205174 588810 240618
rect 588190 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 588190 204854 588810 204938
rect 588190 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 588190 169174 588810 204618
rect 588190 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 588190 168854 588810 168938
rect 588190 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 588190 133174 588810 168618
rect 588190 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 588190 132854 588810 132938
rect 588190 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 588190 97174 588810 132618
rect 588190 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 588190 96854 588810 96938
rect 588190 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 588190 61174 588810 96618
rect 588190 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 588190 60854 588810 60938
rect 588190 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 588190 25174 588810 60618
rect 588190 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect 588190 24854 588810 24938
rect 588190 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect 588190 -3226 588810 24618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 589770 694894
rect 589150 694574 589770 694658
rect 589150 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 589770 694574
rect 589150 658894 589770 694338
rect 589150 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 589770 658894
rect 589150 658574 589770 658658
rect 589150 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 589770 658574
rect 589150 622894 589770 658338
rect 589150 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 589770 622894
rect 589150 622574 589770 622658
rect 589150 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 589770 622574
rect 589150 586894 589770 622338
rect 589150 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 589770 586894
rect 589150 586574 589770 586658
rect 589150 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 589770 586574
rect 589150 550894 589770 586338
rect 589150 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 589770 550894
rect 589150 550574 589770 550658
rect 589150 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 589770 550574
rect 589150 514894 589770 550338
rect 589150 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 589770 514894
rect 589150 514574 589770 514658
rect 589150 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 589770 514574
rect 589150 478894 589770 514338
rect 589150 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 589770 478894
rect 589150 478574 589770 478658
rect 589150 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 589770 478574
rect 589150 442894 589770 478338
rect 589150 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 589770 442894
rect 589150 442574 589770 442658
rect 589150 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 589770 442574
rect 589150 406894 589770 442338
rect 589150 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 589770 406894
rect 589150 406574 589770 406658
rect 589150 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 589770 406574
rect 589150 370894 589770 406338
rect 589150 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 589770 370894
rect 589150 370574 589770 370658
rect 589150 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 589770 370574
rect 589150 334894 589770 370338
rect 589150 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 589770 334894
rect 589150 334574 589770 334658
rect 589150 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 589770 334574
rect 589150 298894 589770 334338
rect 589150 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 589770 298894
rect 589150 298574 589770 298658
rect 589150 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 589770 298574
rect 589150 262894 589770 298338
rect 589150 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 589770 262894
rect 589150 262574 589770 262658
rect 589150 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 589770 262574
rect 589150 226894 589770 262338
rect 589150 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 589770 226894
rect 589150 226574 589770 226658
rect 589150 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 589770 226574
rect 589150 190894 589770 226338
rect 589150 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 589770 190894
rect 589150 190574 589770 190658
rect 589150 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 589770 190574
rect 589150 154894 589770 190338
rect 589150 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 589770 154894
rect 589150 154574 589770 154658
rect 589150 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 589770 154574
rect 589150 118894 589770 154338
rect 589150 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 589770 118894
rect 589150 118574 589770 118658
rect 589150 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 589770 118574
rect 589150 82894 589770 118338
rect 589150 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 589770 82894
rect 589150 82574 589770 82658
rect 589150 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 589770 82574
rect 589150 46894 589770 82338
rect 589150 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 589770 46894
rect 589150 46574 589770 46658
rect 589150 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 589770 46574
rect 589150 10894 589770 46338
rect 589150 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 589770 10894
rect 589150 10574 589770 10658
rect 589150 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 589770 10574
rect 589150 -4186 589770 10338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect 590110 676574 590730 676658
rect 590110 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect 590110 640894 590730 676338
rect 590110 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect 590110 640574 590730 640658
rect 590110 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect 590110 604894 590730 640338
rect 590110 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect 590110 604574 590730 604658
rect 590110 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect 590110 568894 590730 604338
rect 590110 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect 590110 568574 590730 568658
rect 590110 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect 590110 532894 590730 568338
rect 590110 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect 590110 532574 590730 532658
rect 590110 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect 590110 496894 590730 532338
rect 590110 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect 590110 496574 590730 496658
rect 590110 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect 590110 460894 590730 496338
rect 590110 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect 590110 460574 590730 460658
rect 590110 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect 590110 424894 590730 460338
rect 590110 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 590110 424574 590730 424658
rect 590110 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 590110 388894 590730 424338
rect 590110 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 590110 388574 590730 388658
rect 590110 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 590110 352894 590730 388338
rect 590110 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 590110 352574 590730 352658
rect 590110 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 590110 316894 590730 352338
rect 590110 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 590110 316574 590730 316658
rect 590110 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 590110 280894 590730 316338
rect 590110 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 590110 280574 590730 280658
rect 590110 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 590110 244894 590730 280338
rect 590110 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 590110 244574 590730 244658
rect 590110 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 590110 208894 590730 244338
rect 590110 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 590110 208574 590730 208658
rect 590110 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 590110 172894 590730 208338
rect 590110 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 590110 172574 590730 172658
rect 590110 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 590110 136894 590730 172338
rect 590110 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 590110 136574 590730 136658
rect 590110 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 590110 100894 590730 136338
rect 590110 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 590110 100574 590730 100658
rect 590110 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 590110 64894 590730 100338
rect 590110 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 590110 64574 590730 64658
rect 590110 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 590110 28894 590730 64338
rect 590110 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect 590110 28574 590730 28658
rect 590110 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect 590110 -5146 590730 28338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 591690 698614
rect 591070 698294 591690 698378
rect 591070 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 591690 698294
rect 591070 662614 591690 698058
rect 591070 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 591690 662614
rect 591070 662294 591690 662378
rect 591070 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 591690 662294
rect 591070 626614 591690 662058
rect 591070 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 591690 626614
rect 591070 626294 591690 626378
rect 591070 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 591690 626294
rect 591070 590614 591690 626058
rect 591070 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 591690 590614
rect 591070 590294 591690 590378
rect 591070 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 591690 590294
rect 591070 554614 591690 590058
rect 591070 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 591690 554614
rect 591070 554294 591690 554378
rect 591070 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 591690 554294
rect 591070 518614 591690 554058
rect 591070 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 591690 518614
rect 591070 518294 591690 518378
rect 591070 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 591690 518294
rect 591070 482614 591690 518058
rect 591070 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 591690 482614
rect 591070 482294 591690 482378
rect 591070 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 591690 482294
rect 591070 446614 591690 482058
rect 591070 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 591690 446614
rect 591070 446294 591690 446378
rect 591070 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 591690 446294
rect 591070 410614 591690 446058
rect 591070 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 591690 410614
rect 591070 410294 591690 410378
rect 591070 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 591690 410294
rect 591070 374614 591690 410058
rect 591070 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 591690 374614
rect 591070 374294 591690 374378
rect 591070 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 591690 374294
rect 591070 338614 591690 374058
rect 591070 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 591690 338614
rect 591070 338294 591690 338378
rect 591070 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 591690 338294
rect 591070 302614 591690 338058
rect 591070 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 591690 302614
rect 591070 302294 591690 302378
rect 591070 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 591690 302294
rect 591070 266614 591690 302058
rect 591070 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 591690 266614
rect 591070 266294 591690 266378
rect 591070 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 591690 266294
rect 591070 230614 591690 266058
rect 591070 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 591690 230614
rect 591070 230294 591690 230378
rect 591070 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 591690 230294
rect 591070 194614 591690 230058
rect 591070 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 591690 194614
rect 591070 194294 591690 194378
rect 591070 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 591690 194294
rect 591070 158614 591690 194058
rect 591070 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 591690 158614
rect 591070 158294 591690 158378
rect 591070 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 591690 158294
rect 591070 122614 591690 158058
rect 591070 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 591690 122614
rect 591070 122294 591690 122378
rect 591070 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 591690 122294
rect 591070 86614 591690 122058
rect 591070 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 591690 86614
rect 591070 86294 591690 86378
rect 591070 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 591690 86294
rect 591070 50614 591690 86058
rect 591070 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 591690 50614
rect 591070 50294 591690 50378
rect 591070 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 591690 50294
rect 591070 14614 591690 50058
rect 591070 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 591690 14614
rect 591070 14294 591690 14378
rect 591070 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 591690 14294
rect 591070 -6106 591690 14058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect 592030 680294 592650 680378
rect 592030 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect 592030 644614 592650 680058
rect 592030 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect 592030 644294 592650 644378
rect 592030 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect 592030 608614 592650 644058
rect 592030 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect 592030 608294 592650 608378
rect 592030 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect 592030 572614 592650 608058
rect 592030 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect 592030 572294 592650 572378
rect 592030 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect 592030 536614 592650 572058
rect 592030 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect 592030 536294 592650 536378
rect 592030 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect 592030 500614 592650 536058
rect 592030 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect 592030 500294 592650 500378
rect 592030 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect 592030 464614 592650 500058
rect 592030 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect 592030 464294 592650 464378
rect 592030 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect 592030 428614 592650 464058
rect 592030 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 592030 428294 592650 428378
rect 592030 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 592030 392614 592650 428058
rect 592030 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 592030 392294 592650 392378
rect 592030 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 592030 356614 592650 392058
rect 592030 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 592030 356294 592650 356378
rect 592030 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 592030 320614 592650 356058
rect 592030 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 592030 320294 592650 320378
rect 592030 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 592030 284614 592650 320058
rect 592030 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 592030 284294 592650 284378
rect 592030 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 592030 248614 592650 284058
rect 592030 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 592030 248294 592650 248378
rect 592030 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 592030 212614 592650 248058
rect 592030 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 592030 212294 592650 212378
rect 592030 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 592030 176614 592650 212058
rect 592030 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 592030 176294 592650 176378
rect 592030 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 592030 140614 592650 176058
rect 592030 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 592030 140294 592650 140378
rect 592030 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 592030 104614 592650 140058
rect 592030 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 592030 104294 592650 104378
rect 592030 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 592030 68614 592650 104058
rect 592030 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 592030 68294 592650 68378
rect 592030 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 592030 32614 592650 68058
rect 592030 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect 592030 32294 592650 32378
rect 592030 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect 570954 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 571574 -7066
rect 570954 -7386 571574 -7302
rect 570954 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 571574 -7386
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 680378 -8458 680614
rect -8374 680378 -8138 680614
rect -8694 680058 -8458 680294
rect -8374 680058 -8138 680294
rect -8694 644378 -8458 644614
rect -8374 644378 -8138 644614
rect -8694 644058 -8458 644294
rect -8374 644058 -8138 644294
rect -8694 608378 -8458 608614
rect -8374 608378 -8138 608614
rect -8694 608058 -8458 608294
rect -8374 608058 -8138 608294
rect -8694 572378 -8458 572614
rect -8374 572378 -8138 572614
rect -8694 572058 -8458 572294
rect -8374 572058 -8138 572294
rect -8694 536378 -8458 536614
rect -8374 536378 -8138 536614
rect -8694 536058 -8458 536294
rect -8374 536058 -8138 536294
rect -8694 500378 -8458 500614
rect -8374 500378 -8138 500614
rect -8694 500058 -8458 500294
rect -8374 500058 -8138 500294
rect -8694 464378 -8458 464614
rect -8374 464378 -8138 464614
rect -8694 464058 -8458 464294
rect -8374 464058 -8138 464294
rect -8694 428378 -8458 428614
rect -8374 428378 -8138 428614
rect -8694 428058 -8458 428294
rect -8374 428058 -8138 428294
rect -8694 392378 -8458 392614
rect -8374 392378 -8138 392614
rect -8694 392058 -8458 392294
rect -8374 392058 -8138 392294
rect -8694 356378 -8458 356614
rect -8374 356378 -8138 356614
rect -8694 356058 -8458 356294
rect -8374 356058 -8138 356294
rect -8694 320378 -8458 320614
rect -8374 320378 -8138 320614
rect -8694 320058 -8458 320294
rect -8374 320058 -8138 320294
rect -8694 284378 -8458 284614
rect -8374 284378 -8138 284614
rect -8694 284058 -8458 284294
rect -8374 284058 -8138 284294
rect -8694 248378 -8458 248614
rect -8374 248378 -8138 248614
rect -8694 248058 -8458 248294
rect -8374 248058 -8138 248294
rect -8694 212378 -8458 212614
rect -8374 212378 -8138 212614
rect -8694 212058 -8458 212294
rect -8374 212058 -8138 212294
rect -8694 176378 -8458 176614
rect -8374 176378 -8138 176614
rect -8694 176058 -8458 176294
rect -8374 176058 -8138 176294
rect -8694 140378 -8458 140614
rect -8374 140378 -8138 140614
rect -8694 140058 -8458 140294
rect -8374 140058 -8138 140294
rect -8694 104378 -8458 104614
rect -8374 104378 -8138 104614
rect -8694 104058 -8458 104294
rect -8374 104058 -8138 104294
rect -8694 68378 -8458 68614
rect -8374 68378 -8138 68614
rect -8694 68058 -8458 68294
rect -8374 68058 -8138 68294
rect -8694 32378 -8458 32614
rect -8374 32378 -8138 32614
rect -8694 32058 -8458 32294
rect -8374 32058 -8138 32294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12986 710362 13222 710598
rect 13306 710362 13542 710598
rect 12986 710042 13222 710278
rect 13306 710042 13542 710278
rect -7734 698378 -7498 698614
rect -7414 698378 -7178 698614
rect -7734 698058 -7498 698294
rect -7414 698058 -7178 698294
rect -7734 662378 -7498 662614
rect -7414 662378 -7178 662614
rect -7734 662058 -7498 662294
rect -7414 662058 -7178 662294
rect -7734 626378 -7498 626614
rect -7414 626378 -7178 626614
rect -7734 626058 -7498 626294
rect -7414 626058 -7178 626294
rect -7734 590378 -7498 590614
rect -7414 590378 -7178 590614
rect -7734 590058 -7498 590294
rect -7414 590058 -7178 590294
rect -7734 554378 -7498 554614
rect -7414 554378 -7178 554614
rect -7734 554058 -7498 554294
rect -7414 554058 -7178 554294
rect -7734 518378 -7498 518614
rect -7414 518378 -7178 518614
rect -7734 518058 -7498 518294
rect -7414 518058 -7178 518294
rect -7734 482378 -7498 482614
rect -7414 482378 -7178 482614
rect -7734 482058 -7498 482294
rect -7414 482058 -7178 482294
rect -7734 446378 -7498 446614
rect -7414 446378 -7178 446614
rect -7734 446058 -7498 446294
rect -7414 446058 -7178 446294
rect -7734 410378 -7498 410614
rect -7414 410378 -7178 410614
rect -7734 410058 -7498 410294
rect -7414 410058 -7178 410294
rect -7734 374378 -7498 374614
rect -7414 374378 -7178 374614
rect -7734 374058 -7498 374294
rect -7414 374058 -7178 374294
rect -7734 338378 -7498 338614
rect -7414 338378 -7178 338614
rect -7734 338058 -7498 338294
rect -7414 338058 -7178 338294
rect -7734 302378 -7498 302614
rect -7414 302378 -7178 302614
rect -7734 302058 -7498 302294
rect -7414 302058 -7178 302294
rect -7734 266378 -7498 266614
rect -7414 266378 -7178 266614
rect -7734 266058 -7498 266294
rect -7414 266058 -7178 266294
rect -7734 230378 -7498 230614
rect -7414 230378 -7178 230614
rect -7734 230058 -7498 230294
rect -7414 230058 -7178 230294
rect -7734 194378 -7498 194614
rect -7414 194378 -7178 194614
rect -7734 194058 -7498 194294
rect -7414 194058 -7178 194294
rect -7734 158378 -7498 158614
rect -7414 158378 -7178 158614
rect -7734 158058 -7498 158294
rect -7414 158058 -7178 158294
rect -7734 122378 -7498 122614
rect -7414 122378 -7178 122614
rect -7734 122058 -7498 122294
rect -7414 122058 -7178 122294
rect -7734 86378 -7498 86614
rect -7414 86378 -7178 86614
rect -7734 86058 -7498 86294
rect -7414 86058 -7178 86294
rect -7734 50378 -7498 50614
rect -7414 50378 -7178 50614
rect -7734 50058 -7498 50294
rect -7414 50058 -7178 50294
rect -7734 14378 -7498 14614
rect -7414 14378 -7178 14614
rect -7734 14058 -7498 14294
rect -7414 14058 -7178 14294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 676658 -6538 676894
rect -6454 676658 -6218 676894
rect -6774 676338 -6538 676574
rect -6454 676338 -6218 676574
rect -6774 640658 -6538 640894
rect -6454 640658 -6218 640894
rect -6774 640338 -6538 640574
rect -6454 640338 -6218 640574
rect -6774 604658 -6538 604894
rect -6454 604658 -6218 604894
rect -6774 604338 -6538 604574
rect -6454 604338 -6218 604574
rect -6774 568658 -6538 568894
rect -6454 568658 -6218 568894
rect -6774 568338 -6538 568574
rect -6454 568338 -6218 568574
rect -6774 532658 -6538 532894
rect -6454 532658 -6218 532894
rect -6774 532338 -6538 532574
rect -6454 532338 -6218 532574
rect -6774 496658 -6538 496894
rect -6454 496658 -6218 496894
rect -6774 496338 -6538 496574
rect -6454 496338 -6218 496574
rect -6774 460658 -6538 460894
rect -6454 460658 -6218 460894
rect -6774 460338 -6538 460574
rect -6454 460338 -6218 460574
rect -6774 424658 -6538 424894
rect -6454 424658 -6218 424894
rect -6774 424338 -6538 424574
rect -6454 424338 -6218 424574
rect -6774 388658 -6538 388894
rect -6454 388658 -6218 388894
rect -6774 388338 -6538 388574
rect -6454 388338 -6218 388574
rect -6774 352658 -6538 352894
rect -6454 352658 -6218 352894
rect -6774 352338 -6538 352574
rect -6454 352338 -6218 352574
rect -6774 316658 -6538 316894
rect -6454 316658 -6218 316894
rect -6774 316338 -6538 316574
rect -6454 316338 -6218 316574
rect -6774 280658 -6538 280894
rect -6454 280658 -6218 280894
rect -6774 280338 -6538 280574
rect -6454 280338 -6218 280574
rect -6774 244658 -6538 244894
rect -6454 244658 -6218 244894
rect -6774 244338 -6538 244574
rect -6454 244338 -6218 244574
rect -6774 208658 -6538 208894
rect -6454 208658 -6218 208894
rect -6774 208338 -6538 208574
rect -6454 208338 -6218 208574
rect -6774 172658 -6538 172894
rect -6454 172658 -6218 172894
rect -6774 172338 -6538 172574
rect -6454 172338 -6218 172574
rect -6774 136658 -6538 136894
rect -6454 136658 -6218 136894
rect -6774 136338 -6538 136574
rect -6454 136338 -6218 136574
rect -6774 100658 -6538 100894
rect -6454 100658 -6218 100894
rect -6774 100338 -6538 100574
rect -6454 100338 -6218 100574
rect -6774 64658 -6538 64894
rect -6454 64658 -6218 64894
rect -6774 64338 -6538 64574
rect -6454 64338 -6218 64574
rect -6774 28658 -6538 28894
rect -6454 28658 -6218 28894
rect -6774 28338 -6538 28574
rect -6454 28338 -6218 28574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 9266 708442 9502 708678
rect 9586 708442 9822 708678
rect 9266 708122 9502 708358
rect 9586 708122 9822 708358
rect -5814 694658 -5578 694894
rect -5494 694658 -5258 694894
rect -5814 694338 -5578 694574
rect -5494 694338 -5258 694574
rect -5814 658658 -5578 658894
rect -5494 658658 -5258 658894
rect -5814 658338 -5578 658574
rect -5494 658338 -5258 658574
rect -5814 622658 -5578 622894
rect -5494 622658 -5258 622894
rect -5814 622338 -5578 622574
rect -5494 622338 -5258 622574
rect -5814 586658 -5578 586894
rect -5494 586658 -5258 586894
rect -5814 586338 -5578 586574
rect -5494 586338 -5258 586574
rect -5814 550658 -5578 550894
rect -5494 550658 -5258 550894
rect -5814 550338 -5578 550574
rect -5494 550338 -5258 550574
rect -5814 514658 -5578 514894
rect -5494 514658 -5258 514894
rect -5814 514338 -5578 514574
rect -5494 514338 -5258 514574
rect -5814 478658 -5578 478894
rect -5494 478658 -5258 478894
rect -5814 478338 -5578 478574
rect -5494 478338 -5258 478574
rect -5814 442658 -5578 442894
rect -5494 442658 -5258 442894
rect -5814 442338 -5578 442574
rect -5494 442338 -5258 442574
rect -5814 406658 -5578 406894
rect -5494 406658 -5258 406894
rect -5814 406338 -5578 406574
rect -5494 406338 -5258 406574
rect -5814 370658 -5578 370894
rect -5494 370658 -5258 370894
rect -5814 370338 -5578 370574
rect -5494 370338 -5258 370574
rect -5814 334658 -5578 334894
rect -5494 334658 -5258 334894
rect -5814 334338 -5578 334574
rect -5494 334338 -5258 334574
rect -5814 298658 -5578 298894
rect -5494 298658 -5258 298894
rect -5814 298338 -5578 298574
rect -5494 298338 -5258 298574
rect -5814 262658 -5578 262894
rect -5494 262658 -5258 262894
rect -5814 262338 -5578 262574
rect -5494 262338 -5258 262574
rect -5814 226658 -5578 226894
rect -5494 226658 -5258 226894
rect -5814 226338 -5578 226574
rect -5494 226338 -5258 226574
rect -5814 190658 -5578 190894
rect -5494 190658 -5258 190894
rect -5814 190338 -5578 190574
rect -5494 190338 -5258 190574
rect -5814 154658 -5578 154894
rect -5494 154658 -5258 154894
rect -5814 154338 -5578 154574
rect -5494 154338 -5258 154574
rect -5814 118658 -5578 118894
rect -5494 118658 -5258 118894
rect -5814 118338 -5578 118574
rect -5494 118338 -5258 118574
rect -5814 82658 -5578 82894
rect -5494 82658 -5258 82894
rect -5814 82338 -5578 82574
rect -5494 82338 -5258 82574
rect -5814 46658 -5578 46894
rect -5494 46658 -5258 46894
rect -5814 46338 -5578 46574
rect -5494 46338 -5258 46574
rect -5814 10658 -5578 10894
rect -5494 10658 -5258 10894
rect -5814 10338 -5578 10574
rect -5494 10338 -5258 10574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 672938 -4618 673174
rect -4534 672938 -4298 673174
rect -4854 672618 -4618 672854
rect -4534 672618 -4298 672854
rect -4854 636938 -4618 637174
rect -4534 636938 -4298 637174
rect -4854 636618 -4618 636854
rect -4534 636618 -4298 636854
rect -4854 600938 -4618 601174
rect -4534 600938 -4298 601174
rect -4854 600618 -4618 600854
rect -4534 600618 -4298 600854
rect -4854 564938 -4618 565174
rect -4534 564938 -4298 565174
rect -4854 564618 -4618 564854
rect -4534 564618 -4298 564854
rect -4854 528938 -4618 529174
rect -4534 528938 -4298 529174
rect -4854 528618 -4618 528854
rect -4534 528618 -4298 528854
rect -4854 492938 -4618 493174
rect -4534 492938 -4298 493174
rect -4854 492618 -4618 492854
rect -4534 492618 -4298 492854
rect -4854 456938 -4618 457174
rect -4534 456938 -4298 457174
rect -4854 456618 -4618 456854
rect -4534 456618 -4298 456854
rect -4854 420938 -4618 421174
rect -4534 420938 -4298 421174
rect -4854 420618 -4618 420854
rect -4534 420618 -4298 420854
rect -4854 384938 -4618 385174
rect -4534 384938 -4298 385174
rect -4854 384618 -4618 384854
rect -4534 384618 -4298 384854
rect -4854 348938 -4618 349174
rect -4534 348938 -4298 349174
rect -4854 348618 -4618 348854
rect -4534 348618 -4298 348854
rect -4854 312938 -4618 313174
rect -4534 312938 -4298 313174
rect -4854 312618 -4618 312854
rect -4534 312618 -4298 312854
rect -4854 276938 -4618 277174
rect -4534 276938 -4298 277174
rect -4854 276618 -4618 276854
rect -4534 276618 -4298 276854
rect -4854 240938 -4618 241174
rect -4534 240938 -4298 241174
rect -4854 240618 -4618 240854
rect -4534 240618 -4298 240854
rect -4854 204938 -4618 205174
rect -4534 204938 -4298 205174
rect -4854 204618 -4618 204854
rect -4534 204618 -4298 204854
rect -4854 168938 -4618 169174
rect -4534 168938 -4298 169174
rect -4854 168618 -4618 168854
rect -4534 168618 -4298 168854
rect -4854 132938 -4618 133174
rect -4534 132938 -4298 133174
rect -4854 132618 -4618 132854
rect -4534 132618 -4298 132854
rect -4854 96938 -4618 97174
rect -4534 96938 -4298 97174
rect -4854 96618 -4618 96854
rect -4534 96618 -4298 96854
rect -4854 60938 -4618 61174
rect -4534 60938 -4298 61174
rect -4854 60618 -4618 60854
rect -4534 60618 -4298 60854
rect -4854 24938 -4618 25174
rect -4534 24938 -4298 25174
rect -4854 24618 -4618 24854
rect -4534 24618 -4298 24854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 5546 706522 5782 706758
rect 5866 706522 6102 706758
rect 5546 706202 5782 706438
rect 5866 706202 6102 706438
rect -3894 690938 -3658 691174
rect -3574 690938 -3338 691174
rect -3894 690618 -3658 690854
rect -3574 690618 -3338 690854
rect -3894 654938 -3658 655174
rect -3574 654938 -3338 655174
rect -3894 654618 -3658 654854
rect -3574 654618 -3338 654854
rect -3894 618938 -3658 619174
rect -3574 618938 -3338 619174
rect -3894 618618 -3658 618854
rect -3574 618618 -3338 618854
rect -3894 582938 -3658 583174
rect -3574 582938 -3338 583174
rect -3894 582618 -3658 582854
rect -3574 582618 -3338 582854
rect -3894 546938 -3658 547174
rect -3574 546938 -3338 547174
rect -3894 546618 -3658 546854
rect -3574 546618 -3338 546854
rect -3894 510938 -3658 511174
rect -3574 510938 -3338 511174
rect -3894 510618 -3658 510854
rect -3574 510618 -3338 510854
rect -3894 474938 -3658 475174
rect -3574 474938 -3338 475174
rect -3894 474618 -3658 474854
rect -3574 474618 -3338 474854
rect -3894 438938 -3658 439174
rect -3574 438938 -3338 439174
rect -3894 438618 -3658 438854
rect -3574 438618 -3338 438854
rect -3894 402938 -3658 403174
rect -3574 402938 -3338 403174
rect -3894 402618 -3658 402854
rect -3574 402618 -3338 402854
rect -3894 366938 -3658 367174
rect -3574 366938 -3338 367174
rect -3894 366618 -3658 366854
rect -3574 366618 -3338 366854
rect -3894 330938 -3658 331174
rect -3574 330938 -3338 331174
rect -3894 330618 -3658 330854
rect -3574 330618 -3338 330854
rect -3894 294938 -3658 295174
rect -3574 294938 -3338 295174
rect -3894 294618 -3658 294854
rect -3574 294618 -3338 294854
rect -3894 258938 -3658 259174
rect -3574 258938 -3338 259174
rect -3894 258618 -3658 258854
rect -3574 258618 -3338 258854
rect -3894 222938 -3658 223174
rect -3574 222938 -3338 223174
rect -3894 222618 -3658 222854
rect -3574 222618 -3338 222854
rect -3894 186938 -3658 187174
rect -3574 186938 -3338 187174
rect -3894 186618 -3658 186854
rect -3574 186618 -3338 186854
rect -3894 150938 -3658 151174
rect -3574 150938 -3338 151174
rect -3894 150618 -3658 150854
rect -3574 150618 -3338 150854
rect -3894 114938 -3658 115174
rect -3574 114938 -3338 115174
rect -3894 114618 -3658 114854
rect -3574 114618 -3338 114854
rect -3894 78938 -3658 79174
rect -3574 78938 -3338 79174
rect -3894 78618 -3658 78854
rect -3574 78618 -3338 78854
rect -3894 42938 -3658 43174
rect -3574 42938 -3338 43174
rect -3894 42618 -3658 42854
rect -3574 42618 -3338 42854
rect -3894 6938 -3658 7174
rect -3574 6938 -3338 7174
rect -3894 6618 -3658 6854
rect -3574 6618 -3338 6854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 30986 711322 31222 711558
rect 31306 711322 31542 711558
rect 30986 711002 31222 711238
rect 31306 711002 31542 711238
rect 27266 709402 27502 709638
rect 27586 709402 27822 709638
rect 27266 709082 27502 709318
rect 27586 709082 27822 709318
rect 23546 707482 23782 707718
rect 23866 707482 24102 707718
rect 23546 707162 23782 707398
rect 23866 707162 24102 707398
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 48986 710362 49222 710598
rect 49306 710362 49542 710598
rect 48986 710042 49222 710278
rect 49306 710042 49542 710278
rect 45266 708442 45502 708678
rect 45586 708442 45822 708678
rect 45266 708122 45502 708358
rect 45586 708122 45822 708358
rect 41546 706522 41782 706758
rect 41866 706522 42102 706758
rect 41546 706202 41782 706438
rect 41866 706202 42102 706438
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 66986 711322 67222 711558
rect 67306 711322 67542 711558
rect 66986 711002 67222 711238
rect 67306 711002 67542 711238
rect 63266 709402 63502 709638
rect 63586 709402 63822 709638
rect 63266 709082 63502 709318
rect 63586 709082 63822 709318
rect 59546 707482 59782 707718
rect 59866 707482 60102 707718
rect 59546 707162 59782 707398
rect 59866 707162 60102 707398
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 84986 710362 85222 710598
rect 85306 710362 85542 710598
rect 84986 710042 85222 710278
rect 85306 710042 85542 710278
rect 81266 708442 81502 708678
rect 81586 708442 81822 708678
rect 81266 708122 81502 708358
rect 81586 708122 81822 708358
rect 77546 706522 77782 706758
rect 77866 706522 78102 706758
rect 77546 706202 77782 706438
rect 77866 706202 78102 706438
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 102986 711322 103222 711558
rect 103306 711322 103542 711558
rect 102986 711002 103222 711238
rect 103306 711002 103542 711238
rect 99266 709402 99502 709638
rect 99586 709402 99822 709638
rect 99266 709082 99502 709318
rect 99586 709082 99822 709318
rect 95546 707482 95782 707718
rect 95866 707482 96102 707718
rect 95546 707162 95782 707398
rect 95866 707162 96102 707398
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 120986 710362 121222 710598
rect 121306 710362 121542 710598
rect 120986 710042 121222 710278
rect 121306 710042 121542 710278
rect 117266 708442 117502 708678
rect 117586 708442 117822 708678
rect 117266 708122 117502 708358
rect 117586 708122 117822 708358
rect 113546 706522 113782 706758
rect 113866 706522 114102 706758
rect 113546 706202 113782 706438
rect 113866 706202 114102 706438
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 138986 711322 139222 711558
rect 139306 711322 139542 711558
rect 138986 711002 139222 711238
rect 139306 711002 139542 711238
rect 135266 709402 135502 709638
rect 135586 709402 135822 709638
rect 135266 709082 135502 709318
rect 135586 709082 135822 709318
rect 131546 707482 131782 707718
rect 131866 707482 132102 707718
rect 131546 707162 131782 707398
rect 131866 707162 132102 707398
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 156986 710362 157222 710598
rect 157306 710362 157542 710598
rect 156986 710042 157222 710278
rect 157306 710042 157542 710278
rect 153266 708442 153502 708678
rect 153586 708442 153822 708678
rect 153266 708122 153502 708358
rect 153586 708122 153822 708358
rect 149546 706522 149782 706758
rect 149866 706522 150102 706758
rect 149546 706202 149782 706438
rect 149866 706202 150102 706438
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 174986 711322 175222 711558
rect 175306 711322 175542 711558
rect 174986 711002 175222 711238
rect 175306 711002 175542 711238
rect 171266 709402 171502 709638
rect 171586 709402 171822 709638
rect 171266 709082 171502 709318
rect 171586 709082 171822 709318
rect 167546 707482 167782 707718
rect 167866 707482 168102 707718
rect 167546 707162 167782 707398
rect 167866 707162 168102 707398
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 192986 710362 193222 710598
rect 193306 710362 193542 710598
rect 192986 710042 193222 710278
rect 193306 710042 193542 710278
rect 189266 708442 189502 708678
rect 189586 708442 189822 708678
rect 189266 708122 189502 708358
rect 189586 708122 189822 708358
rect 185546 706522 185782 706758
rect 185866 706522 186102 706758
rect 185546 706202 185782 706438
rect 185866 706202 186102 706438
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 210986 711322 211222 711558
rect 211306 711322 211542 711558
rect 210986 711002 211222 711238
rect 211306 711002 211542 711238
rect 207266 709402 207502 709638
rect 207586 709402 207822 709638
rect 207266 709082 207502 709318
rect 207586 709082 207822 709318
rect 203546 707482 203782 707718
rect 203866 707482 204102 707718
rect 203546 707162 203782 707398
rect 203866 707162 204102 707398
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 228986 710362 229222 710598
rect 229306 710362 229542 710598
rect 228986 710042 229222 710278
rect 229306 710042 229542 710278
rect 225266 708442 225502 708678
rect 225586 708442 225822 708678
rect 225266 708122 225502 708358
rect 225586 708122 225822 708358
rect 221546 706522 221782 706758
rect 221866 706522 222102 706758
rect 221546 706202 221782 706438
rect 221866 706202 222102 706438
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 246986 711322 247222 711558
rect 247306 711322 247542 711558
rect 246986 711002 247222 711238
rect 247306 711002 247542 711238
rect 243266 709402 243502 709638
rect 243586 709402 243822 709638
rect 243266 709082 243502 709318
rect 243586 709082 243822 709318
rect 239546 707482 239782 707718
rect 239866 707482 240102 707718
rect 239546 707162 239782 707398
rect 239866 707162 240102 707398
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 264986 710362 265222 710598
rect 265306 710362 265542 710598
rect 264986 710042 265222 710278
rect 265306 710042 265542 710278
rect 261266 708442 261502 708678
rect 261586 708442 261822 708678
rect 261266 708122 261502 708358
rect 261586 708122 261822 708358
rect 257546 706522 257782 706758
rect 257866 706522 258102 706758
rect 257546 706202 257782 706438
rect 257866 706202 258102 706438
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 282986 711322 283222 711558
rect 283306 711322 283542 711558
rect 282986 711002 283222 711238
rect 283306 711002 283542 711238
rect 279266 709402 279502 709638
rect 279586 709402 279822 709638
rect 279266 709082 279502 709318
rect 279586 709082 279822 709318
rect 275546 707482 275782 707718
rect 275866 707482 276102 707718
rect 275546 707162 275782 707398
rect 275866 707162 276102 707398
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 300986 710362 301222 710598
rect 301306 710362 301542 710598
rect 300986 710042 301222 710278
rect 301306 710042 301542 710278
rect 297266 708442 297502 708678
rect 297586 708442 297822 708678
rect 297266 708122 297502 708358
rect 297586 708122 297822 708358
rect 293546 706522 293782 706758
rect 293866 706522 294102 706758
rect 293546 706202 293782 706438
rect 293866 706202 294102 706438
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 318986 711322 319222 711558
rect 319306 711322 319542 711558
rect 318986 711002 319222 711238
rect 319306 711002 319542 711238
rect 315266 709402 315502 709638
rect 315586 709402 315822 709638
rect 315266 709082 315502 709318
rect 315586 709082 315822 709318
rect 311546 707482 311782 707718
rect 311866 707482 312102 707718
rect 311546 707162 311782 707398
rect 311866 707162 312102 707398
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 336986 710362 337222 710598
rect 337306 710362 337542 710598
rect 336986 710042 337222 710278
rect 337306 710042 337542 710278
rect 333266 708442 333502 708678
rect 333586 708442 333822 708678
rect 333266 708122 333502 708358
rect 333586 708122 333822 708358
rect 329546 706522 329782 706758
rect 329866 706522 330102 706758
rect 329546 706202 329782 706438
rect 329866 706202 330102 706438
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 354986 711322 355222 711558
rect 355306 711322 355542 711558
rect 354986 711002 355222 711238
rect 355306 711002 355542 711238
rect 351266 709402 351502 709638
rect 351586 709402 351822 709638
rect 351266 709082 351502 709318
rect 351586 709082 351822 709318
rect 347546 707482 347782 707718
rect 347866 707482 348102 707718
rect 347546 707162 347782 707398
rect 347866 707162 348102 707398
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 372986 710362 373222 710598
rect 373306 710362 373542 710598
rect 372986 710042 373222 710278
rect 373306 710042 373542 710278
rect 369266 708442 369502 708678
rect 369586 708442 369822 708678
rect 369266 708122 369502 708358
rect 369586 708122 369822 708358
rect 365546 706522 365782 706758
rect 365866 706522 366102 706758
rect 365546 706202 365782 706438
rect 365866 706202 366102 706438
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 390986 711322 391222 711558
rect 391306 711322 391542 711558
rect 390986 711002 391222 711238
rect 391306 711002 391542 711238
rect 387266 709402 387502 709638
rect 387586 709402 387822 709638
rect 387266 709082 387502 709318
rect 387586 709082 387822 709318
rect 383546 707482 383782 707718
rect 383866 707482 384102 707718
rect 383546 707162 383782 707398
rect 383866 707162 384102 707398
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 408986 710362 409222 710598
rect 409306 710362 409542 710598
rect 408986 710042 409222 710278
rect 409306 710042 409542 710278
rect 405266 708442 405502 708678
rect 405586 708442 405822 708678
rect 405266 708122 405502 708358
rect 405586 708122 405822 708358
rect 401546 706522 401782 706758
rect 401866 706522 402102 706758
rect 401546 706202 401782 706438
rect 401866 706202 402102 706438
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 426986 711322 427222 711558
rect 427306 711322 427542 711558
rect 426986 711002 427222 711238
rect 427306 711002 427542 711238
rect 423266 709402 423502 709638
rect 423586 709402 423822 709638
rect 423266 709082 423502 709318
rect 423586 709082 423822 709318
rect 419546 707482 419782 707718
rect 419866 707482 420102 707718
rect 419546 707162 419782 707398
rect 419866 707162 420102 707398
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 444986 710362 445222 710598
rect 445306 710362 445542 710598
rect 444986 710042 445222 710278
rect 445306 710042 445542 710278
rect 441266 708442 441502 708678
rect 441586 708442 441822 708678
rect 441266 708122 441502 708358
rect 441586 708122 441822 708358
rect 437546 706522 437782 706758
rect 437866 706522 438102 706758
rect 437546 706202 437782 706438
rect 437866 706202 438102 706438
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 462986 711322 463222 711558
rect 463306 711322 463542 711558
rect 462986 711002 463222 711238
rect 463306 711002 463542 711238
rect 459266 709402 459502 709638
rect 459586 709402 459822 709638
rect 459266 709082 459502 709318
rect 459586 709082 459822 709318
rect 455546 707482 455782 707718
rect 455866 707482 456102 707718
rect 455546 707162 455782 707398
rect 455866 707162 456102 707398
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 480986 710362 481222 710598
rect 481306 710362 481542 710598
rect 480986 710042 481222 710278
rect 481306 710042 481542 710278
rect 477266 708442 477502 708678
rect 477586 708442 477822 708678
rect 477266 708122 477502 708358
rect 477586 708122 477822 708358
rect 473546 706522 473782 706758
rect 473866 706522 474102 706758
rect 473546 706202 473782 706438
rect 473866 706202 474102 706438
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 498986 711322 499222 711558
rect 499306 711322 499542 711558
rect 498986 711002 499222 711238
rect 499306 711002 499542 711238
rect 495266 709402 495502 709638
rect 495586 709402 495822 709638
rect 495266 709082 495502 709318
rect 495586 709082 495822 709318
rect 491546 707482 491782 707718
rect 491866 707482 492102 707718
rect 491546 707162 491782 707398
rect 491866 707162 492102 707398
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 516986 710362 517222 710598
rect 517306 710362 517542 710598
rect 516986 710042 517222 710278
rect 517306 710042 517542 710278
rect 513266 708442 513502 708678
rect 513586 708442 513822 708678
rect 513266 708122 513502 708358
rect 513586 708122 513822 708358
rect 509546 706522 509782 706758
rect 509866 706522 510102 706758
rect 509546 706202 509782 706438
rect 509866 706202 510102 706438
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 534986 711322 535222 711558
rect 535306 711322 535542 711558
rect 534986 711002 535222 711238
rect 535306 711002 535542 711238
rect 531266 709402 531502 709638
rect 531586 709402 531822 709638
rect 531266 709082 531502 709318
rect 531586 709082 531822 709318
rect 527546 707482 527782 707718
rect 527866 707482 528102 707718
rect 527546 707162 527782 707398
rect 527866 707162 528102 707398
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 552986 710362 553222 710598
rect 553306 710362 553542 710598
rect 552986 710042 553222 710278
rect 553306 710042 553542 710278
rect 549266 708442 549502 708678
rect 549586 708442 549822 708678
rect 549266 708122 549502 708358
rect 549586 708122 549822 708358
rect 545546 706522 545782 706758
rect 545866 706522 546102 706758
rect 545546 706202 545782 706438
rect 545866 706202 546102 706438
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 570986 711322 571222 711558
rect 571306 711322 571542 711558
rect 570986 711002 571222 711238
rect 571306 711002 571542 711238
rect 567266 709402 567502 709638
rect 567586 709402 567822 709638
rect 567266 709082 567502 709318
rect 567586 709082 567822 709318
rect 563546 707482 563782 707718
rect 563866 707482 564102 707718
rect 563546 707162 563782 707398
rect 563866 707162 564102 707398
rect 559826 705562 560062 705798
rect 560146 705562 560382 705798
rect 559826 705242 560062 705478
rect 560146 705242 560382 705478
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect 8250 687218 8486 687454
rect 8250 686898 8486 687134
rect 38970 687218 39206 687454
rect 38970 686898 39206 687134
rect 69690 687218 69926 687454
rect 69690 686898 69926 687134
rect 100410 687218 100646 687454
rect 100410 686898 100646 687134
rect 131130 687218 131366 687454
rect 131130 686898 131366 687134
rect 161850 687218 162086 687454
rect 161850 686898 162086 687134
rect 192570 687218 192806 687454
rect 192570 686898 192806 687134
rect 223290 687218 223526 687454
rect 223290 686898 223526 687134
rect 254010 687218 254246 687454
rect 254010 686898 254246 687134
rect 284730 687218 284966 687454
rect 284730 686898 284966 687134
rect 315450 687218 315686 687454
rect 315450 686898 315686 687134
rect 346170 687218 346406 687454
rect 346170 686898 346406 687134
rect 376890 687218 377126 687454
rect 376890 686898 377126 687134
rect 407610 687218 407846 687454
rect 407610 686898 407846 687134
rect 438330 687218 438566 687454
rect 438330 686898 438566 687134
rect 469050 687218 469286 687454
rect 469050 686898 469286 687134
rect 499770 687218 500006 687454
rect 499770 686898 500006 687134
rect 530490 687218 530726 687454
rect 530490 686898 530726 687134
rect 561210 687218 561446 687454
rect 561210 686898 561446 687134
rect 567266 676658 567502 676894
rect 567586 676658 567822 676894
rect 567266 676338 567502 676574
rect 567586 676338 567822 676574
rect 23610 669218 23846 669454
rect 23610 668898 23846 669134
rect 54330 669218 54566 669454
rect 54330 668898 54566 669134
rect 85050 669218 85286 669454
rect 85050 668898 85286 669134
rect 115770 669218 116006 669454
rect 115770 668898 116006 669134
rect 146490 669218 146726 669454
rect 146490 668898 146726 669134
rect 177210 669218 177446 669454
rect 177210 668898 177446 669134
rect 207930 669218 208166 669454
rect 207930 668898 208166 669134
rect 238650 669218 238886 669454
rect 238650 668898 238886 669134
rect 269370 669218 269606 669454
rect 269370 668898 269606 669134
rect 300090 669218 300326 669454
rect 300090 668898 300326 669134
rect 330810 669218 331046 669454
rect 330810 668898 331046 669134
rect 361530 669218 361766 669454
rect 361530 668898 361766 669134
rect 392250 669218 392486 669454
rect 392250 668898 392486 669134
rect 422970 669218 423206 669454
rect 422970 668898 423206 669134
rect 453690 669218 453926 669454
rect 453690 668898 453926 669134
rect 484410 669218 484646 669454
rect 484410 668898 484646 669134
rect 515130 669218 515366 669454
rect 515130 668898 515366 669134
rect 545850 669218 546086 669454
rect 545850 668898 546086 669134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect 8250 651218 8486 651454
rect 8250 650898 8486 651134
rect 38970 651218 39206 651454
rect 38970 650898 39206 651134
rect 69690 651218 69926 651454
rect 69690 650898 69926 651134
rect 100410 651218 100646 651454
rect 100410 650898 100646 651134
rect 131130 651218 131366 651454
rect 131130 650898 131366 651134
rect 161850 651218 162086 651454
rect 161850 650898 162086 651134
rect 192570 651218 192806 651454
rect 192570 650898 192806 651134
rect 223290 651218 223526 651454
rect 223290 650898 223526 651134
rect 254010 651218 254246 651454
rect 254010 650898 254246 651134
rect 284730 651218 284966 651454
rect 284730 650898 284966 651134
rect 315450 651218 315686 651454
rect 315450 650898 315686 651134
rect 346170 651218 346406 651454
rect 346170 650898 346406 651134
rect 376890 651218 377126 651454
rect 376890 650898 377126 651134
rect 407610 651218 407846 651454
rect 407610 650898 407846 651134
rect 438330 651218 438566 651454
rect 438330 650898 438566 651134
rect 469050 651218 469286 651454
rect 469050 650898 469286 651134
rect 499770 651218 500006 651454
rect 499770 650898 500006 651134
rect 530490 651218 530726 651454
rect 530490 650898 530726 651134
rect 561210 651218 561446 651454
rect 561210 650898 561446 651134
rect 567266 640658 567502 640894
rect 567586 640658 567822 640894
rect 567266 640338 567502 640574
rect 567586 640338 567822 640574
rect 23610 633218 23846 633454
rect 23610 632898 23846 633134
rect 54330 633218 54566 633454
rect 54330 632898 54566 633134
rect 85050 633218 85286 633454
rect 85050 632898 85286 633134
rect 115770 633218 116006 633454
rect 115770 632898 116006 633134
rect 146490 633218 146726 633454
rect 146490 632898 146726 633134
rect 177210 633218 177446 633454
rect 177210 632898 177446 633134
rect 207930 633218 208166 633454
rect 207930 632898 208166 633134
rect 238650 633218 238886 633454
rect 238650 632898 238886 633134
rect 269370 633218 269606 633454
rect 269370 632898 269606 633134
rect 300090 633218 300326 633454
rect 300090 632898 300326 633134
rect 330810 633218 331046 633454
rect 330810 632898 331046 633134
rect 361530 633218 361766 633454
rect 361530 632898 361766 633134
rect 392250 633218 392486 633454
rect 392250 632898 392486 633134
rect 422970 633218 423206 633454
rect 422970 632898 423206 633134
rect 453690 633218 453926 633454
rect 453690 632898 453926 633134
rect 484410 633218 484646 633454
rect 484410 632898 484646 633134
rect 515130 633218 515366 633454
rect 515130 632898 515366 633134
rect 545850 633218 546086 633454
rect 545850 632898 546086 633134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect 8250 615218 8486 615454
rect 8250 614898 8486 615134
rect 38970 615218 39206 615454
rect 38970 614898 39206 615134
rect 69690 615218 69926 615454
rect 69690 614898 69926 615134
rect 100410 615218 100646 615454
rect 100410 614898 100646 615134
rect 131130 615218 131366 615454
rect 131130 614898 131366 615134
rect 161850 615218 162086 615454
rect 161850 614898 162086 615134
rect 192570 615218 192806 615454
rect 192570 614898 192806 615134
rect 223290 615218 223526 615454
rect 223290 614898 223526 615134
rect 254010 615218 254246 615454
rect 254010 614898 254246 615134
rect 284730 615218 284966 615454
rect 284730 614898 284966 615134
rect 315450 615218 315686 615454
rect 315450 614898 315686 615134
rect 346170 615218 346406 615454
rect 346170 614898 346406 615134
rect 376890 615218 377126 615454
rect 376890 614898 377126 615134
rect 407610 615218 407846 615454
rect 407610 614898 407846 615134
rect 438330 615218 438566 615454
rect 438330 614898 438566 615134
rect 469050 615218 469286 615454
rect 469050 614898 469286 615134
rect 499770 615218 500006 615454
rect 499770 614898 500006 615134
rect 530490 615218 530726 615454
rect 530490 614898 530726 615134
rect 561210 615218 561446 615454
rect 561210 614898 561446 615134
rect 567266 604658 567502 604894
rect 567586 604658 567822 604894
rect 567266 604338 567502 604574
rect 567586 604338 567822 604574
rect 23610 597218 23846 597454
rect 23610 596898 23846 597134
rect 54330 597218 54566 597454
rect 54330 596898 54566 597134
rect 85050 597218 85286 597454
rect 85050 596898 85286 597134
rect 115770 597218 116006 597454
rect 115770 596898 116006 597134
rect 146490 597218 146726 597454
rect 146490 596898 146726 597134
rect 177210 597218 177446 597454
rect 177210 596898 177446 597134
rect 207930 597218 208166 597454
rect 207930 596898 208166 597134
rect 238650 597218 238886 597454
rect 238650 596898 238886 597134
rect 269370 597218 269606 597454
rect 269370 596898 269606 597134
rect 300090 597218 300326 597454
rect 300090 596898 300326 597134
rect 330810 597218 331046 597454
rect 330810 596898 331046 597134
rect 361530 597218 361766 597454
rect 361530 596898 361766 597134
rect 392250 597218 392486 597454
rect 392250 596898 392486 597134
rect 422970 597218 423206 597454
rect 422970 596898 423206 597134
rect 453690 597218 453926 597454
rect 453690 596898 453926 597134
rect 484410 597218 484646 597454
rect 484410 596898 484646 597134
rect 515130 597218 515366 597454
rect 515130 596898 515366 597134
rect 545850 597218 546086 597454
rect 545850 596898 546086 597134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect 8250 579218 8486 579454
rect 8250 578898 8486 579134
rect 38970 579218 39206 579454
rect 38970 578898 39206 579134
rect 69690 579218 69926 579454
rect 69690 578898 69926 579134
rect 100410 579218 100646 579454
rect 100410 578898 100646 579134
rect 131130 579218 131366 579454
rect 131130 578898 131366 579134
rect 161850 579218 162086 579454
rect 161850 578898 162086 579134
rect 192570 579218 192806 579454
rect 192570 578898 192806 579134
rect 223290 579218 223526 579454
rect 223290 578898 223526 579134
rect 254010 579218 254246 579454
rect 254010 578898 254246 579134
rect 284730 579218 284966 579454
rect 284730 578898 284966 579134
rect 315450 579218 315686 579454
rect 315450 578898 315686 579134
rect 346170 579218 346406 579454
rect 346170 578898 346406 579134
rect 376890 579218 377126 579454
rect 376890 578898 377126 579134
rect 407610 579218 407846 579454
rect 407610 578898 407846 579134
rect 438330 579218 438566 579454
rect 438330 578898 438566 579134
rect 469050 579218 469286 579454
rect 469050 578898 469286 579134
rect 499770 579218 500006 579454
rect 499770 578898 500006 579134
rect 530490 579218 530726 579454
rect 530490 578898 530726 579134
rect 561210 579218 561446 579454
rect 561210 578898 561446 579134
rect 567266 568658 567502 568894
rect 567586 568658 567822 568894
rect 567266 568338 567502 568574
rect 567586 568338 567822 568574
rect 23610 561218 23846 561454
rect 23610 560898 23846 561134
rect 54330 561218 54566 561454
rect 54330 560898 54566 561134
rect 85050 561218 85286 561454
rect 85050 560898 85286 561134
rect 115770 561218 116006 561454
rect 115770 560898 116006 561134
rect 146490 561218 146726 561454
rect 146490 560898 146726 561134
rect 177210 561218 177446 561454
rect 177210 560898 177446 561134
rect 207930 561218 208166 561454
rect 207930 560898 208166 561134
rect 238650 561218 238886 561454
rect 238650 560898 238886 561134
rect 269370 561218 269606 561454
rect 269370 560898 269606 561134
rect 300090 561218 300326 561454
rect 300090 560898 300326 561134
rect 330810 561218 331046 561454
rect 330810 560898 331046 561134
rect 361530 561218 361766 561454
rect 361530 560898 361766 561134
rect 392250 561218 392486 561454
rect 392250 560898 392486 561134
rect 422970 561218 423206 561454
rect 422970 560898 423206 561134
rect 453690 561218 453926 561454
rect 453690 560898 453926 561134
rect 484410 561218 484646 561454
rect 484410 560898 484646 561134
rect 515130 561218 515366 561454
rect 515130 560898 515366 561134
rect 545850 561218 546086 561454
rect 545850 560898 546086 561134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect 8250 543218 8486 543454
rect 8250 542898 8486 543134
rect 38970 543218 39206 543454
rect 38970 542898 39206 543134
rect 69690 543218 69926 543454
rect 69690 542898 69926 543134
rect 100410 543218 100646 543454
rect 100410 542898 100646 543134
rect 131130 543218 131366 543454
rect 131130 542898 131366 543134
rect 161850 543218 162086 543454
rect 161850 542898 162086 543134
rect 192570 543218 192806 543454
rect 192570 542898 192806 543134
rect 223290 543218 223526 543454
rect 223290 542898 223526 543134
rect 254010 543218 254246 543454
rect 254010 542898 254246 543134
rect 284730 543218 284966 543454
rect 284730 542898 284966 543134
rect 315450 543218 315686 543454
rect 315450 542898 315686 543134
rect 346170 543218 346406 543454
rect 346170 542898 346406 543134
rect 376890 543218 377126 543454
rect 376890 542898 377126 543134
rect 407610 543218 407846 543454
rect 407610 542898 407846 543134
rect 438330 543218 438566 543454
rect 438330 542898 438566 543134
rect 469050 543218 469286 543454
rect 469050 542898 469286 543134
rect 499770 543218 500006 543454
rect 499770 542898 500006 543134
rect 530490 543218 530726 543454
rect 530490 542898 530726 543134
rect 561210 543218 561446 543454
rect 561210 542898 561446 543134
rect 567266 532658 567502 532894
rect 567586 532658 567822 532894
rect 567266 532338 567502 532574
rect 567586 532338 567822 532574
rect 23610 525218 23846 525454
rect 23610 524898 23846 525134
rect 54330 525218 54566 525454
rect 54330 524898 54566 525134
rect 85050 525218 85286 525454
rect 85050 524898 85286 525134
rect 115770 525218 116006 525454
rect 115770 524898 116006 525134
rect 146490 525218 146726 525454
rect 146490 524898 146726 525134
rect 177210 525218 177446 525454
rect 177210 524898 177446 525134
rect 207930 525218 208166 525454
rect 207930 524898 208166 525134
rect 238650 525218 238886 525454
rect 238650 524898 238886 525134
rect 269370 525218 269606 525454
rect 269370 524898 269606 525134
rect 300090 525218 300326 525454
rect 300090 524898 300326 525134
rect 330810 525218 331046 525454
rect 330810 524898 331046 525134
rect 361530 525218 361766 525454
rect 361530 524898 361766 525134
rect 392250 525218 392486 525454
rect 392250 524898 392486 525134
rect 422970 525218 423206 525454
rect 422970 524898 423206 525134
rect 453690 525218 453926 525454
rect 453690 524898 453926 525134
rect 484410 525218 484646 525454
rect 484410 524898 484646 525134
rect 515130 525218 515366 525454
rect 515130 524898 515366 525134
rect 545850 525218 546086 525454
rect 545850 524898 546086 525134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect 8250 507218 8486 507454
rect 8250 506898 8486 507134
rect 38970 507218 39206 507454
rect 38970 506898 39206 507134
rect 69690 507218 69926 507454
rect 69690 506898 69926 507134
rect 100410 507218 100646 507454
rect 100410 506898 100646 507134
rect 131130 507218 131366 507454
rect 131130 506898 131366 507134
rect 161850 507218 162086 507454
rect 161850 506898 162086 507134
rect 192570 507218 192806 507454
rect 192570 506898 192806 507134
rect 223290 507218 223526 507454
rect 223290 506898 223526 507134
rect 254010 507218 254246 507454
rect 254010 506898 254246 507134
rect 284730 507218 284966 507454
rect 284730 506898 284966 507134
rect 315450 507218 315686 507454
rect 315450 506898 315686 507134
rect 346170 507218 346406 507454
rect 346170 506898 346406 507134
rect 376890 507218 377126 507454
rect 376890 506898 377126 507134
rect 407610 507218 407846 507454
rect 407610 506898 407846 507134
rect 438330 507218 438566 507454
rect 438330 506898 438566 507134
rect 469050 507218 469286 507454
rect 469050 506898 469286 507134
rect 499770 507218 500006 507454
rect 499770 506898 500006 507134
rect 530490 507218 530726 507454
rect 530490 506898 530726 507134
rect 561210 507218 561446 507454
rect 561210 506898 561446 507134
rect 567266 496658 567502 496894
rect 567586 496658 567822 496894
rect 567266 496338 567502 496574
rect 567586 496338 567822 496574
rect 23610 489218 23846 489454
rect 23610 488898 23846 489134
rect 54330 489218 54566 489454
rect 54330 488898 54566 489134
rect 85050 489218 85286 489454
rect 85050 488898 85286 489134
rect 115770 489218 116006 489454
rect 115770 488898 116006 489134
rect 146490 489218 146726 489454
rect 146490 488898 146726 489134
rect 177210 489218 177446 489454
rect 177210 488898 177446 489134
rect 207930 489218 208166 489454
rect 207930 488898 208166 489134
rect 238650 489218 238886 489454
rect 238650 488898 238886 489134
rect 269370 489218 269606 489454
rect 269370 488898 269606 489134
rect 300090 489218 300326 489454
rect 300090 488898 300326 489134
rect 330810 489218 331046 489454
rect 330810 488898 331046 489134
rect 361530 489218 361766 489454
rect 361530 488898 361766 489134
rect 392250 489218 392486 489454
rect 392250 488898 392486 489134
rect 422970 489218 423206 489454
rect 422970 488898 423206 489134
rect 453690 489218 453926 489454
rect 453690 488898 453926 489134
rect 484410 489218 484646 489454
rect 484410 488898 484646 489134
rect 515130 489218 515366 489454
rect 515130 488898 515366 489134
rect 545850 489218 546086 489454
rect 545850 488898 546086 489134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect 8250 471218 8486 471454
rect 8250 470898 8486 471134
rect 38970 471218 39206 471454
rect 38970 470898 39206 471134
rect 69690 471218 69926 471454
rect 69690 470898 69926 471134
rect 100410 471218 100646 471454
rect 100410 470898 100646 471134
rect 131130 471218 131366 471454
rect 131130 470898 131366 471134
rect 161850 471218 162086 471454
rect 161850 470898 162086 471134
rect 192570 471218 192806 471454
rect 192570 470898 192806 471134
rect 223290 471218 223526 471454
rect 223290 470898 223526 471134
rect 254010 471218 254246 471454
rect 254010 470898 254246 471134
rect 284730 471218 284966 471454
rect 284730 470898 284966 471134
rect 315450 471218 315686 471454
rect 315450 470898 315686 471134
rect 346170 471218 346406 471454
rect 346170 470898 346406 471134
rect 376890 471218 377126 471454
rect 376890 470898 377126 471134
rect 407610 471218 407846 471454
rect 407610 470898 407846 471134
rect 438330 471218 438566 471454
rect 438330 470898 438566 471134
rect 469050 471218 469286 471454
rect 469050 470898 469286 471134
rect 499770 471218 500006 471454
rect 499770 470898 500006 471134
rect 530490 471218 530726 471454
rect 530490 470898 530726 471134
rect 561210 471218 561446 471454
rect 561210 470898 561446 471134
rect 567266 460658 567502 460894
rect 567586 460658 567822 460894
rect 567266 460338 567502 460574
rect 567586 460338 567822 460574
rect 23610 453218 23846 453454
rect 23610 452898 23846 453134
rect 54330 453218 54566 453454
rect 54330 452898 54566 453134
rect 85050 453218 85286 453454
rect 85050 452898 85286 453134
rect 115770 453218 116006 453454
rect 115770 452898 116006 453134
rect 146490 453218 146726 453454
rect 146490 452898 146726 453134
rect 177210 453218 177446 453454
rect 177210 452898 177446 453134
rect 207930 453218 208166 453454
rect 207930 452898 208166 453134
rect 238650 453218 238886 453454
rect 238650 452898 238886 453134
rect 269370 453218 269606 453454
rect 269370 452898 269606 453134
rect 300090 453218 300326 453454
rect 300090 452898 300326 453134
rect 330810 453218 331046 453454
rect 330810 452898 331046 453134
rect 361530 453218 361766 453454
rect 361530 452898 361766 453134
rect 392250 453218 392486 453454
rect 392250 452898 392486 453134
rect 422970 453218 423206 453454
rect 422970 452898 423206 453134
rect 453690 453218 453926 453454
rect 453690 452898 453926 453134
rect 484410 453218 484646 453454
rect 484410 452898 484646 453134
rect 515130 453218 515366 453454
rect 515130 452898 515366 453134
rect 545850 453218 546086 453454
rect 545850 452898 546086 453134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect 8250 435218 8486 435454
rect 8250 434898 8486 435134
rect 38970 435218 39206 435454
rect 38970 434898 39206 435134
rect 69690 435218 69926 435454
rect 69690 434898 69926 435134
rect 100410 435218 100646 435454
rect 100410 434898 100646 435134
rect 131130 435218 131366 435454
rect 131130 434898 131366 435134
rect 161850 435218 162086 435454
rect 161850 434898 162086 435134
rect 192570 435218 192806 435454
rect 192570 434898 192806 435134
rect 223290 435218 223526 435454
rect 223290 434898 223526 435134
rect 254010 435218 254246 435454
rect 254010 434898 254246 435134
rect 284730 435218 284966 435454
rect 284730 434898 284966 435134
rect 315450 435218 315686 435454
rect 315450 434898 315686 435134
rect 346170 435218 346406 435454
rect 346170 434898 346406 435134
rect 376890 435218 377126 435454
rect 376890 434898 377126 435134
rect 407610 435218 407846 435454
rect 407610 434898 407846 435134
rect 438330 435218 438566 435454
rect 438330 434898 438566 435134
rect 469050 435218 469286 435454
rect 469050 434898 469286 435134
rect 499770 435218 500006 435454
rect 499770 434898 500006 435134
rect 530490 435218 530726 435454
rect 530490 434898 530726 435134
rect 561210 435218 561446 435454
rect 561210 434898 561446 435134
rect 567266 424658 567502 424894
rect 567586 424658 567822 424894
rect 567266 424338 567502 424574
rect 567586 424338 567822 424574
rect 23610 417218 23846 417454
rect 23610 416898 23846 417134
rect 54330 417218 54566 417454
rect 54330 416898 54566 417134
rect 85050 417218 85286 417454
rect 85050 416898 85286 417134
rect 115770 417218 116006 417454
rect 115770 416898 116006 417134
rect 146490 417218 146726 417454
rect 146490 416898 146726 417134
rect 177210 417218 177446 417454
rect 177210 416898 177446 417134
rect 207930 417218 208166 417454
rect 207930 416898 208166 417134
rect 238650 417218 238886 417454
rect 238650 416898 238886 417134
rect 269370 417218 269606 417454
rect 269370 416898 269606 417134
rect 300090 417218 300326 417454
rect 300090 416898 300326 417134
rect 330810 417218 331046 417454
rect 330810 416898 331046 417134
rect 361530 417218 361766 417454
rect 361530 416898 361766 417134
rect 392250 417218 392486 417454
rect 392250 416898 392486 417134
rect 422970 417218 423206 417454
rect 422970 416898 423206 417134
rect 453690 417218 453926 417454
rect 453690 416898 453926 417134
rect 484410 417218 484646 417454
rect 484410 416898 484646 417134
rect 515130 417218 515366 417454
rect 515130 416898 515366 417134
rect 545850 417218 546086 417454
rect 545850 416898 546086 417134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect 8250 399218 8486 399454
rect 8250 398898 8486 399134
rect 38970 399218 39206 399454
rect 38970 398898 39206 399134
rect 69690 399218 69926 399454
rect 69690 398898 69926 399134
rect 100410 399218 100646 399454
rect 100410 398898 100646 399134
rect 131130 399218 131366 399454
rect 131130 398898 131366 399134
rect 161850 399218 162086 399454
rect 161850 398898 162086 399134
rect 192570 399218 192806 399454
rect 192570 398898 192806 399134
rect 223290 399218 223526 399454
rect 223290 398898 223526 399134
rect 254010 399218 254246 399454
rect 254010 398898 254246 399134
rect 284730 399218 284966 399454
rect 284730 398898 284966 399134
rect 315450 399218 315686 399454
rect 315450 398898 315686 399134
rect 346170 399218 346406 399454
rect 346170 398898 346406 399134
rect 376890 399218 377126 399454
rect 376890 398898 377126 399134
rect 407610 399218 407846 399454
rect 407610 398898 407846 399134
rect 438330 399218 438566 399454
rect 438330 398898 438566 399134
rect 469050 399218 469286 399454
rect 469050 398898 469286 399134
rect 499770 399218 500006 399454
rect 499770 398898 500006 399134
rect 530490 399218 530726 399454
rect 530490 398898 530726 399134
rect 561210 399218 561446 399454
rect 561210 398898 561446 399134
rect 567266 388658 567502 388894
rect 567586 388658 567822 388894
rect 567266 388338 567502 388574
rect 567586 388338 567822 388574
rect 23610 381218 23846 381454
rect 23610 380898 23846 381134
rect 54330 381218 54566 381454
rect 54330 380898 54566 381134
rect 85050 381218 85286 381454
rect 85050 380898 85286 381134
rect 115770 381218 116006 381454
rect 115770 380898 116006 381134
rect 146490 381218 146726 381454
rect 146490 380898 146726 381134
rect 177210 381218 177446 381454
rect 177210 380898 177446 381134
rect 207930 381218 208166 381454
rect 207930 380898 208166 381134
rect 238650 381218 238886 381454
rect 238650 380898 238886 381134
rect 269370 381218 269606 381454
rect 269370 380898 269606 381134
rect 300090 381218 300326 381454
rect 300090 380898 300326 381134
rect 330810 381218 331046 381454
rect 330810 380898 331046 381134
rect 361530 381218 361766 381454
rect 361530 380898 361766 381134
rect 392250 381218 392486 381454
rect 392250 380898 392486 381134
rect 422970 381218 423206 381454
rect 422970 380898 423206 381134
rect 453690 381218 453926 381454
rect 453690 380898 453926 381134
rect 484410 381218 484646 381454
rect 484410 380898 484646 381134
rect 515130 381218 515366 381454
rect 515130 380898 515366 381134
rect 545850 381218 546086 381454
rect 545850 380898 546086 381134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect 8250 363218 8486 363454
rect 8250 362898 8486 363134
rect 38970 363218 39206 363454
rect 38970 362898 39206 363134
rect 69690 363218 69926 363454
rect 69690 362898 69926 363134
rect 100410 363218 100646 363454
rect 100410 362898 100646 363134
rect 131130 363218 131366 363454
rect 131130 362898 131366 363134
rect 161850 363218 162086 363454
rect 161850 362898 162086 363134
rect 192570 363218 192806 363454
rect 192570 362898 192806 363134
rect 223290 363218 223526 363454
rect 223290 362898 223526 363134
rect 254010 363218 254246 363454
rect 254010 362898 254246 363134
rect 284730 363218 284966 363454
rect 284730 362898 284966 363134
rect 315450 363218 315686 363454
rect 315450 362898 315686 363134
rect 346170 363218 346406 363454
rect 346170 362898 346406 363134
rect 376890 363218 377126 363454
rect 376890 362898 377126 363134
rect 407610 363218 407846 363454
rect 407610 362898 407846 363134
rect 438330 363218 438566 363454
rect 438330 362898 438566 363134
rect 469050 363218 469286 363454
rect 469050 362898 469286 363134
rect 499770 363218 500006 363454
rect 499770 362898 500006 363134
rect 530490 363218 530726 363454
rect 530490 362898 530726 363134
rect 561210 363218 561446 363454
rect 561210 362898 561446 363134
rect 567266 352658 567502 352894
rect 567586 352658 567822 352894
rect 567266 352338 567502 352574
rect 567586 352338 567822 352574
rect 23610 345218 23846 345454
rect 23610 344898 23846 345134
rect 54330 345218 54566 345454
rect 54330 344898 54566 345134
rect 85050 345218 85286 345454
rect 85050 344898 85286 345134
rect 115770 345218 116006 345454
rect 115770 344898 116006 345134
rect 146490 345218 146726 345454
rect 146490 344898 146726 345134
rect 177210 345218 177446 345454
rect 177210 344898 177446 345134
rect 207930 345218 208166 345454
rect 207930 344898 208166 345134
rect 238650 345218 238886 345454
rect 238650 344898 238886 345134
rect 269370 345218 269606 345454
rect 269370 344898 269606 345134
rect 300090 345218 300326 345454
rect 300090 344898 300326 345134
rect 330810 345218 331046 345454
rect 330810 344898 331046 345134
rect 361530 345218 361766 345454
rect 361530 344898 361766 345134
rect 392250 345218 392486 345454
rect 392250 344898 392486 345134
rect 422970 345218 423206 345454
rect 422970 344898 423206 345134
rect 453690 345218 453926 345454
rect 453690 344898 453926 345134
rect 484410 345218 484646 345454
rect 484410 344898 484646 345134
rect 515130 345218 515366 345454
rect 515130 344898 515366 345134
rect 545850 345218 546086 345454
rect 545850 344898 546086 345134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect 8250 327218 8486 327454
rect 8250 326898 8486 327134
rect 38970 327218 39206 327454
rect 38970 326898 39206 327134
rect 69690 327218 69926 327454
rect 69690 326898 69926 327134
rect 100410 327218 100646 327454
rect 100410 326898 100646 327134
rect 131130 327218 131366 327454
rect 131130 326898 131366 327134
rect 161850 327218 162086 327454
rect 161850 326898 162086 327134
rect 192570 327218 192806 327454
rect 192570 326898 192806 327134
rect 223290 327218 223526 327454
rect 223290 326898 223526 327134
rect 254010 327218 254246 327454
rect 254010 326898 254246 327134
rect 284730 327218 284966 327454
rect 284730 326898 284966 327134
rect 315450 327218 315686 327454
rect 315450 326898 315686 327134
rect 346170 327218 346406 327454
rect 346170 326898 346406 327134
rect 376890 327218 377126 327454
rect 376890 326898 377126 327134
rect 407610 327218 407846 327454
rect 407610 326898 407846 327134
rect 438330 327218 438566 327454
rect 438330 326898 438566 327134
rect 469050 327218 469286 327454
rect 469050 326898 469286 327134
rect 499770 327218 500006 327454
rect 499770 326898 500006 327134
rect 530490 327218 530726 327454
rect 530490 326898 530726 327134
rect 561210 327218 561446 327454
rect 561210 326898 561446 327134
rect 567266 316658 567502 316894
rect 567586 316658 567822 316894
rect 567266 316338 567502 316574
rect 567586 316338 567822 316574
rect 23610 309218 23846 309454
rect 23610 308898 23846 309134
rect 54330 309218 54566 309454
rect 54330 308898 54566 309134
rect 85050 309218 85286 309454
rect 85050 308898 85286 309134
rect 115770 309218 116006 309454
rect 115770 308898 116006 309134
rect 146490 309218 146726 309454
rect 146490 308898 146726 309134
rect 177210 309218 177446 309454
rect 177210 308898 177446 309134
rect 207930 309218 208166 309454
rect 207930 308898 208166 309134
rect 238650 309218 238886 309454
rect 238650 308898 238886 309134
rect 269370 309218 269606 309454
rect 269370 308898 269606 309134
rect 300090 309218 300326 309454
rect 300090 308898 300326 309134
rect 330810 309218 331046 309454
rect 330810 308898 331046 309134
rect 361530 309218 361766 309454
rect 361530 308898 361766 309134
rect 392250 309218 392486 309454
rect 392250 308898 392486 309134
rect 422970 309218 423206 309454
rect 422970 308898 423206 309134
rect 453690 309218 453926 309454
rect 453690 308898 453926 309134
rect 484410 309218 484646 309454
rect 484410 308898 484646 309134
rect 515130 309218 515366 309454
rect 515130 308898 515366 309134
rect 545850 309218 546086 309454
rect 545850 308898 546086 309134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect 8250 291218 8486 291454
rect 8250 290898 8486 291134
rect 38970 291218 39206 291454
rect 38970 290898 39206 291134
rect 69690 291218 69926 291454
rect 69690 290898 69926 291134
rect 100410 291218 100646 291454
rect 100410 290898 100646 291134
rect 131130 291218 131366 291454
rect 131130 290898 131366 291134
rect 161850 291218 162086 291454
rect 161850 290898 162086 291134
rect 192570 291218 192806 291454
rect 192570 290898 192806 291134
rect 223290 291218 223526 291454
rect 223290 290898 223526 291134
rect 254010 291218 254246 291454
rect 254010 290898 254246 291134
rect 284730 291218 284966 291454
rect 284730 290898 284966 291134
rect 315450 291218 315686 291454
rect 315450 290898 315686 291134
rect 346170 291218 346406 291454
rect 346170 290898 346406 291134
rect 376890 291218 377126 291454
rect 376890 290898 377126 291134
rect 407610 291218 407846 291454
rect 407610 290898 407846 291134
rect 438330 291218 438566 291454
rect 438330 290898 438566 291134
rect 469050 291218 469286 291454
rect 469050 290898 469286 291134
rect 499770 291218 500006 291454
rect 499770 290898 500006 291134
rect 530490 291218 530726 291454
rect 530490 290898 530726 291134
rect 561210 291218 561446 291454
rect 561210 290898 561446 291134
rect 567266 280658 567502 280894
rect 567586 280658 567822 280894
rect 567266 280338 567502 280574
rect 567586 280338 567822 280574
rect 23610 273218 23846 273454
rect 23610 272898 23846 273134
rect 54330 273218 54566 273454
rect 54330 272898 54566 273134
rect 85050 273218 85286 273454
rect 85050 272898 85286 273134
rect 115770 273218 116006 273454
rect 115770 272898 116006 273134
rect 146490 273218 146726 273454
rect 146490 272898 146726 273134
rect 177210 273218 177446 273454
rect 177210 272898 177446 273134
rect 207930 273218 208166 273454
rect 207930 272898 208166 273134
rect 238650 273218 238886 273454
rect 238650 272898 238886 273134
rect 269370 273218 269606 273454
rect 269370 272898 269606 273134
rect 300090 273218 300326 273454
rect 300090 272898 300326 273134
rect 330810 273218 331046 273454
rect 330810 272898 331046 273134
rect 361530 273218 361766 273454
rect 361530 272898 361766 273134
rect 392250 273218 392486 273454
rect 392250 272898 392486 273134
rect 422970 273218 423206 273454
rect 422970 272898 423206 273134
rect 453690 273218 453926 273454
rect 453690 272898 453926 273134
rect 484410 273218 484646 273454
rect 484410 272898 484646 273134
rect 515130 273218 515366 273454
rect 515130 272898 515366 273134
rect 545850 273218 546086 273454
rect 545850 272898 546086 273134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect 8250 255218 8486 255454
rect 8250 254898 8486 255134
rect 38970 255218 39206 255454
rect 38970 254898 39206 255134
rect 69690 255218 69926 255454
rect 69690 254898 69926 255134
rect 100410 255218 100646 255454
rect 100410 254898 100646 255134
rect 131130 255218 131366 255454
rect 131130 254898 131366 255134
rect 161850 255218 162086 255454
rect 161850 254898 162086 255134
rect 192570 255218 192806 255454
rect 192570 254898 192806 255134
rect 223290 255218 223526 255454
rect 223290 254898 223526 255134
rect 254010 255218 254246 255454
rect 254010 254898 254246 255134
rect 284730 255218 284966 255454
rect 284730 254898 284966 255134
rect 315450 255218 315686 255454
rect 315450 254898 315686 255134
rect 346170 255218 346406 255454
rect 346170 254898 346406 255134
rect 376890 255218 377126 255454
rect 376890 254898 377126 255134
rect 407610 255218 407846 255454
rect 407610 254898 407846 255134
rect 438330 255218 438566 255454
rect 438330 254898 438566 255134
rect 469050 255218 469286 255454
rect 469050 254898 469286 255134
rect 499770 255218 500006 255454
rect 499770 254898 500006 255134
rect 530490 255218 530726 255454
rect 530490 254898 530726 255134
rect 561210 255218 561446 255454
rect 561210 254898 561446 255134
rect 567266 244658 567502 244894
rect 567586 244658 567822 244894
rect 567266 244338 567502 244574
rect 567586 244338 567822 244574
rect 23610 237218 23846 237454
rect 23610 236898 23846 237134
rect 54330 237218 54566 237454
rect 54330 236898 54566 237134
rect 85050 237218 85286 237454
rect 85050 236898 85286 237134
rect 115770 237218 116006 237454
rect 115770 236898 116006 237134
rect 146490 237218 146726 237454
rect 146490 236898 146726 237134
rect 177210 237218 177446 237454
rect 177210 236898 177446 237134
rect 207930 237218 208166 237454
rect 207930 236898 208166 237134
rect 238650 237218 238886 237454
rect 238650 236898 238886 237134
rect 269370 237218 269606 237454
rect 269370 236898 269606 237134
rect 300090 237218 300326 237454
rect 300090 236898 300326 237134
rect 330810 237218 331046 237454
rect 330810 236898 331046 237134
rect 361530 237218 361766 237454
rect 361530 236898 361766 237134
rect 392250 237218 392486 237454
rect 392250 236898 392486 237134
rect 422970 237218 423206 237454
rect 422970 236898 423206 237134
rect 453690 237218 453926 237454
rect 453690 236898 453926 237134
rect 484410 237218 484646 237454
rect 484410 236898 484646 237134
rect 515130 237218 515366 237454
rect 515130 236898 515366 237134
rect 545850 237218 546086 237454
rect 545850 236898 546086 237134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect 8250 219218 8486 219454
rect 8250 218898 8486 219134
rect 38970 219218 39206 219454
rect 38970 218898 39206 219134
rect 69690 219218 69926 219454
rect 69690 218898 69926 219134
rect 100410 219218 100646 219454
rect 100410 218898 100646 219134
rect 131130 219218 131366 219454
rect 131130 218898 131366 219134
rect 161850 219218 162086 219454
rect 161850 218898 162086 219134
rect 192570 219218 192806 219454
rect 192570 218898 192806 219134
rect 223290 219218 223526 219454
rect 223290 218898 223526 219134
rect 254010 219218 254246 219454
rect 254010 218898 254246 219134
rect 284730 219218 284966 219454
rect 284730 218898 284966 219134
rect 315450 219218 315686 219454
rect 315450 218898 315686 219134
rect 346170 219218 346406 219454
rect 346170 218898 346406 219134
rect 376890 219218 377126 219454
rect 376890 218898 377126 219134
rect 407610 219218 407846 219454
rect 407610 218898 407846 219134
rect 438330 219218 438566 219454
rect 438330 218898 438566 219134
rect 469050 219218 469286 219454
rect 469050 218898 469286 219134
rect 499770 219218 500006 219454
rect 499770 218898 500006 219134
rect 530490 219218 530726 219454
rect 530490 218898 530726 219134
rect 561210 219218 561446 219454
rect 561210 218898 561446 219134
rect 567266 208658 567502 208894
rect 567586 208658 567822 208894
rect 567266 208338 567502 208574
rect 567586 208338 567822 208574
rect 23610 201218 23846 201454
rect 23610 200898 23846 201134
rect 54330 201218 54566 201454
rect 54330 200898 54566 201134
rect 85050 201218 85286 201454
rect 85050 200898 85286 201134
rect 115770 201218 116006 201454
rect 115770 200898 116006 201134
rect 146490 201218 146726 201454
rect 146490 200898 146726 201134
rect 177210 201218 177446 201454
rect 177210 200898 177446 201134
rect 207930 201218 208166 201454
rect 207930 200898 208166 201134
rect 238650 201218 238886 201454
rect 238650 200898 238886 201134
rect 269370 201218 269606 201454
rect 269370 200898 269606 201134
rect 300090 201218 300326 201454
rect 300090 200898 300326 201134
rect 330810 201218 331046 201454
rect 330810 200898 331046 201134
rect 361530 201218 361766 201454
rect 361530 200898 361766 201134
rect 392250 201218 392486 201454
rect 392250 200898 392486 201134
rect 422970 201218 423206 201454
rect 422970 200898 423206 201134
rect 453690 201218 453926 201454
rect 453690 200898 453926 201134
rect 484410 201218 484646 201454
rect 484410 200898 484646 201134
rect 515130 201218 515366 201454
rect 515130 200898 515366 201134
rect 545850 201218 546086 201454
rect 545850 200898 546086 201134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect 8250 183218 8486 183454
rect 8250 182898 8486 183134
rect 38970 183218 39206 183454
rect 38970 182898 39206 183134
rect 69690 183218 69926 183454
rect 69690 182898 69926 183134
rect 100410 183218 100646 183454
rect 100410 182898 100646 183134
rect 131130 183218 131366 183454
rect 131130 182898 131366 183134
rect 161850 183218 162086 183454
rect 161850 182898 162086 183134
rect 192570 183218 192806 183454
rect 192570 182898 192806 183134
rect 223290 183218 223526 183454
rect 223290 182898 223526 183134
rect 254010 183218 254246 183454
rect 254010 182898 254246 183134
rect 284730 183218 284966 183454
rect 284730 182898 284966 183134
rect 315450 183218 315686 183454
rect 315450 182898 315686 183134
rect 346170 183218 346406 183454
rect 346170 182898 346406 183134
rect 376890 183218 377126 183454
rect 376890 182898 377126 183134
rect 407610 183218 407846 183454
rect 407610 182898 407846 183134
rect 438330 183218 438566 183454
rect 438330 182898 438566 183134
rect 469050 183218 469286 183454
rect 469050 182898 469286 183134
rect 499770 183218 500006 183454
rect 499770 182898 500006 183134
rect 530490 183218 530726 183454
rect 530490 182898 530726 183134
rect 561210 183218 561446 183454
rect 561210 182898 561446 183134
rect 567266 172658 567502 172894
rect 567586 172658 567822 172894
rect 567266 172338 567502 172574
rect 567586 172338 567822 172574
rect 23610 165218 23846 165454
rect 23610 164898 23846 165134
rect 54330 165218 54566 165454
rect 54330 164898 54566 165134
rect 85050 165218 85286 165454
rect 85050 164898 85286 165134
rect 115770 165218 116006 165454
rect 115770 164898 116006 165134
rect 146490 165218 146726 165454
rect 146490 164898 146726 165134
rect 177210 165218 177446 165454
rect 177210 164898 177446 165134
rect 207930 165218 208166 165454
rect 207930 164898 208166 165134
rect 238650 165218 238886 165454
rect 238650 164898 238886 165134
rect 269370 165218 269606 165454
rect 269370 164898 269606 165134
rect 300090 165218 300326 165454
rect 300090 164898 300326 165134
rect 330810 165218 331046 165454
rect 330810 164898 331046 165134
rect 361530 165218 361766 165454
rect 361530 164898 361766 165134
rect 392250 165218 392486 165454
rect 392250 164898 392486 165134
rect 422970 165218 423206 165454
rect 422970 164898 423206 165134
rect 453690 165218 453926 165454
rect 453690 164898 453926 165134
rect 484410 165218 484646 165454
rect 484410 164898 484646 165134
rect 515130 165218 515366 165454
rect 515130 164898 515366 165134
rect 545850 165218 546086 165454
rect 545850 164898 546086 165134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect 8250 147218 8486 147454
rect 8250 146898 8486 147134
rect 38970 147218 39206 147454
rect 38970 146898 39206 147134
rect 69690 147218 69926 147454
rect 69690 146898 69926 147134
rect 100410 147218 100646 147454
rect 100410 146898 100646 147134
rect 131130 147218 131366 147454
rect 131130 146898 131366 147134
rect 161850 147218 162086 147454
rect 161850 146898 162086 147134
rect 192570 147218 192806 147454
rect 192570 146898 192806 147134
rect 223290 147218 223526 147454
rect 223290 146898 223526 147134
rect 254010 147218 254246 147454
rect 254010 146898 254246 147134
rect 284730 147218 284966 147454
rect 284730 146898 284966 147134
rect 315450 147218 315686 147454
rect 315450 146898 315686 147134
rect 346170 147218 346406 147454
rect 346170 146898 346406 147134
rect 376890 147218 377126 147454
rect 376890 146898 377126 147134
rect 407610 147218 407846 147454
rect 407610 146898 407846 147134
rect 438330 147218 438566 147454
rect 438330 146898 438566 147134
rect 469050 147218 469286 147454
rect 469050 146898 469286 147134
rect 499770 147218 500006 147454
rect 499770 146898 500006 147134
rect 530490 147218 530726 147454
rect 530490 146898 530726 147134
rect 561210 147218 561446 147454
rect 561210 146898 561446 147134
rect 567266 136658 567502 136894
rect 567586 136658 567822 136894
rect 567266 136338 567502 136574
rect 567586 136338 567822 136574
rect 23610 129218 23846 129454
rect 23610 128898 23846 129134
rect 54330 129218 54566 129454
rect 54330 128898 54566 129134
rect 85050 129218 85286 129454
rect 85050 128898 85286 129134
rect 115770 129218 116006 129454
rect 115770 128898 116006 129134
rect 146490 129218 146726 129454
rect 146490 128898 146726 129134
rect 177210 129218 177446 129454
rect 177210 128898 177446 129134
rect 207930 129218 208166 129454
rect 207930 128898 208166 129134
rect 238650 129218 238886 129454
rect 238650 128898 238886 129134
rect 269370 129218 269606 129454
rect 269370 128898 269606 129134
rect 300090 129218 300326 129454
rect 300090 128898 300326 129134
rect 330810 129218 331046 129454
rect 330810 128898 331046 129134
rect 361530 129218 361766 129454
rect 361530 128898 361766 129134
rect 392250 129218 392486 129454
rect 392250 128898 392486 129134
rect 422970 129218 423206 129454
rect 422970 128898 423206 129134
rect 453690 129218 453926 129454
rect 453690 128898 453926 129134
rect 484410 129218 484646 129454
rect 484410 128898 484646 129134
rect 515130 129218 515366 129454
rect 515130 128898 515366 129134
rect 545850 129218 546086 129454
rect 545850 128898 546086 129134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect 8250 111218 8486 111454
rect 8250 110898 8486 111134
rect 38970 111218 39206 111454
rect 38970 110898 39206 111134
rect 69690 111218 69926 111454
rect 69690 110898 69926 111134
rect 100410 111218 100646 111454
rect 100410 110898 100646 111134
rect 131130 111218 131366 111454
rect 131130 110898 131366 111134
rect 161850 111218 162086 111454
rect 161850 110898 162086 111134
rect 192570 111218 192806 111454
rect 192570 110898 192806 111134
rect 223290 111218 223526 111454
rect 223290 110898 223526 111134
rect 254010 111218 254246 111454
rect 254010 110898 254246 111134
rect 284730 111218 284966 111454
rect 284730 110898 284966 111134
rect 315450 111218 315686 111454
rect 315450 110898 315686 111134
rect 346170 111218 346406 111454
rect 346170 110898 346406 111134
rect 376890 111218 377126 111454
rect 376890 110898 377126 111134
rect 407610 111218 407846 111454
rect 407610 110898 407846 111134
rect 438330 111218 438566 111454
rect 438330 110898 438566 111134
rect 469050 111218 469286 111454
rect 469050 110898 469286 111134
rect 499770 111218 500006 111454
rect 499770 110898 500006 111134
rect 530490 111218 530726 111454
rect 530490 110898 530726 111134
rect 561210 111218 561446 111454
rect 561210 110898 561446 111134
rect 567266 100658 567502 100894
rect 567586 100658 567822 100894
rect 567266 100338 567502 100574
rect 567586 100338 567822 100574
rect 23610 93218 23846 93454
rect 23610 92898 23846 93134
rect 54330 93218 54566 93454
rect 54330 92898 54566 93134
rect 85050 93218 85286 93454
rect 85050 92898 85286 93134
rect 115770 93218 116006 93454
rect 115770 92898 116006 93134
rect 146490 93218 146726 93454
rect 146490 92898 146726 93134
rect 177210 93218 177446 93454
rect 177210 92898 177446 93134
rect 207930 93218 208166 93454
rect 207930 92898 208166 93134
rect 238650 93218 238886 93454
rect 238650 92898 238886 93134
rect 269370 93218 269606 93454
rect 269370 92898 269606 93134
rect 300090 93218 300326 93454
rect 300090 92898 300326 93134
rect 330810 93218 331046 93454
rect 330810 92898 331046 93134
rect 361530 93218 361766 93454
rect 361530 92898 361766 93134
rect 392250 93218 392486 93454
rect 392250 92898 392486 93134
rect 422970 93218 423206 93454
rect 422970 92898 423206 93134
rect 453690 93218 453926 93454
rect 453690 92898 453926 93134
rect 484410 93218 484646 93454
rect 484410 92898 484646 93134
rect 515130 93218 515366 93454
rect 515130 92898 515366 93134
rect 545850 93218 546086 93454
rect 545850 92898 546086 93134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect 8250 75218 8486 75454
rect 8250 74898 8486 75134
rect 38970 75218 39206 75454
rect 38970 74898 39206 75134
rect 69690 75218 69926 75454
rect 69690 74898 69926 75134
rect 100410 75218 100646 75454
rect 100410 74898 100646 75134
rect 131130 75218 131366 75454
rect 131130 74898 131366 75134
rect 161850 75218 162086 75454
rect 161850 74898 162086 75134
rect 192570 75218 192806 75454
rect 192570 74898 192806 75134
rect 223290 75218 223526 75454
rect 223290 74898 223526 75134
rect 254010 75218 254246 75454
rect 254010 74898 254246 75134
rect 284730 75218 284966 75454
rect 284730 74898 284966 75134
rect 315450 75218 315686 75454
rect 315450 74898 315686 75134
rect 346170 75218 346406 75454
rect 346170 74898 346406 75134
rect 376890 75218 377126 75454
rect 376890 74898 377126 75134
rect 407610 75218 407846 75454
rect 407610 74898 407846 75134
rect 438330 75218 438566 75454
rect 438330 74898 438566 75134
rect 469050 75218 469286 75454
rect 469050 74898 469286 75134
rect 499770 75218 500006 75454
rect 499770 74898 500006 75134
rect 530490 75218 530726 75454
rect 530490 74898 530726 75134
rect 561210 75218 561446 75454
rect 561210 74898 561446 75134
rect 567266 64658 567502 64894
rect 567586 64658 567822 64894
rect 567266 64338 567502 64574
rect 567586 64338 567822 64574
rect 23610 57218 23846 57454
rect 23610 56898 23846 57134
rect 54330 57218 54566 57454
rect 54330 56898 54566 57134
rect 85050 57218 85286 57454
rect 85050 56898 85286 57134
rect 115770 57218 116006 57454
rect 115770 56898 116006 57134
rect 146490 57218 146726 57454
rect 146490 56898 146726 57134
rect 177210 57218 177446 57454
rect 177210 56898 177446 57134
rect 207930 57218 208166 57454
rect 207930 56898 208166 57134
rect 238650 57218 238886 57454
rect 238650 56898 238886 57134
rect 269370 57218 269606 57454
rect 269370 56898 269606 57134
rect 300090 57218 300326 57454
rect 300090 56898 300326 57134
rect 330810 57218 331046 57454
rect 330810 56898 331046 57134
rect 361530 57218 361766 57454
rect 361530 56898 361766 57134
rect 392250 57218 392486 57454
rect 392250 56898 392486 57134
rect 422970 57218 423206 57454
rect 422970 56898 423206 57134
rect 453690 57218 453926 57454
rect 453690 56898 453926 57134
rect 484410 57218 484646 57454
rect 484410 56898 484646 57134
rect 515130 57218 515366 57454
rect 515130 56898 515366 57134
rect 545850 57218 546086 57454
rect 545850 56898 546086 57134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect 8250 39218 8486 39454
rect 8250 38898 8486 39134
rect 38970 39218 39206 39454
rect 38970 38898 39206 39134
rect 69690 39218 69926 39454
rect 69690 38898 69926 39134
rect 100410 39218 100646 39454
rect 100410 38898 100646 39134
rect 131130 39218 131366 39454
rect 131130 38898 131366 39134
rect 161850 39218 162086 39454
rect 161850 38898 162086 39134
rect 192570 39218 192806 39454
rect 192570 38898 192806 39134
rect 223290 39218 223526 39454
rect 223290 38898 223526 39134
rect 254010 39218 254246 39454
rect 254010 38898 254246 39134
rect 284730 39218 284966 39454
rect 284730 38898 284966 39134
rect 315450 39218 315686 39454
rect 315450 38898 315686 39134
rect 346170 39218 346406 39454
rect 346170 38898 346406 39134
rect 376890 39218 377126 39454
rect 376890 38898 377126 39134
rect 407610 39218 407846 39454
rect 407610 38898 407846 39134
rect 438330 39218 438566 39454
rect 438330 38898 438566 39134
rect 469050 39218 469286 39454
rect 469050 38898 469286 39134
rect 499770 39218 500006 39454
rect 499770 38898 500006 39134
rect 530490 39218 530726 39454
rect 530490 38898 530726 39134
rect 561210 39218 561446 39454
rect 561210 38898 561446 39134
rect 567266 28658 567502 28894
rect 567586 28658 567822 28894
rect 567266 28338 567502 28574
rect 567586 28338 567822 28574
rect 23610 21218 23846 21454
rect 23610 20898 23846 21134
rect 54330 21218 54566 21454
rect 54330 20898 54566 21134
rect 85050 21218 85286 21454
rect 85050 20898 85286 21134
rect 115770 21218 116006 21454
rect 115770 20898 116006 21134
rect 146490 21218 146726 21454
rect 146490 20898 146726 21134
rect 177210 21218 177446 21454
rect 177210 20898 177446 21134
rect 207930 21218 208166 21454
rect 207930 20898 208166 21134
rect 238650 21218 238886 21454
rect 238650 20898 238886 21134
rect 269370 21218 269606 21454
rect 269370 20898 269606 21134
rect 300090 21218 300326 21454
rect 300090 20898 300326 21134
rect 330810 21218 331046 21454
rect 330810 20898 331046 21134
rect 361530 21218 361766 21454
rect 361530 20898 361766 21134
rect 392250 21218 392486 21454
rect 392250 20898 392486 21134
rect 422970 21218 423206 21454
rect 422970 20898 423206 21134
rect 453690 21218 453926 21454
rect 453690 20898 453926 21134
rect 484410 21218 484646 21454
rect 484410 20898 484646 21134
rect 515130 21218 515366 21454
rect 515130 20898 515366 21134
rect 545850 21218 546086 21454
rect 545850 20898 546086 21134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect 8250 3218 8486 3454
rect 8250 2898 8486 3134
rect 38970 3218 39206 3454
rect 38970 2898 39206 3134
rect 69690 3218 69926 3454
rect 69690 2898 69926 3134
rect 100410 3218 100646 3454
rect 100410 2898 100646 3134
rect 131130 3218 131366 3454
rect 131130 2898 131366 3134
rect 161850 3218 162086 3454
rect 161850 2898 162086 3134
rect 192570 3218 192806 3454
rect 192570 2898 192806 3134
rect 223290 3218 223526 3454
rect 223290 2898 223526 3134
rect 254010 3218 254246 3454
rect 254010 2898 254246 3134
rect 284730 3218 284966 3454
rect 284730 2898 284966 3134
rect 315450 3218 315686 3454
rect 315450 2898 315686 3134
rect 346170 3218 346406 3454
rect 346170 2898 346406 3134
rect 376890 3218 377126 3454
rect 376890 2898 377126 3134
rect 407610 3218 407846 3454
rect 407610 2898 407846 3134
rect 438330 3218 438566 3454
rect 438330 2898 438566 3134
rect 469050 3218 469286 3454
rect 469050 2898 469286 3134
rect 499770 3218 500006 3454
rect 499770 2898 500006 3134
rect 530490 3218 530726 3454
rect 530490 2898 530726 3134
rect 561210 3218 561446 3454
rect 561210 2898 561446 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 5546 -2502 5782 -2266
rect 5866 -2502 6102 -2266
rect 5546 -2822 5782 -2586
rect 5866 -2822 6102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 9266 -4422 9502 -4186
rect 9586 -4422 9822 -4186
rect 9266 -4742 9502 -4506
rect 9586 -4742 9822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 23546 -3462 23782 -3226
rect 23866 -3462 24102 -3226
rect 23546 -3782 23782 -3546
rect 23866 -3782 24102 -3546
rect 27266 -5382 27502 -5146
rect 27586 -5382 27822 -5146
rect 27266 -5702 27502 -5466
rect 27586 -5702 27822 -5466
rect 12986 -6342 13222 -6106
rect 13306 -6342 13542 -6106
rect 12986 -6662 13222 -6426
rect 13306 -6662 13542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 41546 -2502 41782 -2266
rect 41866 -2502 42102 -2266
rect 41546 -2822 41782 -2586
rect 41866 -2822 42102 -2586
rect 45266 -4422 45502 -4186
rect 45586 -4422 45822 -4186
rect 45266 -4742 45502 -4506
rect 45586 -4742 45822 -4506
rect 30986 -7302 31222 -7066
rect 31306 -7302 31542 -7066
rect 30986 -7622 31222 -7386
rect 31306 -7622 31542 -7386
rect 59546 -3462 59782 -3226
rect 59866 -3462 60102 -3226
rect 59546 -3782 59782 -3546
rect 59866 -3782 60102 -3546
rect 63266 -5382 63502 -5146
rect 63586 -5382 63822 -5146
rect 63266 -5702 63502 -5466
rect 63586 -5702 63822 -5466
rect 48986 -6342 49222 -6106
rect 49306 -6342 49542 -6106
rect 48986 -6662 49222 -6426
rect 49306 -6662 49542 -6426
rect 77546 -2502 77782 -2266
rect 77866 -2502 78102 -2266
rect 77546 -2822 77782 -2586
rect 77866 -2822 78102 -2586
rect 81266 -4422 81502 -4186
rect 81586 -4422 81822 -4186
rect 81266 -4742 81502 -4506
rect 81586 -4742 81822 -4506
rect 66986 -7302 67222 -7066
rect 67306 -7302 67542 -7066
rect 66986 -7622 67222 -7386
rect 67306 -7622 67542 -7386
rect 95546 -3462 95782 -3226
rect 95866 -3462 96102 -3226
rect 95546 -3782 95782 -3546
rect 95866 -3782 96102 -3546
rect 99266 -5382 99502 -5146
rect 99586 -5382 99822 -5146
rect 99266 -5702 99502 -5466
rect 99586 -5702 99822 -5466
rect 84986 -6342 85222 -6106
rect 85306 -6342 85542 -6106
rect 84986 -6662 85222 -6426
rect 85306 -6662 85542 -6426
rect 113546 -2502 113782 -2266
rect 113866 -2502 114102 -2266
rect 113546 -2822 113782 -2586
rect 113866 -2822 114102 -2586
rect 117266 -4422 117502 -4186
rect 117586 -4422 117822 -4186
rect 117266 -4742 117502 -4506
rect 117586 -4742 117822 -4506
rect 102986 -7302 103222 -7066
rect 103306 -7302 103542 -7066
rect 102986 -7622 103222 -7386
rect 103306 -7622 103542 -7386
rect 131546 -3462 131782 -3226
rect 131866 -3462 132102 -3226
rect 131546 -3782 131782 -3546
rect 131866 -3782 132102 -3546
rect 135266 -5382 135502 -5146
rect 135586 -5382 135822 -5146
rect 135266 -5702 135502 -5466
rect 135586 -5702 135822 -5466
rect 120986 -6342 121222 -6106
rect 121306 -6342 121542 -6106
rect 120986 -6662 121222 -6426
rect 121306 -6662 121542 -6426
rect 149546 -2502 149782 -2266
rect 149866 -2502 150102 -2266
rect 149546 -2822 149782 -2586
rect 149866 -2822 150102 -2586
rect 153266 -4422 153502 -4186
rect 153586 -4422 153822 -4186
rect 153266 -4742 153502 -4506
rect 153586 -4742 153822 -4506
rect 138986 -7302 139222 -7066
rect 139306 -7302 139542 -7066
rect 138986 -7622 139222 -7386
rect 139306 -7622 139542 -7386
rect 167546 -3462 167782 -3226
rect 167866 -3462 168102 -3226
rect 167546 -3782 167782 -3546
rect 167866 -3782 168102 -3546
rect 171266 -5382 171502 -5146
rect 171586 -5382 171822 -5146
rect 171266 -5702 171502 -5466
rect 171586 -5702 171822 -5466
rect 156986 -6342 157222 -6106
rect 157306 -6342 157542 -6106
rect 156986 -6662 157222 -6426
rect 157306 -6662 157542 -6426
rect 185546 -2502 185782 -2266
rect 185866 -2502 186102 -2266
rect 185546 -2822 185782 -2586
rect 185866 -2822 186102 -2586
rect 189266 -4422 189502 -4186
rect 189586 -4422 189822 -4186
rect 189266 -4742 189502 -4506
rect 189586 -4742 189822 -4506
rect 174986 -7302 175222 -7066
rect 175306 -7302 175542 -7066
rect 174986 -7622 175222 -7386
rect 175306 -7622 175542 -7386
rect 203546 -3462 203782 -3226
rect 203866 -3462 204102 -3226
rect 203546 -3782 203782 -3546
rect 203866 -3782 204102 -3546
rect 207266 -5382 207502 -5146
rect 207586 -5382 207822 -5146
rect 207266 -5702 207502 -5466
rect 207586 -5702 207822 -5466
rect 192986 -6342 193222 -6106
rect 193306 -6342 193542 -6106
rect 192986 -6662 193222 -6426
rect 193306 -6662 193542 -6426
rect 221546 -2502 221782 -2266
rect 221866 -2502 222102 -2266
rect 221546 -2822 221782 -2586
rect 221866 -2822 222102 -2586
rect 225266 -4422 225502 -4186
rect 225586 -4422 225822 -4186
rect 225266 -4742 225502 -4506
rect 225586 -4742 225822 -4506
rect 210986 -7302 211222 -7066
rect 211306 -7302 211542 -7066
rect 210986 -7622 211222 -7386
rect 211306 -7622 211542 -7386
rect 239546 -3462 239782 -3226
rect 239866 -3462 240102 -3226
rect 239546 -3782 239782 -3546
rect 239866 -3782 240102 -3546
rect 243266 -5382 243502 -5146
rect 243586 -5382 243822 -5146
rect 243266 -5702 243502 -5466
rect 243586 -5702 243822 -5466
rect 228986 -6342 229222 -6106
rect 229306 -6342 229542 -6106
rect 228986 -6662 229222 -6426
rect 229306 -6662 229542 -6426
rect 257546 -2502 257782 -2266
rect 257866 -2502 258102 -2266
rect 257546 -2822 257782 -2586
rect 257866 -2822 258102 -2586
rect 261266 -4422 261502 -4186
rect 261586 -4422 261822 -4186
rect 261266 -4742 261502 -4506
rect 261586 -4742 261822 -4506
rect 246986 -7302 247222 -7066
rect 247306 -7302 247542 -7066
rect 246986 -7622 247222 -7386
rect 247306 -7622 247542 -7386
rect 275546 -3462 275782 -3226
rect 275866 -3462 276102 -3226
rect 275546 -3782 275782 -3546
rect 275866 -3782 276102 -3546
rect 279266 -5382 279502 -5146
rect 279586 -5382 279822 -5146
rect 279266 -5702 279502 -5466
rect 279586 -5702 279822 -5466
rect 264986 -6342 265222 -6106
rect 265306 -6342 265542 -6106
rect 264986 -6662 265222 -6426
rect 265306 -6662 265542 -6426
rect 293546 -2502 293782 -2266
rect 293866 -2502 294102 -2266
rect 293546 -2822 293782 -2586
rect 293866 -2822 294102 -2586
rect 297266 -4422 297502 -4186
rect 297586 -4422 297822 -4186
rect 297266 -4742 297502 -4506
rect 297586 -4742 297822 -4506
rect 282986 -7302 283222 -7066
rect 283306 -7302 283542 -7066
rect 282986 -7622 283222 -7386
rect 283306 -7622 283542 -7386
rect 311546 -3462 311782 -3226
rect 311866 -3462 312102 -3226
rect 311546 -3782 311782 -3546
rect 311866 -3782 312102 -3546
rect 315266 -5382 315502 -5146
rect 315586 -5382 315822 -5146
rect 315266 -5702 315502 -5466
rect 315586 -5702 315822 -5466
rect 300986 -6342 301222 -6106
rect 301306 -6342 301542 -6106
rect 300986 -6662 301222 -6426
rect 301306 -6662 301542 -6426
rect 329546 -2502 329782 -2266
rect 329866 -2502 330102 -2266
rect 329546 -2822 329782 -2586
rect 329866 -2822 330102 -2586
rect 333266 -4422 333502 -4186
rect 333586 -4422 333822 -4186
rect 333266 -4742 333502 -4506
rect 333586 -4742 333822 -4506
rect 318986 -7302 319222 -7066
rect 319306 -7302 319542 -7066
rect 318986 -7622 319222 -7386
rect 319306 -7622 319542 -7386
rect 347546 -3462 347782 -3226
rect 347866 -3462 348102 -3226
rect 347546 -3782 347782 -3546
rect 347866 -3782 348102 -3546
rect 351266 -5382 351502 -5146
rect 351586 -5382 351822 -5146
rect 351266 -5702 351502 -5466
rect 351586 -5702 351822 -5466
rect 336986 -6342 337222 -6106
rect 337306 -6342 337542 -6106
rect 336986 -6662 337222 -6426
rect 337306 -6662 337542 -6426
rect 365546 -2502 365782 -2266
rect 365866 -2502 366102 -2266
rect 365546 -2822 365782 -2586
rect 365866 -2822 366102 -2586
rect 369266 -4422 369502 -4186
rect 369586 -4422 369822 -4186
rect 369266 -4742 369502 -4506
rect 369586 -4742 369822 -4506
rect 354986 -7302 355222 -7066
rect 355306 -7302 355542 -7066
rect 354986 -7622 355222 -7386
rect 355306 -7622 355542 -7386
rect 383546 -3462 383782 -3226
rect 383866 -3462 384102 -3226
rect 383546 -3782 383782 -3546
rect 383866 -3782 384102 -3546
rect 387266 -5382 387502 -5146
rect 387586 -5382 387822 -5146
rect 387266 -5702 387502 -5466
rect 387586 -5702 387822 -5466
rect 372986 -6342 373222 -6106
rect 373306 -6342 373542 -6106
rect 372986 -6662 373222 -6426
rect 373306 -6662 373542 -6426
rect 401546 -2502 401782 -2266
rect 401866 -2502 402102 -2266
rect 401546 -2822 401782 -2586
rect 401866 -2822 402102 -2586
rect 405266 -4422 405502 -4186
rect 405586 -4422 405822 -4186
rect 405266 -4742 405502 -4506
rect 405586 -4742 405822 -4506
rect 390986 -7302 391222 -7066
rect 391306 -7302 391542 -7066
rect 390986 -7622 391222 -7386
rect 391306 -7622 391542 -7386
rect 419546 -3462 419782 -3226
rect 419866 -3462 420102 -3226
rect 419546 -3782 419782 -3546
rect 419866 -3782 420102 -3546
rect 423266 -5382 423502 -5146
rect 423586 -5382 423822 -5146
rect 423266 -5702 423502 -5466
rect 423586 -5702 423822 -5466
rect 408986 -6342 409222 -6106
rect 409306 -6342 409542 -6106
rect 408986 -6662 409222 -6426
rect 409306 -6662 409542 -6426
rect 437546 -2502 437782 -2266
rect 437866 -2502 438102 -2266
rect 437546 -2822 437782 -2586
rect 437866 -2822 438102 -2586
rect 441266 -4422 441502 -4186
rect 441586 -4422 441822 -4186
rect 441266 -4742 441502 -4506
rect 441586 -4742 441822 -4506
rect 426986 -7302 427222 -7066
rect 427306 -7302 427542 -7066
rect 426986 -7622 427222 -7386
rect 427306 -7622 427542 -7386
rect 455546 -3462 455782 -3226
rect 455866 -3462 456102 -3226
rect 455546 -3782 455782 -3546
rect 455866 -3782 456102 -3546
rect 459266 -5382 459502 -5146
rect 459586 -5382 459822 -5146
rect 459266 -5702 459502 -5466
rect 459586 -5702 459822 -5466
rect 444986 -6342 445222 -6106
rect 445306 -6342 445542 -6106
rect 444986 -6662 445222 -6426
rect 445306 -6662 445542 -6426
rect 473546 -2502 473782 -2266
rect 473866 -2502 474102 -2266
rect 473546 -2822 473782 -2586
rect 473866 -2822 474102 -2586
rect 477266 -4422 477502 -4186
rect 477586 -4422 477822 -4186
rect 477266 -4742 477502 -4506
rect 477586 -4742 477822 -4506
rect 462986 -7302 463222 -7066
rect 463306 -7302 463542 -7066
rect 462986 -7622 463222 -7386
rect 463306 -7622 463542 -7386
rect 491546 -3462 491782 -3226
rect 491866 -3462 492102 -3226
rect 491546 -3782 491782 -3546
rect 491866 -3782 492102 -3546
rect 495266 -5382 495502 -5146
rect 495586 -5382 495822 -5146
rect 495266 -5702 495502 -5466
rect 495586 -5702 495822 -5466
rect 480986 -6342 481222 -6106
rect 481306 -6342 481542 -6106
rect 480986 -6662 481222 -6426
rect 481306 -6662 481542 -6426
rect 509546 -2502 509782 -2266
rect 509866 -2502 510102 -2266
rect 509546 -2822 509782 -2586
rect 509866 -2822 510102 -2586
rect 513266 -4422 513502 -4186
rect 513586 -4422 513822 -4186
rect 513266 -4742 513502 -4506
rect 513586 -4742 513822 -4506
rect 498986 -7302 499222 -7066
rect 499306 -7302 499542 -7066
rect 498986 -7622 499222 -7386
rect 499306 -7622 499542 -7386
rect 527546 -3462 527782 -3226
rect 527866 -3462 528102 -3226
rect 527546 -3782 527782 -3546
rect 527866 -3782 528102 -3546
rect 531266 -5382 531502 -5146
rect 531586 -5382 531822 -5146
rect 531266 -5702 531502 -5466
rect 531586 -5702 531822 -5466
rect 516986 -6342 517222 -6106
rect 517306 -6342 517542 -6106
rect 516986 -6662 517222 -6426
rect 517306 -6662 517542 -6426
rect 545546 -2502 545782 -2266
rect 545866 -2502 546102 -2266
rect 545546 -2822 545782 -2586
rect 545866 -2822 546102 -2586
rect 549266 -4422 549502 -4186
rect 549586 -4422 549822 -4186
rect 549266 -4742 549502 -4506
rect 549586 -4742 549822 -4506
rect 534986 -7302 535222 -7066
rect 535306 -7302 535542 -7066
rect 534986 -7622 535222 -7386
rect 535306 -7622 535542 -7386
rect 563546 -3462 563782 -3226
rect 563866 -3462 564102 -3226
rect 563546 -3782 563782 -3546
rect 563866 -3782 564102 -3546
rect 567266 -5382 567502 -5146
rect 567586 -5382 567822 -5146
rect 567266 -5702 567502 -5466
rect 567586 -5702 567822 -5466
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 581546 706522 581782 706758
rect 581866 706522 582102 706758
rect 581546 706202 581782 706438
rect 581866 706202 582102 706438
rect 570986 680378 571222 680614
rect 571306 680378 571542 680614
rect 570986 680058 571222 680294
rect 571306 680058 571542 680294
rect 570986 644378 571222 644614
rect 571306 644378 571542 644614
rect 570986 644058 571222 644294
rect 571306 644058 571542 644294
rect 570986 608378 571222 608614
rect 571306 608378 571542 608614
rect 570986 608058 571222 608294
rect 571306 608058 571542 608294
rect 570986 572378 571222 572614
rect 571306 572378 571542 572614
rect 570986 572058 571222 572294
rect 571306 572058 571542 572294
rect 570986 536378 571222 536614
rect 571306 536378 571542 536614
rect 570986 536058 571222 536294
rect 571306 536058 571542 536294
rect 570986 500378 571222 500614
rect 571306 500378 571542 500614
rect 570986 500058 571222 500294
rect 571306 500058 571542 500294
rect 570986 464378 571222 464614
rect 571306 464378 571542 464614
rect 570986 464058 571222 464294
rect 571306 464058 571542 464294
rect 570986 428378 571222 428614
rect 571306 428378 571542 428614
rect 570986 428058 571222 428294
rect 571306 428058 571542 428294
rect 570986 392378 571222 392614
rect 571306 392378 571542 392614
rect 570986 392058 571222 392294
rect 571306 392058 571542 392294
rect 570986 356378 571222 356614
rect 571306 356378 571542 356614
rect 570986 356058 571222 356294
rect 571306 356058 571542 356294
rect 570986 320378 571222 320614
rect 571306 320378 571542 320614
rect 570986 320058 571222 320294
rect 571306 320058 571542 320294
rect 570986 284378 571222 284614
rect 571306 284378 571542 284614
rect 570986 284058 571222 284294
rect 571306 284058 571542 284294
rect 570986 248378 571222 248614
rect 571306 248378 571542 248614
rect 570986 248058 571222 248294
rect 571306 248058 571542 248294
rect 570986 212378 571222 212614
rect 571306 212378 571542 212614
rect 570986 212058 571222 212294
rect 571306 212058 571542 212294
rect 570986 176378 571222 176614
rect 571306 176378 571542 176614
rect 570986 176058 571222 176294
rect 571306 176058 571542 176294
rect 570986 140378 571222 140614
rect 571306 140378 571542 140614
rect 570986 140058 571222 140294
rect 571306 140058 571542 140294
rect 570986 104378 571222 104614
rect 571306 104378 571542 104614
rect 570986 104058 571222 104294
rect 571306 104058 571542 104294
rect 570986 68378 571222 68614
rect 571306 68378 571542 68614
rect 570986 68058 571222 68294
rect 571306 68058 571542 68294
rect 570986 32378 571222 32614
rect 571306 32378 571542 32614
rect 570986 32058 571222 32294
rect 571306 32058 571542 32294
rect 552986 -6342 553222 -6106
rect 553306 -6342 553542 -6106
rect 552986 -6662 553222 -6426
rect 553306 -6662 553542 -6426
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 690938 587498 691174
rect 587582 690938 587818 691174
rect 587262 690618 587498 690854
rect 587582 690618 587818 690854
rect 587262 654938 587498 655174
rect 587582 654938 587818 655174
rect 587262 654618 587498 654854
rect 587582 654618 587818 654854
rect 587262 618938 587498 619174
rect 587582 618938 587818 619174
rect 587262 618618 587498 618854
rect 587582 618618 587818 618854
rect 587262 582938 587498 583174
rect 587582 582938 587818 583174
rect 587262 582618 587498 582854
rect 587582 582618 587818 582854
rect 587262 546938 587498 547174
rect 587582 546938 587818 547174
rect 587262 546618 587498 546854
rect 587582 546618 587818 546854
rect 587262 510938 587498 511174
rect 587582 510938 587818 511174
rect 587262 510618 587498 510854
rect 587582 510618 587818 510854
rect 587262 474938 587498 475174
rect 587582 474938 587818 475174
rect 587262 474618 587498 474854
rect 587582 474618 587818 474854
rect 587262 438938 587498 439174
rect 587582 438938 587818 439174
rect 587262 438618 587498 438854
rect 587582 438618 587818 438854
rect 587262 402938 587498 403174
rect 587582 402938 587818 403174
rect 587262 402618 587498 402854
rect 587582 402618 587818 402854
rect 587262 366938 587498 367174
rect 587582 366938 587818 367174
rect 587262 366618 587498 366854
rect 587582 366618 587818 366854
rect 587262 330938 587498 331174
rect 587582 330938 587818 331174
rect 587262 330618 587498 330854
rect 587582 330618 587818 330854
rect 587262 294938 587498 295174
rect 587582 294938 587818 295174
rect 587262 294618 587498 294854
rect 587582 294618 587818 294854
rect 587262 258938 587498 259174
rect 587582 258938 587818 259174
rect 587262 258618 587498 258854
rect 587582 258618 587818 258854
rect 587262 222938 587498 223174
rect 587582 222938 587818 223174
rect 587262 222618 587498 222854
rect 587582 222618 587818 222854
rect 587262 186938 587498 187174
rect 587582 186938 587818 187174
rect 587262 186618 587498 186854
rect 587582 186618 587818 186854
rect 587262 150938 587498 151174
rect 587582 150938 587818 151174
rect 587262 150618 587498 150854
rect 587582 150618 587818 150854
rect 587262 114938 587498 115174
rect 587582 114938 587818 115174
rect 587262 114618 587498 114854
rect 587582 114618 587818 114854
rect 587262 78938 587498 79174
rect 587582 78938 587818 79174
rect 587262 78618 587498 78854
rect 587582 78618 587818 78854
rect 587262 42938 587498 43174
rect 587582 42938 587818 43174
rect 587262 42618 587498 42854
rect 587582 42618 587818 42854
rect 587262 6938 587498 7174
rect 587582 6938 587818 7174
rect 587262 6618 587498 6854
rect 587582 6618 587818 6854
rect 581546 -2502 581782 -2266
rect 581866 -2502 582102 -2266
rect 581546 -2822 581782 -2586
rect 581866 -2822 582102 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 672938 588458 673174
rect 588542 672938 588778 673174
rect 588222 672618 588458 672854
rect 588542 672618 588778 672854
rect 588222 636938 588458 637174
rect 588542 636938 588778 637174
rect 588222 636618 588458 636854
rect 588542 636618 588778 636854
rect 588222 600938 588458 601174
rect 588542 600938 588778 601174
rect 588222 600618 588458 600854
rect 588542 600618 588778 600854
rect 588222 564938 588458 565174
rect 588542 564938 588778 565174
rect 588222 564618 588458 564854
rect 588542 564618 588778 564854
rect 588222 528938 588458 529174
rect 588542 528938 588778 529174
rect 588222 528618 588458 528854
rect 588542 528618 588778 528854
rect 588222 492938 588458 493174
rect 588542 492938 588778 493174
rect 588222 492618 588458 492854
rect 588542 492618 588778 492854
rect 588222 456938 588458 457174
rect 588542 456938 588778 457174
rect 588222 456618 588458 456854
rect 588542 456618 588778 456854
rect 588222 420938 588458 421174
rect 588542 420938 588778 421174
rect 588222 420618 588458 420854
rect 588542 420618 588778 420854
rect 588222 384938 588458 385174
rect 588542 384938 588778 385174
rect 588222 384618 588458 384854
rect 588542 384618 588778 384854
rect 588222 348938 588458 349174
rect 588542 348938 588778 349174
rect 588222 348618 588458 348854
rect 588542 348618 588778 348854
rect 588222 312938 588458 313174
rect 588542 312938 588778 313174
rect 588222 312618 588458 312854
rect 588542 312618 588778 312854
rect 588222 276938 588458 277174
rect 588542 276938 588778 277174
rect 588222 276618 588458 276854
rect 588542 276618 588778 276854
rect 588222 240938 588458 241174
rect 588542 240938 588778 241174
rect 588222 240618 588458 240854
rect 588542 240618 588778 240854
rect 588222 204938 588458 205174
rect 588542 204938 588778 205174
rect 588222 204618 588458 204854
rect 588542 204618 588778 204854
rect 588222 168938 588458 169174
rect 588542 168938 588778 169174
rect 588222 168618 588458 168854
rect 588542 168618 588778 168854
rect 588222 132938 588458 133174
rect 588542 132938 588778 133174
rect 588222 132618 588458 132854
rect 588542 132618 588778 132854
rect 588222 96938 588458 97174
rect 588542 96938 588778 97174
rect 588222 96618 588458 96854
rect 588542 96618 588778 96854
rect 588222 60938 588458 61174
rect 588542 60938 588778 61174
rect 588222 60618 588458 60854
rect 588542 60618 588778 60854
rect 588222 24938 588458 25174
rect 588542 24938 588778 25174
rect 588222 24618 588458 24854
rect 588542 24618 588778 24854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 694658 589418 694894
rect 589502 694658 589738 694894
rect 589182 694338 589418 694574
rect 589502 694338 589738 694574
rect 589182 658658 589418 658894
rect 589502 658658 589738 658894
rect 589182 658338 589418 658574
rect 589502 658338 589738 658574
rect 589182 622658 589418 622894
rect 589502 622658 589738 622894
rect 589182 622338 589418 622574
rect 589502 622338 589738 622574
rect 589182 586658 589418 586894
rect 589502 586658 589738 586894
rect 589182 586338 589418 586574
rect 589502 586338 589738 586574
rect 589182 550658 589418 550894
rect 589502 550658 589738 550894
rect 589182 550338 589418 550574
rect 589502 550338 589738 550574
rect 589182 514658 589418 514894
rect 589502 514658 589738 514894
rect 589182 514338 589418 514574
rect 589502 514338 589738 514574
rect 589182 478658 589418 478894
rect 589502 478658 589738 478894
rect 589182 478338 589418 478574
rect 589502 478338 589738 478574
rect 589182 442658 589418 442894
rect 589502 442658 589738 442894
rect 589182 442338 589418 442574
rect 589502 442338 589738 442574
rect 589182 406658 589418 406894
rect 589502 406658 589738 406894
rect 589182 406338 589418 406574
rect 589502 406338 589738 406574
rect 589182 370658 589418 370894
rect 589502 370658 589738 370894
rect 589182 370338 589418 370574
rect 589502 370338 589738 370574
rect 589182 334658 589418 334894
rect 589502 334658 589738 334894
rect 589182 334338 589418 334574
rect 589502 334338 589738 334574
rect 589182 298658 589418 298894
rect 589502 298658 589738 298894
rect 589182 298338 589418 298574
rect 589502 298338 589738 298574
rect 589182 262658 589418 262894
rect 589502 262658 589738 262894
rect 589182 262338 589418 262574
rect 589502 262338 589738 262574
rect 589182 226658 589418 226894
rect 589502 226658 589738 226894
rect 589182 226338 589418 226574
rect 589502 226338 589738 226574
rect 589182 190658 589418 190894
rect 589502 190658 589738 190894
rect 589182 190338 589418 190574
rect 589502 190338 589738 190574
rect 589182 154658 589418 154894
rect 589502 154658 589738 154894
rect 589182 154338 589418 154574
rect 589502 154338 589738 154574
rect 589182 118658 589418 118894
rect 589502 118658 589738 118894
rect 589182 118338 589418 118574
rect 589502 118338 589738 118574
rect 589182 82658 589418 82894
rect 589502 82658 589738 82894
rect 589182 82338 589418 82574
rect 589502 82338 589738 82574
rect 589182 46658 589418 46894
rect 589502 46658 589738 46894
rect 589182 46338 589418 46574
rect 589502 46338 589738 46574
rect 589182 10658 589418 10894
rect 589502 10658 589738 10894
rect 589182 10338 589418 10574
rect 589502 10338 589738 10574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 676658 590378 676894
rect 590462 676658 590698 676894
rect 590142 676338 590378 676574
rect 590462 676338 590698 676574
rect 590142 640658 590378 640894
rect 590462 640658 590698 640894
rect 590142 640338 590378 640574
rect 590462 640338 590698 640574
rect 590142 604658 590378 604894
rect 590462 604658 590698 604894
rect 590142 604338 590378 604574
rect 590462 604338 590698 604574
rect 590142 568658 590378 568894
rect 590462 568658 590698 568894
rect 590142 568338 590378 568574
rect 590462 568338 590698 568574
rect 590142 532658 590378 532894
rect 590462 532658 590698 532894
rect 590142 532338 590378 532574
rect 590462 532338 590698 532574
rect 590142 496658 590378 496894
rect 590462 496658 590698 496894
rect 590142 496338 590378 496574
rect 590462 496338 590698 496574
rect 590142 460658 590378 460894
rect 590462 460658 590698 460894
rect 590142 460338 590378 460574
rect 590462 460338 590698 460574
rect 590142 424658 590378 424894
rect 590462 424658 590698 424894
rect 590142 424338 590378 424574
rect 590462 424338 590698 424574
rect 590142 388658 590378 388894
rect 590462 388658 590698 388894
rect 590142 388338 590378 388574
rect 590462 388338 590698 388574
rect 590142 352658 590378 352894
rect 590462 352658 590698 352894
rect 590142 352338 590378 352574
rect 590462 352338 590698 352574
rect 590142 316658 590378 316894
rect 590462 316658 590698 316894
rect 590142 316338 590378 316574
rect 590462 316338 590698 316574
rect 590142 280658 590378 280894
rect 590462 280658 590698 280894
rect 590142 280338 590378 280574
rect 590462 280338 590698 280574
rect 590142 244658 590378 244894
rect 590462 244658 590698 244894
rect 590142 244338 590378 244574
rect 590462 244338 590698 244574
rect 590142 208658 590378 208894
rect 590462 208658 590698 208894
rect 590142 208338 590378 208574
rect 590462 208338 590698 208574
rect 590142 172658 590378 172894
rect 590462 172658 590698 172894
rect 590142 172338 590378 172574
rect 590462 172338 590698 172574
rect 590142 136658 590378 136894
rect 590462 136658 590698 136894
rect 590142 136338 590378 136574
rect 590462 136338 590698 136574
rect 590142 100658 590378 100894
rect 590462 100658 590698 100894
rect 590142 100338 590378 100574
rect 590462 100338 590698 100574
rect 590142 64658 590378 64894
rect 590462 64658 590698 64894
rect 590142 64338 590378 64574
rect 590462 64338 590698 64574
rect 590142 28658 590378 28894
rect 590462 28658 590698 28894
rect 590142 28338 590378 28574
rect 590462 28338 590698 28574
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 698378 591338 698614
rect 591422 698378 591658 698614
rect 591102 698058 591338 698294
rect 591422 698058 591658 698294
rect 591102 662378 591338 662614
rect 591422 662378 591658 662614
rect 591102 662058 591338 662294
rect 591422 662058 591658 662294
rect 591102 626378 591338 626614
rect 591422 626378 591658 626614
rect 591102 626058 591338 626294
rect 591422 626058 591658 626294
rect 591102 590378 591338 590614
rect 591422 590378 591658 590614
rect 591102 590058 591338 590294
rect 591422 590058 591658 590294
rect 591102 554378 591338 554614
rect 591422 554378 591658 554614
rect 591102 554058 591338 554294
rect 591422 554058 591658 554294
rect 591102 518378 591338 518614
rect 591422 518378 591658 518614
rect 591102 518058 591338 518294
rect 591422 518058 591658 518294
rect 591102 482378 591338 482614
rect 591422 482378 591658 482614
rect 591102 482058 591338 482294
rect 591422 482058 591658 482294
rect 591102 446378 591338 446614
rect 591422 446378 591658 446614
rect 591102 446058 591338 446294
rect 591422 446058 591658 446294
rect 591102 410378 591338 410614
rect 591422 410378 591658 410614
rect 591102 410058 591338 410294
rect 591422 410058 591658 410294
rect 591102 374378 591338 374614
rect 591422 374378 591658 374614
rect 591102 374058 591338 374294
rect 591422 374058 591658 374294
rect 591102 338378 591338 338614
rect 591422 338378 591658 338614
rect 591102 338058 591338 338294
rect 591422 338058 591658 338294
rect 591102 302378 591338 302614
rect 591422 302378 591658 302614
rect 591102 302058 591338 302294
rect 591422 302058 591658 302294
rect 591102 266378 591338 266614
rect 591422 266378 591658 266614
rect 591102 266058 591338 266294
rect 591422 266058 591658 266294
rect 591102 230378 591338 230614
rect 591422 230378 591658 230614
rect 591102 230058 591338 230294
rect 591422 230058 591658 230294
rect 591102 194378 591338 194614
rect 591422 194378 591658 194614
rect 591102 194058 591338 194294
rect 591422 194058 591658 194294
rect 591102 158378 591338 158614
rect 591422 158378 591658 158614
rect 591102 158058 591338 158294
rect 591422 158058 591658 158294
rect 591102 122378 591338 122614
rect 591422 122378 591658 122614
rect 591102 122058 591338 122294
rect 591422 122058 591658 122294
rect 591102 86378 591338 86614
rect 591422 86378 591658 86614
rect 591102 86058 591338 86294
rect 591422 86058 591658 86294
rect 591102 50378 591338 50614
rect 591422 50378 591658 50614
rect 591102 50058 591338 50294
rect 591422 50058 591658 50294
rect 591102 14378 591338 14614
rect 591422 14378 591658 14614
rect 591102 14058 591338 14294
rect 591422 14058 591658 14294
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 680378 592298 680614
rect 592382 680378 592618 680614
rect 592062 680058 592298 680294
rect 592382 680058 592618 680294
rect 592062 644378 592298 644614
rect 592382 644378 592618 644614
rect 592062 644058 592298 644294
rect 592382 644058 592618 644294
rect 592062 608378 592298 608614
rect 592382 608378 592618 608614
rect 592062 608058 592298 608294
rect 592382 608058 592618 608294
rect 592062 572378 592298 572614
rect 592382 572378 592618 572614
rect 592062 572058 592298 572294
rect 592382 572058 592618 572294
rect 592062 536378 592298 536614
rect 592382 536378 592618 536614
rect 592062 536058 592298 536294
rect 592382 536058 592618 536294
rect 592062 500378 592298 500614
rect 592382 500378 592618 500614
rect 592062 500058 592298 500294
rect 592382 500058 592618 500294
rect 592062 464378 592298 464614
rect 592382 464378 592618 464614
rect 592062 464058 592298 464294
rect 592382 464058 592618 464294
rect 592062 428378 592298 428614
rect 592382 428378 592618 428614
rect 592062 428058 592298 428294
rect 592382 428058 592618 428294
rect 592062 392378 592298 392614
rect 592382 392378 592618 392614
rect 592062 392058 592298 392294
rect 592382 392058 592618 392294
rect 592062 356378 592298 356614
rect 592382 356378 592618 356614
rect 592062 356058 592298 356294
rect 592382 356058 592618 356294
rect 592062 320378 592298 320614
rect 592382 320378 592618 320614
rect 592062 320058 592298 320294
rect 592382 320058 592618 320294
rect 592062 284378 592298 284614
rect 592382 284378 592618 284614
rect 592062 284058 592298 284294
rect 592382 284058 592618 284294
rect 592062 248378 592298 248614
rect 592382 248378 592618 248614
rect 592062 248058 592298 248294
rect 592382 248058 592618 248294
rect 592062 212378 592298 212614
rect 592382 212378 592618 212614
rect 592062 212058 592298 212294
rect 592382 212058 592618 212294
rect 592062 176378 592298 176614
rect 592382 176378 592618 176614
rect 592062 176058 592298 176294
rect 592382 176058 592618 176294
rect 592062 140378 592298 140614
rect 592382 140378 592618 140614
rect 592062 140058 592298 140294
rect 592382 140058 592618 140294
rect 592062 104378 592298 104614
rect 592382 104378 592618 104614
rect 592062 104058 592298 104294
rect 592382 104058 592618 104294
rect 592062 68378 592298 68614
rect 592382 68378 592618 68614
rect 592062 68058 592298 68294
rect 592382 68058 592618 68294
rect 592062 32378 592298 32614
rect 592382 32378 592618 32614
rect 592062 32058 592298 32294
rect 592382 32058 592618 32294
rect 570986 -7302 571222 -7066
rect 571306 -7302 571542 -7066
rect 570986 -7622 571222 -7386
rect 571306 -7622 571542 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 592650 698294
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 590730 694894
rect -6806 694574 590730 694658
rect -6806 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 590730 694574
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 588810 691174
rect -4886 690854 588810 690938
rect -4886 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 588810 690854
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 8250 687454
rect 8486 687218 38970 687454
rect 39206 687218 69690 687454
rect 69926 687218 100410 687454
rect 100646 687218 131130 687454
rect 131366 687218 161850 687454
rect 162086 687218 192570 687454
rect 192806 687218 223290 687454
rect 223526 687218 254010 687454
rect 254246 687218 284730 687454
rect 284966 687218 315450 687454
rect 315686 687218 346170 687454
rect 346406 687218 376890 687454
rect 377126 687218 407610 687454
rect 407846 687218 438330 687454
rect 438566 687218 469050 687454
rect 469286 687218 499770 687454
rect 500006 687218 530490 687454
rect 530726 687218 561210 687454
rect 561446 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 8250 687134
rect 8486 686898 38970 687134
rect 39206 686898 69690 687134
rect 69926 686898 100410 687134
rect 100646 686898 131130 687134
rect 131366 686898 161850 687134
rect 162086 686898 192570 687134
rect 192806 686898 223290 687134
rect 223526 686898 254010 687134
rect 254246 686898 284730 687134
rect 284966 686898 315450 687134
rect 315686 686898 346170 687134
rect 346406 686898 376890 687134
rect 377126 686898 407610 687134
rect 407846 686898 438330 687134
rect 438566 686898 469050 687134
rect 469286 686898 499770 687134
rect 500006 686898 530490 687134
rect 530726 686898 561210 687134
rect 561446 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect -8726 680294 592650 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect -6806 676574 590730 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect -4886 672854 588810 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 23610 669454
rect 23846 669218 54330 669454
rect 54566 669218 85050 669454
rect 85286 669218 115770 669454
rect 116006 669218 146490 669454
rect 146726 669218 177210 669454
rect 177446 669218 207930 669454
rect 208166 669218 238650 669454
rect 238886 669218 269370 669454
rect 269606 669218 300090 669454
rect 300326 669218 330810 669454
rect 331046 669218 361530 669454
rect 361766 669218 392250 669454
rect 392486 669218 422970 669454
rect 423206 669218 453690 669454
rect 453926 669218 484410 669454
rect 484646 669218 515130 669454
rect 515366 669218 545850 669454
rect 546086 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 23610 669134
rect 23846 668898 54330 669134
rect 54566 668898 85050 669134
rect 85286 668898 115770 669134
rect 116006 668898 146490 669134
rect 146726 668898 177210 669134
rect 177446 668898 207930 669134
rect 208166 668898 238650 669134
rect 238886 668898 269370 669134
rect 269606 668898 300090 669134
rect 300326 668898 330810 669134
rect 331046 668898 361530 669134
rect 361766 668898 392250 669134
rect 392486 668898 422970 669134
rect 423206 668898 453690 669134
rect 453926 668898 484410 669134
rect 484646 668898 515130 669134
rect 515366 668898 545850 669134
rect 546086 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 592650 662294
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 590730 658894
rect -6806 658574 590730 658658
rect -6806 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 590730 658574
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 588810 655174
rect -4886 654854 588810 654938
rect -4886 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 588810 654854
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 8250 651454
rect 8486 651218 38970 651454
rect 39206 651218 69690 651454
rect 69926 651218 100410 651454
rect 100646 651218 131130 651454
rect 131366 651218 161850 651454
rect 162086 651218 192570 651454
rect 192806 651218 223290 651454
rect 223526 651218 254010 651454
rect 254246 651218 284730 651454
rect 284966 651218 315450 651454
rect 315686 651218 346170 651454
rect 346406 651218 376890 651454
rect 377126 651218 407610 651454
rect 407846 651218 438330 651454
rect 438566 651218 469050 651454
rect 469286 651218 499770 651454
rect 500006 651218 530490 651454
rect 530726 651218 561210 651454
rect 561446 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 8250 651134
rect 8486 650898 38970 651134
rect 39206 650898 69690 651134
rect 69926 650898 100410 651134
rect 100646 650898 131130 651134
rect 131366 650898 161850 651134
rect 162086 650898 192570 651134
rect 192806 650898 223290 651134
rect 223526 650898 254010 651134
rect 254246 650898 284730 651134
rect 284966 650898 315450 651134
rect 315686 650898 346170 651134
rect 346406 650898 376890 651134
rect 377126 650898 407610 651134
rect 407846 650898 438330 651134
rect 438566 650898 469050 651134
rect 469286 650898 499770 651134
rect 500006 650898 530490 651134
rect 530726 650898 561210 651134
rect 561446 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect -8726 644294 592650 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect -6806 640574 590730 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect -4886 636854 588810 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 23610 633454
rect 23846 633218 54330 633454
rect 54566 633218 85050 633454
rect 85286 633218 115770 633454
rect 116006 633218 146490 633454
rect 146726 633218 177210 633454
rect 177446 633218 207930 633454
rect 208166 633218 238650 633454
rect 238886 633218 269370 633454
rect 269606 633218 300090 633454
rect 300326 633218 330810 633454
rect 331046 633218 361530 633454
rect 361766 633218 392250 633454
rect 392486 633218 422970 633454
rect 423206 633218 453690 633454
rect 453926 633218 484410 633454
rect 484646 633218 515130 633454
rect 515366 633218 545850 633454
rect 546086 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 23610 633134
rect 23846 632898 54330 633134
rect 54566 632898 85050 633134
rect 85286 632898 115770 633134
rect 116006 632898 146490 633134
rect 146726 632898 177210 633134
rect 177446 632898 207930 633134
rect 208166 632898 238650 633134
rect 238886 632898 269370 633134
rect 269606 632898 300090 633134
rect 300326 632898 330810 633134
rect 331046 632898 361530 633134
rect 361766 632898 392250 633134
rect 392486 632898 422970 633134
rect 423206 632898 453690 633134
rect 453926 632898 484410 633134
rect 484646 632898 515130 633134
rect 515366 632898 545850 633134
rect 546086 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 592650 626294
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 590730 622894
rect -6806 622574 590730 622658
rect -6806 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 590730 622574
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 588810 619174
rect -4886 618854 588810 618938
rect -4886 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 588810 618854
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 8250 615454
rect 8486 615218 38970 615454
rect 39206 615218 69690 615454
rect 69926 615218 100410 615454
rect 100646 615218 131130 615454
rect 131366 615218 161850 615454
rect 162086 615218 192570 615454
rect 192806 615218 223290 615454
rect 223526 615218 254010 615454
rect 254246 615218 284730 615454
rect 284966 615218 315450 615454
rect 315686 615218 346170 615454
rect 346406 615218 376890 615454
rect 377126 615218 407610 615454
rect 407846 615218 438330 615454
rect 438566 615218 469050 615454
rect 469286 615218 499770 615454
rect 500006 615218 530490 615454
rect 530726 615218 561210 615454
rect 561446 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 8250 615134
rect 8486 614898 38970 615134
rect 39206 614898 69690 615134
rect 69926 614898 100410 615134
rect 100646 614898 131130 615134
rect 131366 614898 161850 615134
rect 162086 614898 192570 615134
rect 192806 614898 223290 615134
rect 223526 614898 254010 615134
rect 254246 614898 284730 615134
rect 284966 614898 315450 615134
rect 315686 614898 346170 615134
rect 346406 614898 376890 615134
rect 377126 614898 407610 615134
rect 407846 614898 438330 615134
rect 438566 614898 469050 615134
rect 469286 614898 499770 615134
rect 500006 614898 530490 615134
rect 530726 614898 561210 615134
rect 561446 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect -8726 608294 592650 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect -6806 604574 590730 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect -4886 600854 588810 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 23610 597454
rect 23846 597218 54330 597454
rect 54566 597218 85050 597454
rect 85286 597218 115770 597454
rect 116006 597218 146490 597454
rect 146726 597218 177210 597454
rect 177446 597218 207930 597454
rect 208166 597218 238650 597454
rect 238886 597218 269370 597454
rect 269606 597218 300090 597454
rect 300326 597218 330810 597454
rect 331046 597218 361530 597454
rect 361766 597218 392250 597454
rect 392486 597218 422970 597454
rect 423206 597218 453690 597454
rect 453926 597218 484410 597454
rect 484646 597218 515130 597454
rect 515366 597218 545850 597454
rect 546086 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 23610 597134
rect 23846 596898 54330 597134
rect 54566 596898 85050 597134
rect 85286 596898 115770 597134
rect 116006 596898 146490 597134
rect 146726 596898 177210 597134
rect 177446 596898 207930 597134
rect 208166 596898 238650 597134
rect 238886 596898 269370 597134
rect 269606 596898 300090 597134
rect 300326 596898 330810 597134
rect 331046 596898 361530 597134
rect 361766 596898 392250 597134
rect 392486 596898 422970 597134
rect 423206 596898 453690 597134
rect 453926 596898 484410 597134
rect 484646 596898 515130 597134
rect 515366 596898 545850 597134
rect 546086 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 592650 590294
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 590730 586894
rect -6806 586574 590730 586658
rect -6806 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 590730 586574
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 588810 583174
rect -4886 582854 588810 582938
rect -4886 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 588810 582854
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 8250 579454
rect 8486 579218 38970 579454
rect 39206 579218 69690 579454
rect 69926 579218 100410 579454
rect 100646 579218 131130 579454
rect 131366 579218 161850 579454
rect 162086 579218 192570 579454
rect 192806 579218 223290 579454
rect 223526 579218 254010 579454
rect 254246 579218 284730 579454
rect 284966 579218 315450 579454
rect 315686 579218 346170 579454
rect 346406 579218 376890 579454
rect 377126 579218 407610 579454
rect 407846 579218 438330 579454
rect 438566 579218 469050 579454
rect 469286 579218 499770 579454
rect 500006 579218 530490 579454
rect 530726 579218 561210 579454
rect 561446 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 8250 579134
rect 8486 578898 38970 579134
rect 39206 578898 69690 579134
rect 69926 578898 100410 579134
rect 100646 578898 131130 579134
rect 131366 578898 161850 579134
rect 162086 578898 192570 579134
rect 192806 578898 223290 579134
rect 223526 578898 254010 579134
rect 254246 578898 284730 579134
rect 284966 578898 315450 579134
rect 315686 578898 346170 579134
rect 346406 578898 376890 579134
rect 377126 578898 407610 579134
rect 407846 578898 438330 579134
rect 438566 578898 469050 579134
rect 469286 578898 499770 579134
rect 500006 578898 530490 579134
rect 530726 578898 561210 579134
rect 561446 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect -8726 572294 592650 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect -6806 568574 590730 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect -4886 564854 588810 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect -4886 564586 588810 564618
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 23610 561454
rect 23846 561218 54330 561454
rect 54566 561218 85050 561454
rect 85286 561218 115770 561454
rect 116006 561218 146490 561454
rect 146726 561218 177210 561454
rect 177446 561218 207930 561454
rect 208166 561218 238650 561454
rect 238886 561218 269370 561454
rect 269606 561218 300090 561454
rect 300326 561218 330810 561454
rect 331046 561218 361530 561454
rect 361766 561218 392250 561454
rect 392486 561218 422970 561454
rect 423206 561218 453690 561454
rect 453926 561218 484410 561454
rect 484646 561218 515130 561454
rect 515366 561218 545850 561454
rect 546086 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 23610 561134
rect 23846 560898 54330 561134
rect 54566 560898 85050 561134
rect 85286 560898 115770 561134
rect 116006 560898 146490 561134
rect 146726 560898 177210 561134
rect 177446 560898 207930 561134
rect 208166 560898 238650 561134
rect 238886 560898 269370 561134
rect 269606 560898 300090 561134
rect 300326 560898 330810 561134
rect 331046 560898 361530 561134
rect 361766 560898 392250 561134
rect 392486 560898 422970 561134
rect 423206 560898 453690 561134
rect 453926 560898 484410 561134
rect 484646 560898 515130 561134
rect 515366 560898 545850 561134
rect 546086 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 592650 554294
rect -8726 554026 592650 554058
rect -6806 550894 590730 550926
rect -6806 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 590730 550894
rect -6806 550574 590730 550658
rect -6806 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 590730 550574
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 588810 547174
rect -4886 546854 588810 546938
rect -4886 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 588810 546854
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 8250 543454
rect 8486 543218 38970 543454
rect 39206 543218 69690 543454
rect 69926 543218 100410 543454
rect 100646 543218 131130 543454
rect 131366 543218 161850 543454
rect 162086 543218 192570 543454
rect 192806 543218 223290 543454
rect 223526 543218 254010 543454
rect 254246 543218 284730 543454
rect 284966 543218 315450 543454
rect 315686 543218 346170 543454
rect 346406 543218 376890 543454
rect 377126 543218 407610 543454
rect 407846 543218 438330 543454
rect 438566 543218 469050 543454
rect 469286 543218 499770 543454
rect 500006 543218 530490 543454
rect 530726 543218 561210 543454
rect 561446 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 8250 543134
rect 8486 542898 38970 543134
rect 39206 542898 69690 543134
rect 69926 542898 100410 543134
rect 100646 542898 131130 543134
rect 131366 542898 161850 543134
rect 162086 542898 192570 543134
rect 192806 542898 223290 543134
rect 223526 542898 254010 543134
rect 254246 542898 284730 543134
rect 284966 542898 315450 543134
rect 315686 542898 346170 543134
rect 346406 542898 376890 543134
rect 377126 542898 407610 543134
rect 407846 542898 438330 543134
rect 438566 542898 469050 543134
rect 469286 542898 499770 543134
rect 500006 542898 530490 543134
rect 530726 542898 561210 543134
rect 561446 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect -8726 536294 592650 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect -6806 532574 590730 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect -4886 528854 588810 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 23610 525454
rect 23846 525218 54330 525454
rect 54566 525218 85050 525454
rect 85286 525218 115770 525454
rect 116006 525218 146490 525454
rect 146726 525218 177210 525454
rect 177446 525218 207930 525454
rect 208166 525218 238650 525454
rect 238886 525218 269370 525454
rect 269606 525218 300090 525454
rect 300326 525218 330810 525454
rect 331046 525218 361530 525454
rect 361766 525218 392250 525454
rect 392486 525218 422970 525454
rect 423206 525218 453690 525454
rect 453926 525218 484410 525454
rect 484646 525218 515130 525454
rect 515366 525218 545850 525454
rect 546086 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 23610 525134
rect 23846 524898 54330 525134
rect 54566 524898 85050 525134
rect 85286 524898 115770 525134
rect 116006 524898 146490 525134
rect 146726 524898 177210 525134
rect 177446 524898 207930 525134
rect 208166 524898 238650 525134
rect 238886 524898 269370 525134
rect 269606 524898 300090 525134
rect 300326 524898 330810 525134
rect 331046 524898 361530 525134
rect 361766 524898 392250 525134
rect 392486 524898 422970 525134
rect 423206 524898 453690 525134
rect 453926 524898 484410 525134
rect 484646 524898 515130 525134
rect 515366 524898 545850 525134
rect 546086 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 592650 518294
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 590730 514894
rect -6806 514574 590730 514658
rect -6806 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 590730 514574
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 588810 511174
rect -4886 510854 588810 510938
rect -4886 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 588810 510854
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 8250 507454
rect 8486 507218 38970 507454
rect 39206 507218 69690 507454
rect 69926 507218 100410 507454
rect 100646 507218 131130 507454
rect 131366 507218 161850 507454
rect 162086 507218 192570 507454
rect 192806 507218 223290 507454
rect 223526 507218 254010 507454
rect 254246 507218 284730 507454
rect 284966 507218 315450 507454
rect 315686 507218 346170 507454
rect 346406 507218 376890 507454
rect 377126 507218 407610 507454
rect 407846 507218 438330 507454
rect 438566 507218 469050 507454
rect 469286 507218 499770 507454
rect 500006 507218 530490 507454
rect 530726 507218 561210 507454
rect 561446 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 8250 507134
rect 8486 506898 38970 507134
rect 39206 506898 69690 507134
rect 69926 506898 100410 507134
rect 100646 506898 131130 507134
rect 131366 506898 161850 507134
rect 162086 506898 192570 507134
rect 192806 506898 223290 507134
rect 223526 506898 254010 507134
rect 254246 506898 284730 507134
rect 284966 506898 315450 507134
rect 315686 506898 346170 507134
rect 346406 506898 376890 507134
rect 377126 506898 407610 507134
rect 407846 506898 438330 507134
rect 438566 506898 469050 507134
rect 469286 506898 499770 507134
rect 500006 506898 530490 507134
rect 530726 506898 561210 507134
rect 561446 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect -8726 500294 592650 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect -6806 496574 590730 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect -4886 492854 588810 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 23610 489454
rect 23846 489218 54330 489454
rect 54566 489218 85050 489454
rect 85286 489218 115770 489454
rect 116006 489218 146490 489454
rect 146726 489218 177210 489454
rect 177446 489218 207930 489454
rect 208166 489218 238650 489454
rect 238886 489218 269370 489454
rect 269606 489218 300090 489454
rect 300326 489218 330810 489454
rect 331046 489218 361530 489454
rect 361766 489218 392250 489454
rect 392486 489218 422970 489454
rect 423206 489218 453690 489454
rect 453926 489218 484410 489454
rect 484646 489218 515130 489454
rect 515366 489218 545850 489454
rect 546086 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 23610 489134
rect 23846 488898 54330 489134
rect 54566 488898 85050 489134
rect 85286 488898 115770 489134
rect 116006 488898 146490 489134
rect 146726 488898 177210 489134
rect 177446 488898 207930 489134
rect 208166 488898 238650 489134
rect 238886 488898 269370 489134
rect 269606 488898 300090 489134
rect 300326 488898 330810 489134
rect 331046 488898 361530 489134
rect 361766 488898 392250 489134
rect 392486 488898 422970 489134
rect 423206 488898 453690 489134
rect 453926 488898 484410 489134
rect 484646 488898 515130 489134
rect 515366 488898 545850 489134
rect 546086 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 592650 482294
rect -8726 482026 592650 482058
rect -6806 478894 590730 478926
rect -6806 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 590730 478894
rect -6806 478574 590730 478658
rect -6806 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 590730 478574
rect -6806 478306 590730 478338
rect -4886 475174 588810 475206
rect -4886 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 588810 475174
rect -4886 474854 588810 474938
rect -4886 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 588810 474854
rect -4886 474586 588810 474618
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 8250 471454
rect 8486 471218 38970 471454
rect 39206 471218 69690 471454
rect 69926 471218 100410 471454
rect 100646 471218 131130 471454
rect 131366 471218 161850 471454
rect 162086 471218 192570 471454
rect 192806 471218 223290 471454
rect 223526 471218 254010 471454
rect 254246 471218 284730 471454
rect 284966 471218 315450 471454
rect 315686 471218 346170 471454
rect 346406 471218 376890 471454
rect 377126 471218 407610 471454
rect 407846 471218 438330 471454
rect 438566 471218 469050 471454
rect 469286 471218 499770 471454
rect 500006 471218 530490 471454
rect 530726 471218 561210 471454
rect 561446 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 8250 471134
rect 8486 470898 38970 471134
rect 39206 470898 69690 471134
rect 69926 470898 100410 471134
rect 100646 470898 131130 471134
rect 131366 470898 161850 471134
rect 162086 470898 192570 471134
rect 192806 470898 223290 471134
rect 223526 470898 254010 471134
rect 254246 470898 284730 471134
rect 284966 470898 315450 471134
rect 315686 470898 346170 471134
rect 346406 470898 376890 471134
rect 377126 470898 407610 471134
rect 407846 470898 438330 471134
rect 438566 470898 469050 471134
rect 469286 470898 499770 471134
rect 500006 470898 530490 471134
rect 530726 470898 561210 471134
rect 561446 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect -8726 464294 592650 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect -6806 460574 590730 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect -4886 456854 588810 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 23610 453454
rect 23846 453218 54330 453454
rect 54566 453218 85050 453454
rect 85286 453218 115770 453454
rect 116006 453218 146490 453454
rect 146726 453218 177210 453454
rect 177446 453218 207930 453454
rect 208166 453218 238650 453454
rect 238886 453218 269370 453454
rect 269606 453218 300090 453454
rect 300326 453218 330810 453454
rect 331046 453218 361530 453454
rect 361766 453218 392250 453454
rect 392486 453218 422970 453454
rect 423206 453218 453690 453454
rect 453926 453218 484410 453454
rect 484646 453218 515130 453454
rect 515366 453218 545850 453454
rect 546086 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 23610 453134
rect 23846 452898 54330 453134
rect 54566 452898 85050 453134
rect 85286 452898 115770 453134
rect 116006 452898 146490 453134
rect 146726 452898 177210 453134
rect 177446 452898 207930 453134
rect 208166 452898 238650 453134
rect 238886 452898 269370 453134
rect 269606 452898 300090 453134
rect 300326 452898 330810 453134
rect 331046 452898 361530 453134
rect 361766 452898 392250 453134
rect 392486 452898 422970 453134
rect 423206 452898 453690 453134
rect 453926 452898 484410 453134
rect 484646 452898 515130 453134
rect 515366 452898 545850 453134
rect 546086 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 592650 446294
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 590730 442894
rect -6806 442574 590730 442658
rect -6806 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 590730 442574
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 588810 439174
rect -4886 438854 588810 438938
rect -4886 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 588810 438854
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 8250 435454
rect 8486 435218 38970 435454
rect 39206 435218 69690 435454
rect 69926 435218 100410 435454
rect 100646 435218 131130 435454
rect 131366 435218 161850 435454
rect 162086 435218 192570 435454
rect 192806 435218 223290 435454
rect 223526 435218 254010 435454
rect 254246 435218 284730 435454
rect 284966 435218 315450 435454
rect 315686 435218 346170 435454
rect 346406 435218 376890 435454
rect 377126 435218 407610 435454
rect 407846 435218 438330 435454
rect 438566 435218 469050 435454
rect 469286 435218 499770 435454
rect 500006 435218 530490 435454
rect 530726 435218 561210 435454
rect 561446 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 8250 435134
rect 8486 434898 38970 435134
rect 39206 434898 69690 435134
rect 69926 434898 100410 435134
rect 100646 434898 131130 435134
rect 131366 434898 161850 435134
rect 162086 434898 192570 435134
rect 192806 434898 223290 435134
rect 223526 434898 254010 435134
rect 254246 434898 284730 435134
rect 284966 434898 315450 435134
rect 315686 434898 346170 435134
rect 346406 434898 376890 435134
rect 377126 434898 407610 435134
rect 407846 434898 438330 435134
rect 438566 434898 469050 435134
rect 469286 434898 499770 435134
rect 500006 434898 530490 435134
rect 530726 434898 561210 435134
rect 561446 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect -8726 428294 592650 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect -6806 424574 590730 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect -4886 420854 588810 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 23610 417454
rect 23846 417218 54330 417454
rect 54566 417218 85050 417454
rect 85286 417218 115770 417454
rect 116006 417218 146490 417454
rect 146726 417218 177210 417454
rect 177446 417218 207930 417454
rect 208166 417218 238650 417454
rect 238886 417218 269370 417454
rect 269606 417218 300090 417454
rect 300326 417218 330810 417454
rect 331046 417218 361530 417454
rect 361766 417218 392250 417454
rect 392486 417218 422970 417454
rect 423206 417218 453690 417454
rect 453926 417218 484410 417454
rect 484646 417218 515130 417454
rect 515366 417218 545850 417454
rect 546086 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 23610 417134
rect 23846 416898 54330 417134
rect 54566 416898 85050 417134
rect 85286 416898 115770 417134
rect 116006 416898 146490 417134
rect 146726 416898 177210 417134
rect 177446 416898 207930 417134
rect 208166 416898 238650 417134
rect 238886 416898 269370 417134
rect 269606 416898 300090 417134
rect 300326 416898 330810 417134
rect 331046 416898 361530 417134
rect 361766 416898 392250 417134
rect 392486 416898 422970 417134
rect 423206 416898 453690 417134
rect 453926 416898 484410 417134
rect 484646 416898 515130 417134
rect 515366 416898 545850 417134
rect 546086 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 592650 410294
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 590730 406894
rect -6806 406574 590730 406658
rect -6806 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 590730 406574
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 588810 403174
rect -4886 402854 588810 402938
rect -4886 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 588810 402854
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 8250 399454
rect 8486 399218 38970 399454
rect 39206 399218 69690 399454
rect 69926 399218 100410 399454
rect 100646 399218 131130 399454
rect 131366 399218 161850 399454
rect 162086 399218 192570 399454
rect 192806 399218 223290 399454
rect 223526 399218 254010 399454
rect 254246 399218 284730 399454
rect 284966 399218 315450 399454
rect 315686 399218 346170 399454
rect 346406 399218 376890 399454
rect 377126 399218 407610 399454
rect 407846 399218 438330 399454
rect 438566 399218 469050 399454
rect 469286 399218 499770 399454
rect 500006 399218 530490 399454
rect 530726 399218 561210 399454
rect 561446 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 8250 399134
rect 8486 398898 38970 399134
rect 39206 398898 69690 399134
rect 69926 398898 100410 399134
rect 100646 398898 131130 399134
rect 131366 398898 161850 399134
rect 162086 398898 192570 399134
rect 192806 398898 223290 399134
rect 223526 398898 254010 399134
rect 254246 398898 284730 399134
rect 284966 398898 315450 399134
rect 315686 398898 346170 399134
rect 346406 398898 376890 399134
rect 377126 398898 407610 399134
rect 407846 398898 438330 399134
rect 438566 398898 469050 399134
rect 469286 398898 499770 399134
rect 500006 398898 530490 399134
rect 530726 398898 561210 399134
rect 561446 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect -8726 392294 592650 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect -8726 392026 592650 392058
rect -6806 388894 590730 388926
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect -6806 388574 590730 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect -4886 384854 588810 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 23610 381454
rect 23846 381218 54330 381454
rect 54566 381218 85050 381454
rect 85286 381218 115770 381454
rect 116006 381218 146490 381454
rect 146726 381218 177210 381454
rect 177446 381218 207930 381454
rect 208166 381218 238650 381454
rect 238886 381218 269370 381454
rect 269606 381218 300090 381454
rect 300326 381218 330810 381454
rect 331046 381218 361530 381454
rect 361766 381218 392250 381454
rect 392486 381218 422970 381454
rect 423206 381218 453690 381454
rect 453926 381218 484410 381454
rect 484646 381218 515130 381454
rect 515366 381218 545850 381454
rect 546086 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect -2966 381134 586890 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 23610 381134
rect 23846 380898 54330 381134
rect 54566 380898 85050 381134
rect 85286 380898 115770 381134
rect 116006 380898 146490 381134
rect 146726 380898 177210 381134
rect 177446 380898 207930 381134
rect 208166 380898 238650 381134
rect 238886 380898 269370 381134
rect 269606 380898 300090 381134
rect 300326 380898 330810 381134
rect 331046 380898 361530 381134
rect 361766 380898 392250 381134
rect 392486 380898 422970 381134
rect 423206 380898 453690 381134
rect 453926 380898 484410 381134
rect 484646 380898 515130 381134
rect 515366 380898 545850 381134
rect 546086 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 592650 374294
rect -8726 374026 592650 374058
rect -6806 370894 590730 370926
rect -6806 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 590730 370894
rect -6806 370574 590730 370658
rect -6806 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 590730 370574
rect -6806 370306 590730 370338
rect -4886 367174 588810 367206
rect -4886 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 588810 367174
rect -4886 366854 588810 366938
rect -4886 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 588810 366854
rect -4886 366586 588810 366618
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 8250 363454
rect 8486 363218 38970 363454
rect 39206 363218 69690 363454
rect 69926 363218 100410 363454
rect 100646 363218 131130 363454
rect 131366 363218 161850 363454
rect 162086 363218 192570 363454
rect 192806 363218 223290 363454
rect 223526 363218 254010 363454
rect 254246 363218 284730 363454
rect 284966 363218 315450 363454
rect 315686 363218 346170 363454
rect 346406 363218 376890 363454
rect 377126 363218 407610 363454
rect 407846 363218 438330 363454
rect 438566 363218 469050 363454
rect 469286 363218 499770 363454
rect 500006 363218 530490 363454
rect 530726 363218 561210 363454
rect 561446 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 8250 363134
rect 8486 362898 38970 363134
rect 39206 362898 69690 363134
rect 69926 362898 100410 363134
rect 100646 362898 131130 363134
rect 131366 362898 161850 363134
rect 162086 362898 192570 363134
rect 192806 362898 223290 363134
rect 223526 362898 254010 363134
rect 254246 362898 284730 363134
rect 284966 362898 315450 363134
rect 315686 362898 346170 363134
rect 346406 362898 376890 363134
rect 377126 362898 407610 363134
rect 407846 362898 438330 363134
rect 438566 362898 469050 363134
rect 469286 362898 499770 363134
rect 500006 362898 530490 363134
rect 530726 362898 561210 363134
rect 561446 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect -8726 356614 592650 356646
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect -8726 356294 592650 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect -6806 352574 590730 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect -4886 348854 588810 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect -4886 348586 588810 348618
rect -2966 345454 586890 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 23610 345454
rect 23846 345218 54330 345454
rect 54566 345218 85050 345454
rect 85286 345218 115770 345454
rect 116006 345218 146490 345454
rect 146726 345218 177210 345454
rect 177446 345218 207930 345454
rect 208166 345218 238650 345454
rect 238886 345218 269370 345454
rect 269606 345218 300090 345454
rect 300326 345218 330810 345454
rect 331046 345218 361530 345454
rect 361766 345218 392250 345454
rect 392486 345218 422970 345454
rect 423206 345218 453690 345454
rect 453926 345218 484410 345454
rect 484646 345218 515130 345454
rect 515366 345218 545850 345454
rect 546086 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect -2966 345134 586890 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 23610 345134
rect 23846 344898 54330 345134
rect 54566 344898 85050 345134
rect 85286 344898 115770 345134
rect 116006 344898 146490 345134
rect 146726 344898 177210 345134
rect 177446 344898 207930 345134
rect 208166 344898 238650 345134
rect 238886 344898 269370 345134
rect 269606 344898 300090 345134
rect 300326 344898 330810 345134
rect 331046 344898 361530 345134
rect 361766 344898 392250 345134
rect 392486 344898 422970 345134
rect 423206 344898 453690 345134
rect 453926 344898 484410 345134
rect 484646 344898 515130 345134
rect 515366 344898 545850 345134
rect 546086 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect -2966 344866 586890 344898
rect -8726 338614 592650 338646
rect -8726 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 592650 338294
rect -8726 338026 592650 338058
rect -6806 334894 590730 334926
rect -6806 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 590730 334894
rect -6806 334574 590730 334658
rect -6806 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 590730 334574
rect -6806 334306 590730 334338
rect -4886 331174 588810 331206
rect -4886 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 588810 331174
rect -4886 330854 588810 330938
rect -4886 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 588810 330854
rect -4886 330586 588810 330618
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 8250 327454
rect 8486 327218 38970 327454
rect 39206 327218 69690 327454
rect 69926 327218 100410 327454
rect 100646 327218 131130 327454
rect 131366 327218 161850 327454
rect 162086 327218 192570 327454
rect 192806 327218 223290 327454
rect 223526 327218 254010 327454
rect 254246 327218 284730 327454
rect 284966 327218 315450 327454
rect 315686 327218 346170 327454
rect 346406 327218 376890 327454
rect 377126 327218 407610 327454
rect 407846 327218 438330 327454
rect 438566 327218 469050 327454
rect 469286 327218 499770 327454
rect 500006 327218 530490 327454
rect 530726 327218 561210 327454
rect 561446 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 8250 327134
rect 8486 326898 38970 327134
rect 39206 326898 69690 327134
rect 69926 326898 100410 327134
rect 100646 326898 131130 327134
rect 131366 326898 161850 327134
rect 162086 326898 192570 327134
rect 192806 326898 223290 327134
rect 223526 326898 254010 327134
rect 254246 326898 284730 327134
rect 284966 326898 315450 327134
rect 315686 326898 346170 327134
rect 346406 326898 376890 327134
rect 377126 326898 407610 327134
rect 407846 326898 438330 327134
rect 438566 326898 469050 327134
rect 469286 326898 499770 327134
rect 500006 326898 530490 327134
rect 530726 326898 561210 327134
rect 561446 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect -8726 320294 592650 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect -6806 316574 590730 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect -4886 312854 588810 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 23610 309454
rect 23846 309218 54330 309454
rect 54566 309218 85050 309454
rect 85286 309218 115770 309454
rect 116006 309218 146490 309454
rect 146726 309218 177210 309454
rect 177446 309218 207930 309454
rect 208166 309218 238650 309454
rect 238886 309218 269370 309454
rect 269606 309218 300090 309454
rect 300326 309218 330810 309454
rect 331046 309218 361530 309454
rect 361766 309218 392250 309454
rect 392486 309218 422970 309454
rect 423206 309218 453690 309454
rect 453926 309218 484410 309454
rect 484646 309218 515130 309454
rect 515366 309218 545850 309454
rect 546086 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect -2966 309134 586890 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 23610 309134
rect 23846 308898 54330 309134
rect 54566 308898 85050 309134
rect 85286 308898 115770 309134
rect 116006 308898 146490 309134
rect 146726 308898 177210 309134
rect 177446 308898 207930 309134
rect 208166 308898 238650 309134
rect 238886 308898 269370 309134
rect 269606 308898 300090 309134
rect 300326 308898 330810 309134
rect 331046 308898 361530 309134
rect 361766 308898 392250 309134
rect 392486 308898 422970 309134
rect 423206 308898 453690 309134
rect 453926 308898 484410 309134
rect 484646 308898 515130 309134
rect 515366 308898 545850 309134
rect 546086 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect -2966 308866 586890 308898
rect -8726 302614 592650 302646
rect -8726 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 592650 302294
rect -8726 302026 592650 302058
rect -6806 298894 590730 298926
rect -6806 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 590730 298894
rect -6806 298574 590730 298658
rect -6806 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 590730 298574
rect -6806 298306 590730 298338
rect -4886 295174 588810 295206
rect -4886 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 588810 295174
rect -4886 294854 588810 294938
rect -4886 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 588810 294854
rect -4886 294586 588810 294618
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 8250 291454
rect 8486 291218 38970 291454
rect 39206 291218 69690 291454
rect 69926 291218 100410 291454
rect 100646 291218 131130 291454
rect 131366 291218 161850 291454
rect 162086 291218 192570 291454
rect 192806 291218 223290 291454
rect 223526 291218 254010 291454
rect 254246 291218 284730 291454
rect 284966 291218 315450 291454
rect 315686 291218 346170 291454
rect 346406 291218 376890 291454
rect 377126 291218 407610 291454
rect 407846 291218 438330 291454
rect 438566 291218 469050 291454
rect 469286 291218 499770 291454
rect 500006 291218 530490 291454
rect 530726 291218 561210 291454
rect 561446 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 8250 291134
rect 8486 290898 38970 291134
rect 39206 290898 69690 291134
rect 69926 290898 100410 291134
rect 100646 290898 131130 291134
rect 131366 290898 161850 291134
rect 162086 290898 192570 291134
rect 192806 290898 223290 291134
rect 223526 290898 254010 291134
rect 254246 290898 284730 291134
rect 284966 290898 315450 291134
rect 315686 290898 346170 291134
rect 346406 290898 376890 291134
rect 377126 290898 407610 291134
rect 407846 290898 438330 291134
rect 438566 290898 469050 291134
rect 469286 290898 499770 291134
rect 500006 290898 530490 291134
rect 530726 290898 561210 291134
rect 561446 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect -8726 284294 592650 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect -6806 280574 590730 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect -4886 276854 588810 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect -4886 276586 588810 276618
rect -2966 273454 586890 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 23610 273454
rect 23846 273218 54330 273454
rect 54566 273218 85050 273454
rect 85286 273218 115770 273454
rect 116006 273218 146490 273454
rect 146726 273218 177210 273454
rect 177446 273218 207930 273454
rect 208166 273218 238650 273454
rect 238886 273218 269370 273454
rect 269606 273218 300090 273454
rect 300326 273218 330810 273454
rect 331046 273218 361530 273454
rect 361766 273218 392250 273454
rect 392486 273218 422970 273454
rect 423206 273218 453690 273454
rect 453926 273218 484410 273454
rect 484646 273218 515130 273454
rect 515366 273218 545850 273454
rect 546086 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect -2966 273134 586890 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 23610 273134
rect 23846 272898 54330 273134
rect 54566 272898 85050 273134
rect 85286 272898 115770 273134
rect 116006 272898 146490 273134
rect 146726 272898 177210 273134
rect 177446 272898 207930 273134
rect 208166 272898 238650 273134
rect 238886 272898 269370 273134
rect 269606 272898 300090 273134
rect 300326 272898 330810 273134
rect 331046 272898 361530 273134
rect 361766 272898 392250 273134
rect 392486 272898 422970 273134
rect 423206 272898 453690 273134
rect 453926 272898 484410 273134
rect 484646 272898 515130 273134
rect 515366 272898 545850 273134
rect 546086 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 592650 266294
rect -8726 266026 592650 266058
rect -6806 262894 590730 262926
rect -6806 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 590730 262894
rect -6806 262574 590730 262658
rect -6806 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 590730 262574
rect -6806 262306 590730 262338
rect -4886 259174 588810 259206
rect -4886 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 588810 259174
rect -4886 258854 588810 258938
rect -4886 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 588810 258854
rect -4886 258586 588810 258618
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 8250 255454
rect 8486 255218 38970 255454
rect 39206 255218 69690 255454
rect 69926 255218 100410 255454
rect 100646 255218 131130 255454
rect 131366 255218 161850 255454
rect 162086 255218 192570 255454
rect 192806 255218 223290 255454
rect 223526 255218 254010 255454
rect 254246 255218 284730 255454
rect 284966 255218 315450 255454
rect 315686 255218 346170 255454
rect 346406 255218 376890 255454
rect 377126 255218 407610 255454
rect 407846 255218 438330 255454
rect 438566 255218 469050 255454
rect 469286 255218 499770 255454
rect 500006 255218 530490 255454
rect 530726 255218 561210 255454
rect 561446 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 8250 255134
rect 8486 254898 38970 255134
rect 39206 254898 69690 255134
rect 69926 254898 100410 255134
rect 100646 254898 131130 255134
rect 131366 254898 161850 255134
rect 162086 254898 192570 255134
rect 192806 254898 223290 255134
rect 223526 254898 254010 255134
rect 254246 254898 284730 255134
rect 284966 254898 315450 255134
rect 315686 254898 346170 255134
rect 346406 254898 376890 255134
rect 377126 254898 407610 255134
rect 407846 254898 438330 255134
rect 438566 254898 469050 255134
rect 469286 254898 499770 255134
rect 500006 254898 530490 255134
rect 530726 254898 561210 255134
rect 561446 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -8726 248614 592650 248646
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect -8726 248294 592650 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect -6806 244574 590730 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect -4886 240854 588810 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 23610 237454
rect 23846 237218 54330 237454
rect 54566 237218 85050 237454
rect 85286 237218 115770 237454
rect 116006 237218 146490 237454
rect 146726 237218 177210 237454
rect 177446 237218 207930 237454
rect 208166 237218 238650 237454
rect 238886 237218 269370 237454
rect 269606 237218 300090 237454
rect 300326 237218 330810 237454
rect 331046 237218 361530 237454
rect 361766 237218 392250 237454
rect 392486 237218 422970 237454
rect 423206 237218 453690 237454
rect 453926 237218 484410 237454
rect 484646 237218 515130 237454
rect 515366 237218 545850 237454
rect 546086 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect -2966 237134 586890 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 23610 237134
rect 23846 236898 54330 237134
rect 54566 236898 85050 237134
rect 85286 236898 115770 237134
rect 116006 236898 146490 237134
rect 146726 236898 177210 237134
rect 177446 236898 207930 237134
rect 208166 236898 238650 237134
rect 238886 236898 269370 237134
rect 269606 236898 300090 237134
rect 300326 236898 330810 237134
rect 331046 236898 361530 237134
rect 361766 236898 392250 237134
rect 392486 236898 422970 237134
rect 423206 236898 453690 237134
rect 453926 236898 484410 237134
rect 484646 236898 515130 237134
rect 515366 236898 545850 237134
rect 546086 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 592650 230294
rect -8726 230026 592650 230058
rect -6806 226894 590730 226926
rect -6806 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 590730 226894
rect -6806 226574 590730 226658
rect -6806 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 590730 226574
rect -6806 226306 590730 226338
rect -4886 223174 588810 223206
rect -4886 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 588810 223174
rect -4886 222854 588810 222938
rect -4886 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 588810 222854
rect -4886 222586 588810 222618
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 8250 219454
rect 8486 219218 38970 219454
rect 39206 219218 69690 219454
rect 69926 219218 100410 219454
rect 100646 219218 131130 219454
rect 131366 219218 161850 219454
rect 162086 219218 192570 219454
rect 192806 219218 223290 219454
rect 223526 219218 254010 219454
rect 254246 219218 284730 219454
rect 284966 219218 315450 219454
rect 315686 219218 346170 219454
rect 346406 219218 376890 219454
rect 377126 219218 407610 219454
rect 407846 219218 438330 219454
rect 438566 219218 469050 219454
rect 469286 219218 499770 219454
rect 500006 219218 530490 219454
rect 530726 219218 561210 219454
rect 561446 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 8250 219134
rect 8486 218898 38970 219134
rect 39206 218898 69690 219134
rect 69926 218898 100410 219134
rect 100646 218898 131130 219134
rect 131366 218898 161850 219134
rect 162086 218898 192570 219134
rect 192806 218898 223290 219134
rect 223526 218898 254010 219134
rect 254246 218898 284730 219134
rect 284966 218898 315450 219134
rect 315686 218898 346170 219134
rect 346406 218898 376890 219134
rect 377126 218898 407610 219134
rect 407846 218898 438330 219134
rect 438566 218898 469050 219134
rect 469286 218898 499770 219134
rect 500006 218898 530490 219134
rect 530726 218898 561210 219134
rect 561446 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -8726 212614 592650 212646
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect -8726 212294 592650 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect -6806 208574 590730 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect -4886 204854 588810 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 23610 201454
rect 23846 201218 54330 201454
rect 54566 201218 85050 201454
rect 85286 201218 115770 201454
rect 116006 201218 146490 201454
rect 146726 201218 177210 201454
rect 177446 201218 207930 201454
rect 208166 201218 238650 201454
rect 238886 201218 269370 201454
rect 269606 201218 300090 201454
rect 300326 201218 330810 201454
rect 331046 201218 361530 201454
rect 361766 201218 392250 201454
rect 392486 201218 422970 201454
rect 423206 201218 453690 201454
rect 453926 201218 484410 201454
rect 484646 201218 515130 201454
rect 515366 201218 545850 201454
rect 546086 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect -2966 201134 586890 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 23610 201134
rect 23846 200898 54330 201134
rect 54566 200898 85050 201134
rect 85286 200898 115770 201134
rect 116006 200898 146490 201134
rect 146726 200898 177210 201134
rect 177446 200898 207930 201134
rect 208166 200898 238650 201134
rect 238886 200898 269370 201134
rect 269606 200898 300090 201134
rect 300326 200898 330810 201134
rect 331046 200898 361530 201134
rect 361766 200898 392250 201134
rect 392486 200898 422970 201134
rect 423206 200898 453690 201134
rect 453926 200898 484410 201134
rect 484646 200898 515130 201134
rect 515366 200898 545850 201134
rect 546086 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 592650 194294
rect -8726 194026 592650 194058
rect -6806 190894 590730 190926
rect -6806 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 590730 190894
rect -6806 190574 590730 190658
rect -6806 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 590730 190574
rect -6806 190306 590730 190338
rect -4886 187174 588810 187206
rect -4886 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 588810 187174
rect -4886 186854 588810 186938
rect -4886 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 588810 186854
rect -4886 186586 588810 186618
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 8250 183454
rect 8486 183218 38970 183454
rect 39206 183218 69690 183454
rect 69926 183218 100410 183454
rect 100646 183218 131130 183454
rect 131366 183218 161850 183454
rect 162086 183218 192570 183454
rect 192806 183218 223290 183454
rect 223526 183218 254010 183454
rect 254246 183218 284730 183454
rect 284966 183218 315450 183454
rect 315686 183218 346170 183454
rect 346406 183218 376890 183454
rect 377126 183218 407610 183454
rect 407846 183218 438330 183454
rect 438566 183218 469050 183454
rect 469286 183218 499770 183454
rect 500006 183218 530490 183454
rect 530726 183218 561210 183454
rect 561446 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 8250 183134
rect 8486 182898 38970 183134
rect 39206 182898 69690 183134
rect 69926 182898 100410 183134
rect 100646 182898 131130 183134
rect 131366 182898 161850 183134
rect 162086 182898 192570 183134
rect 192806 182898 223290 183134
rect 223526 182898 254010 183134
rect 254246 182898 284730 183134
rect 284966 182898 315450 183134
rect 315686 182898 346170 183134
rect 346406 182898 376890 183134
rect 377126 182898 407610 183134
rect 407846 182898 438330 183134
rect 438566 182898 469050 183134
rect 469286 182898 499770 183134
rect 500006 182898 530490 183134
rect 530726 182898 561210 183134
rect 561446 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect -8726 176614 592650 176646
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect -8726 176294 592650 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect -8726 176026 592650 176058
rect -6806 172894 590730 172926
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect -6806 172574 590730 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect -6806 172306 590730 172338
rect -4886 169174 588810 169206
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect -4886 168854 588810 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect -4886 168586 588810 168618
rect -2966 165454 586890 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 23610 165454
rect 23846 165218 54330 165454
rect 54566 165218 85050 165454
rect 85286 165218 115770 165454
rect 116006 165218 146490 165454
rect 146726 165218 177210 165454
rect 177446 165218 207930 165454
rect 208166 165218 238650 165454
rect 238886 165218 269370 165454
rect 269606 165218 300090 165454
rect 300326 165218 330810 165454
rect 331046 165218 361530 165454
rect 361766 165218 392250 165454
rect 392486 165218 422970 165454
rect 423206 165218 453690 165454
rect 453926 165218 484410 165454
rect 484646 165218 515130 165454
rect 515366 165218 545850 165454
rect 546086 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect -2966 165134 586890 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 23610 165134
rect 23846 164898 54330 165134
rect 54566 164898 85050 165134
rect 85286 164898 115770 165134
rect 116006 164898 146490 165134
rect 146726 164898 177210 165134
rect 177446 164898 207930 165134
rect 208166 164898 238650 165134
rect 238886 164898 269370 165134
rect 269606 164898 300090 165134
rect 300326 164898 330810 165134
rect 331046 164898 361530 165134
rect 361766 164898 392250 165134
rect 392486 164898 422970 165134
rect 423206 164898 453690 165134
rect 453926 164898 484410 165134
rect 484646 164898 515130 165134
rect 515366 164898 545850 165134
rect 546086 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect -2966 164866 586890 164898
rect -8726 158614 592650 158646
rect -8726 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 592650 158294
rect -8726 158026 592650 158058
rect -6806 154894 590730 154926
rect -6806 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 590730 154894
rect -6806 154574 590730 154658
rect -6806 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 590730 154574
rect -6806 154306 590730 154338
rect -4886 151174 588810 151206
rect -4886 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 588810 151174
rect -4886 150854 588810 150938
rect -4886 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 588810 150854
rect -4886 150586 588810 150618
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 8250 147454
rect 8486 147218 38970 147454
rect 39206 147218 69690 147454
rect 69926 147218 100410 147454
rect 100646 147218 131130 147454
rect 131366 147218 161850 147454
rect 162086 147218 192570 147454
rect 192806 147218 223290 147454
rect 223526 147218 254010 147454
rect 254246 147218 284730 147454
rect 284966 147218 315450 147454
rect 315686 147218 346170 147454
rect 346406 147218 376890 147454
rect 377126 147218 407610 147454
rect 407846 147218 438330 147454
rect 438566 147218 469050 147454
rect 469286 147218 499770 147454
rect 500006 147218 530490 147454
rect 530726 147218 561210 147454
rect 561446 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 8250 147134
rect 8486 146898 38970 147134
rect 39206 146898 69690 147134
rect 69926 146898 100410 147134
rect 100646 146898 131130 147134
rect 131366 146898 161850 147134
rect 162086 146898 192570 147134
rect 192806 146898 223290 147134
rect 223526 146898 254010 147134
rect 254246 146898 284730 147134
rect 284966 146898 315450 147134
rect 315686 146898 346170 147134
rect 346406 146898 376890 147134
rect 377126 146898 407610 147134
rect 407846 146898 438330 147134
rect 438566 146898 469050 147134
rect 469286 146898 499770 147134
rect 500006 146898 530490 147134
rect 530726 146898 561210 147134
rect 561446 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -8726 140614 592650 140646
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect -8726 140294 592650 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect -8726 140026 592650 140058
rect -6806 136894 590730 136926
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect -6806 136574 590730 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect -6806 136306 590730 136338
rect -4886 133174 588810 133206
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect -4886 132854 588810 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect -4886 132586 588810 132618
rect -2966 129454 586890 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 23610 129454
rect 23846 129218 54330 129454
rect 54566 129218 85050 129454
rect 85286 129218 115770 129454
rect 116006 129218 146490 129454
rect 146726 129218 177210 129454
rect 177446 129218 207930 129454
rect 208166 129218 238650 129454
rect 238886 129218 269370 129454
rect 269606 129218 300090 129454
rect 300326 129218 330810 129454
rect 331046 129218 361530 129454
rect 361766 129218 392250 129454
rect 392486 129218 422970 129454
rect 423206 129218 453690 129454
rect 453926 129218 484410 129454
rect 484646 129218 515130 129454
rect 515366 129218 545850 129454
rect 546086 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect -2966 129134 586890 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 23610 129134
rect 23846 128898 54330 129134
rect 54566 128898 85050 129134
rect 85286 128898 115770 129134
rect 116006 128898 146490 129134
rect 146726 128898 177210 129134
rect 177446 128898 207930 129134
rect 208166 128898 238650 129134
rect 238886 128898 269370 129134
rect 269606 128898 300090 129134
rect 300326 128898 330810 129134
rect 331046 128898 361530 129134
rect 361766 128898 392250 129134
rect 392486 128898 422970 129134
rect 423206 128898 453690 129134
rect 453926 128898 484410 129134
rect 484646 128898 515130 129134
rect 515366 128898 545850 129134
rect 546086 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect -2966 128866 586890 128898
rect -8726 122614 592650 122646
rect -8726 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 592650 122294
rect -8726 122026 592650 122058
rect -6806 118894 590730 118926
rect -6806 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 590730 118894
rect -6806 118574 590730 118658
rect -6806 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 590730 118574
rect -6806 118306 590730 118338
rect -4886 115174 588810 115206
rect -4886 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 588810 115174
rect -4886 114854 588810 114938
rect -4886 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 588810 114854
rect -4886 114586 588810 114618
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 8250 111454
rect 8486 111218 38970 111454
rect 39206 111218 69690 111454
rect 69926 111218 100410 111454
rect 100646 111218 131130 111454
rect 131366 111218 161850 111454
rect 162086 111218 192570 111454
rect 192806 111218 223290 111454
rect 223526 111218 254010 111454
rect 254246 111218 284730 111454
rect 284966 111218 315450 111454
rect 315686 111218 346170 111454
rect 346406 111218 376890 111454
rect 377126 111218 407610 111454
rect 407846 111218 438330 111454
rect 438566 111218 469050 111454
rect 469286 111218 499770 111454
rect 500006 111218 530490 111454
rect 530726 111218 561210 111454
rect 561446 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 8250 111134
rect 8486 110898 38970 111134
rect 39206 110898 69690 111134
rect 69926 110898 100410 111134
rect 100646 110898 131130 111134
rect 131366 110898 161850 111134
rect 162086 110898 192570 111134
rect 192806 110898 223290 111134
rect 223526 110898 254010 111134
rect 254246 110898 284730 111134
rect 284966 110898 315450 111134
rect 315686 110898 346170 111134
rect 346406 110898 376890 111134
rect 377126 110898 407610 111134
rect 407846 110898 438330 111134
rect 438566 110898 469050 111134
rect 469286 110898 499770 111134
rect 500006 110898 530490 111134
rect 530726 110898 561210 111134
rect 561446 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -8726 104614 592650 104646
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect -8726 104294 592650 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect -8726 104026 592650 104058
rect -6806 100894 590730 100926
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect -6806 100574 590730 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect -6806 100306 590730 100338
rect -4886 97174 588810 97206
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect -4886 96854 588810 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect -4886 96586 588810 96618
rect -2966 93454 586890 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 23610 93454
rect 23846 93218 54330 93454
rect 54566 93218 85050 93454
rect 85286 93218 115770 93454
rect 116006 93218 146490 93454
rect 146726 93218 177210 93454
rect 177446 93218 207930 93454
rect 208166 93218 238650 93454
rect 238886 93218 269370 93454
rect 269606 93218 300090 93454
rect 300326 93218 330810 93454
rect 331046 93218 361530 93454
rect 361766 93218 392250 93454
rect 392486 93218 422970 93454
rect 423206 93218 453690 93454
rect 453926 93218 484410 93454
rect 484646 93218 515130 93454
rect 515366 93218 545850 93454
rect 546086 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect -2966 93134 586890 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 23610 93134
rect 23846 92898 54330 93134
rect 54566 92898 85050 93134
rect 85286 92898 115770 93134
rect 116006 92898 146490 93134
rect 146726 92898 177210 93134
rect 177446 92898 207930 93134
rect 208166 92898 238650 93134
rect 238886 92898 269370 93134
rect 269606 92898 300090 93134
rect 300326 92898 330810 93134
rect 331046 92898 361530 93134
rect 361766 92898 392250 93134
rect 392486 92898 422970 93134
rect 423206 92898 453690 93134
rect 453926 92898 484410 93134
rect 484646 92898 515130 93134
rect 515366 92898 545850 93134
rect 546086 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect -2966 92866 586890 92898
rect -8726 86614 592650 86646
rect -8726 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 592650 86294
rect -8726 86026 592650 86058
rect -6806 82894 590730 82926
rect -6806 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 590730 82894
rect -6806 82574 590730 82658
rect -6806 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 590730 82574
rect -6806 82306 590730 82338
rect -4886 79174 588810 79206
rect -4886 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 588810 79174
rect -4886 78854 588810 78938
rect -4886 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 588810 78854
rect -4886 78586 588810 78618
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 8250 75454
rect 8486 75218 38970 75454
rect 39206 75218 69690 75454
rect 69926 75218 100410 75454
rect 100646 75218 131130 75454
rect 131366 75218 161850 75454
rect 162086 75218 192570 75454
rect 192806 75218 223290 75454
rect 223526 75218 254010 75454
rect 254246 75218 284730 75454
rect 284966 75218 315450 75454
rect 315686 75218 346170 75454
rect 346406 75218 376890 75454
rect 377126 75218 407610 75454
rect 407846 75218 438330 75454
rect 438566 75218 469050 75454
rect 469286 75218 499770 75454
rect 500006 75218 530490 75454
rect 530726 75218 561210 75454
rect 561446 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 8250 75134
rect 8486 74898 38970 75134
rect 39206 74898 69690 75134
rect 69926 74898 100410 75134
rect 100646 74898 131130 75134
rect 131366 74898 161850 75134
rect 162086 74898 192570 75134
rect 192806 74898 223290 75134
rect 223526 74898 254010 75134
rect 254246 74898 284730 75134
rect 284966 74898 315450 75134
rect 315686 74898 346170 75134
rect 346406 74898 376890 75134
rect 377126 74898 407610 75134
rect 407846 74898 438330 75134
rect 438566 74898 469050 75134
rect 469286 74898 499770 75134
rect 500006 74898 530490 75134
rect 530726 74898 561210 75134
rect 561446 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -8726 68614 592650 68646
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect -8726 68294 592650 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect -8726 68026 592650 68058
rect -6806 64894 590730 64926
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect -6806 64574 590730 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect -6806 64306 590730 64338
rect -4886 61174 588810 61206
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect -4886 60854 588810 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect -4886 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 23610 57454
rect 23846 57218 54330 57454
rect 54566 57218 85050 57454
rect 85286 57218 115770 57454
rect 116006 57218 146490 57454
rect 146726 57218 177210 57454
rect 177446 57218 207930 57454
rect 208166 57218 238650 57454
rect 238886 57218 269370 57454
rect 269606 57218 300090 57454
rect 300326 57218 330810 57454
rect 331046 57218 361530 57454
rect 361766 57218 392250 57454
rect 392486 57218 422970 57454
rect 423206 57218 453690 57454
rect 453926 57218 484410 57454
rect 484646 57218 515130 57454
rect 515366 57218 545850 57454
rect 546086 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 23610 57134
rect 23846 56898 54330 57134
rect 54566 56898 85050 57134
rect 85286 56898 115770 57134
rect 116006 56898 146490 57134
rect 146726 56898 177210 57134
rect 177446 56898 207930 57134
rect 208166 56898 238650 57134
rect 238886 56898 269370 57134
rect 269606 56898 300090 57134
rect 300326 56898 330810 57134
rect 331046 56898 361530 57134
rect 361766 56898 392250 57134
rect 392486 56898 422970 57134
rect 423206 56898 453690 57134
rect 453926 56898 484410 57134
rect 484646 56898 515130 57134
rect 515366 56898 545850 57134
rect 546086 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 592650 50294
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 590730 46894
rect -6806 46574 590730 46658
rect -6806 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 590730 46574
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 588810 43174
rect -4886 42854 588810 42938
rect -4886 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 588810 42854
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 8250 39454
rect 8486 39218 38970 39454
rect 39206 39218 69690 39454
rect 69926 39218 100410 39454
rect 100646 39218 131130 39454
rect 131366 39218 161850 39454
rect 162086 39218 192570 39454
rect 192806 39218 223290 39454
rect 223526 39218 254010 39454
rect 254246 39218 284730 39454
rect 284966 39218 315450 39454
rect 315686 39218 346170 39454
rect 346406 39218 376890 39454
rect 377126 39218 407610 39454
rect 407846 39218 438330 39454
rect 438566 39218 469050 39454
rect 469286 39218 499770 39454
rect 500006 39218 530490 39454
rect 530726 39218 561210 39454
rect 561446 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 8250 39134
rect 8486 38898 38970 39134
rect 39206 38898 69690 39134
rect 69926 38898 100410 39134
rect 100646 38898 131130 39134
rect 131366 38898 161850 39134
rect 162086 38898 192570 39134
rect 192806 38898 223290 39134
rect 223526 38898 254010 39134
rect 254246 38898 284730 39134
rect 284966 38898 315450 39134
rect 315686 38898 346170 39134
rect 346406 38898 376890 39134
rect 377126 38898 407610 39134
rect 407846 38898 438330 39134
rect 438566 38898 469050 39134
rect 469286 38898 499770 39134
rect 500006 38898 530490 39134
rect 530726 38898 561210 39134
rect 561446 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect -8726 32294 592650 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect -6806 28574 590730 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect -4886 24854 588810 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 23610 21454
rect 23846 21218 54330 21454
rect 54566 21218 85050 21454
rect 85286 21218 115770 21454
rect 116006 21218 146490 21454
rect 146726 21218 177210 21454
rect 177446 21218 207930 21454
rect 208166 21218 238650 21454
rect 238886 21218 269370 21454
rect 269606 21218 300090 21454
rect 300326 21218 330810 21454
rect 331046 21218 361530 21454
rect 361766 21218 392250 21454
rect 392486 21218 422970 21454
rect 423206 21218 453690 21454
rect 453926 21218 484410 21454
rect 484646 21218 515130 21454
rect 515366 21218 545850 21454
rect 546086 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 23610 21134
rect 23846 20898 54330 21134
rect 54566 20898 85050 21134
rect 85286 20898 115770 21134
rect 116006 20898 146490 21134
rect 146726 20898 177210 21134
rect 177446 20898 207930 21134
rect 208166 20898 238650 21134
rect 238886 20898 269370 21134
rect 269606 20898 300090 21134
rect 300326 20898 330810 21134
rect 331046 20898 361530 21134
rect 361766 20898 392250 21134
rect 392486 20898 422970 21134
rect 423206 20898 453690 21134
rect 453926 20898 484410 21134
rect 484646 20898 515130 21134
rect 515366 20898 545850 21134
rect 546086 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 592650 14294
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 590730 10894
rect -6806 10574 590730 10658
rect -6806 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 590730 10574
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 588810 7174
rect -4886 6854 588810 6938
rect -4886 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 588810 6854
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 8250 3454
rect 8486 3218 38970 3454
rect 39206 3218 69690 3454
rect 69926 3218 100410 3454
rect 100646 3218 131130 3454
rect 131366 3218 161850 3454
rect 162086 3218 192570 3454
rect 192806 3218 223290 3454
rect 223526 3218 254010 3454
rect 254246 3218 284730 3454
rect 284966 3218 315450 3454
rect 315686 3218 346170 3454
rect 346406 3218 376890 3454
rect 377126 3218 407610 3454
rect 407846 3218 438330 3454
rect 438566 3218 469050 3454
rect 469286 3218 499770 3454
rect 500006 3218 530490 3454
rect 530726 3218 561210 3454
rect 561446 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 8250 3134
rect 8486 2898 38970 3134
rect 39206 2898 69690 3134
rect 69926 2898 100410 3134
rect 100646 2898 131130 3134
rect 131366 2898 161850 3134
rect 162086 2898 192570 3134
rect 192806 2898 223290 3134
rect 223526 2898 254010 3134
rect 254246 2898 284730 3134
rect 284966 2898 315450 3134
rect 315686 2898 346170 3134
rect 346406 2898 376890 3134
rect 377126 2898 407610 3134
rect 407846 2898 438330 3134
rect 438566 2898 469050 3134
rect 469286 2898 499770 3134
rect 500006 2898 530490 3134
rect 530726 2898 561210 3134
rect 561446 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use user_proj  mprj
timestamp 1639392407
transform 1 0 4000 0 1 0
box 566 0 559438 700000
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 702000 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 702000 38414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 702000 74414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 702000 110414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 702000 146414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 702000 182414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 702000 218414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 702000 254414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 702000 290414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 702000 326414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 702000 362414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 702000 398414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 702000 434414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 702000 470414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 702000 506414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 702000 542414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 -3814 6134 -2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 41514 -3814 42134 -2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 77514 -3814 78134 -2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 113514 -3814 114134 -2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 149514 -3814 150134 -2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 185514 -3814 186134 -2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 221514 -3814 222134 -2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 257514 -3814 258134 -2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 293514 -3814 294134 -2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 329514 -3814 330134 -2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 365514 -3814 366134 -2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 401514 -3814 402134 -2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 437514 -3814 438134 -2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 473514 -3814 474134 -2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 509514 -3814 510134 -2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 545514 -3814 546134 -2000 8 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 702000 6134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 702000 42134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 702000 78134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 702000 114134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 702000 150134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 702000 186134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 702000 222134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 702000 258134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 702000 294134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 702000 330134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 702000 366134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 702000 402134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 702000 438134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 702000 474134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 702000 510134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 702000 546134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 581514 -3814 582134 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 -5734 9854 -2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 45234 -5734 45854 -2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 81234 -5734 81854 -2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 117234 -5734 117854 -2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 153234 -5734 153854 -2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 189234 -5734 189854 -2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 225234 -5734 225854 -2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 261234 -5734 261854 -2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 297234 -5734 297854 -2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 333234 -5734 333854 -2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 369234 -5734 369854 -2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 405234 -5734 405854 -2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 441234 -5734 441854 -2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 477234 -5734 477854 -2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 513234 -5734 513854 -2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 549234 -5734 549854 -2000 8 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 702000 9854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 702000 45854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 702000 81854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 702000 117854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 702000 153854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 702000 189854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 702000 225854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 702000 261854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 702000 297854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 702000 333854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 702000 369854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 702000 405854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 702000 441854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 702000 477854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 702000 513854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 702000 549854 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 -7654 13574 -2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 48954 -7654 49574 -2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 84954 -7654 85574 -2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 120954 -7654 121574 -2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 156954 -7654 157574 -2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 192954 -7654 193574 -2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 228954 -7654 229574 -2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 264954 -7654 265574 -2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 300954 -7654 301574 -2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 336954 -7654 337574 -2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 372954 -7654 373574 -2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 408954 -7654 409574 -2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 444954 -7654 445574 -2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 480954 -7654 481574 -2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 516954 -7654 517574 -2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 552954 -7654 553574 -2000 8 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 702000 13574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 702000 49574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 702000 85574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 702000 121574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 702000 157574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 702000 193574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 702000 229574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 702000 265574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 702000 301574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 702000 337574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 702000 373574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 702000 409574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 702000 445574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 702000 481574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 702000 517574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 702000 553574 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 -5734 27854 -2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 -5734 63854 -2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 -5734 99854 -2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 -5734 135854 -2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 -5734 171854 -2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 -5734 207854 -2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 -5734 243854 -2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 -5734 279854 -2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 -5734 315854 -2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 -5734 351854 -2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 -5734 387854 -2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 -5734 423854 -2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 -5734 459854 -2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 -5734 495854 -2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 -5734 531854 -2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 702000 27854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 702000 63854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 702000 99854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 702000 135854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 702000 171854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 702000 207854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 702000 243854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 702000 279854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 702000 315854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 702000 351854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 702000 387854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 702000 423854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 702000 459854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 702000 495854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 702000 531854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 -5734 567854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 -7654 31574 -2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 -7654 67574 -2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 -7654 103574 -2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 -7654 139574 -2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 -7654 175574 -2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 -7654 211574 -2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 -7654 247574 -2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 -7654 283574 -2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 -7654 319574 -2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 -7654 355574 -2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 -7654 391574 -2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 -7654 427574 -2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 -7654 463574 -2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 -7654 499574 -2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 -7654 535574 -2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 702000 31574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 702000 67574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 702000 103574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 702000 139574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 702000 175574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 702000 211574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 702000 247574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 702000 283574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 702000 319574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 702000 355574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 702000 391574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 702000 427574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 702000 463574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 702000 499574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 702000 535574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 -7654 571574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 702000 20414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 702000 56414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 702000 92414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 702000 128414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 702000 164414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 702000 200414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 702000 236414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 702000 272414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 702000 308414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 702000 344414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 702000 380414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 702000 416414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 702000 452414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 702000 488414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 702000 524414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 702000 560414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 -3814 24134 -2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 -3814 60134 -2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 -3814 96134 -2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 -3814 132134 -2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 -3814 168134 -2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 -3814 204134 -2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 -3814 240134 -2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 -3814 276134 -2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 -3814 312134 -2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 -3814 348134 -2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 -3814 384134 -2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 -3814 420134 -2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 -3814 456134 -2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 -3814 492134 -2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 -3814 528134 -2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 -3814 564134 -2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 702000 24134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 702000 60134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 702000 96134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 702000 132134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 702000 168134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 702000 204134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 702000 240134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 702000 276134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 702000 312134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 702000 348134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 702000 384134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 702000 420134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 702000 456134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 702000 492134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 702000 528134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 702000 564134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
