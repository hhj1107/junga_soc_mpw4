VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_proj
  CLASS BLOCK ;
  FOREIGN user_proj ;
  ORIGIN 0.000 0.000 ;
  SIZE 821.885 BY 832.605 ;
  PIN i_dout0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.470 828.605 553.750 832.605 ;
    END
  END i_dout0[0]
  PIN i_dout0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 817.885 378.800 821.885 379.400 ;
    END
  END i_dout0[10]
  PIN i_dout0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 817.885 415.520 821.885 416.120 ;
    END
  END i_dout0[11]
  PIN i_dout0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.490 0.000 685.770 4.000 ;
    END
  END i_dout0[12]
  PIN i_dout0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 817.885 451.560 821.885 452.160 ;
    END
  END i_dout0[13]
  PIN i_dout0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 710.330 828.605 710.610 832.605 ;
    END
  END i_dout0[14]
  PIN i_dout0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 705.270 0.000 705.550 4.000 ;
    END
  END i_dout0[15]
  PIN i_dout0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 817.885 499.840 821.885 500.440 ;
    END
  END i_dout0[16]
  PIN i_dout0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 729.190 828.605 729.470 832.605 ;
    END
  END i_dout0[17]
  PIN i_dout0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 817.885 548.120 821.885 548.720 ;
    END
  END i_dout0[18]
  PIN i_dout0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 738.850 828.605 739.130 832.605 ;
    END
  END i_dout0[19]
  PIN i_dout0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 817.885 65.320 821.885 65.920 ;
    END
  END i_dout0[1]
  PIN i_dout0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 748.050 828.605 748.330 832.605 ;
    END
  END i_dout0[20]
  PIN i_dout0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 749.890 0.000 750.170 4.000 ;
    END
  END i_dout0[21]
  PIN i_dout0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 753.110 828.605 753.390 832.605 ;
    END
  END i_dout0[22]
  PIN i_dout0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 817.885 632.440 821.885 633.040 ;
    END
  END i_dout0[23]
  PIN i_dout0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 767.370 828.605 767.650 832.605 ;
    END
  END i_dout0[24]
  PIN i_dout0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 781.630 828.605 781.910 832.605 ;
    END
  END i_dout0[25]
  PIN i_dout0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 817.885 680.720 821.885 681.320 ;
    END
  END i_dout0[26]
  PIN i_dout0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 817.885 741.240 821.885 741.840 ;
    END
  END i_dout0[27]
  PIN i_dout0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 794.510 0.000 794.790 4.000 ;
    END
  END i_dout0[28]
  PIN i_dout0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 817.885 789.520 821.885 790.120 ;
    END
  END i_dout0[29]
  PIN i_dout0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 817.885 101.360 821.885 101.960 ;
    END
  END i_dout0[2]
  PIN i_dout0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 809.230 0.000 809.510 4.000 ;
    END
  END i_dout0[30]
  PIN i_dout0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 819.350 828.605 819.630 832.605 ;
    END
  END i_dout0[31]
  PIN i_dout0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.450 828.605 605.730 832.605 ;
    END
  END i_dout0[3]
  PIN i_dout0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.080 4.000 138.680 ;
    END
  END i_dout0[4]
  PIN i_dout0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 629.370 828.605 629.650 832.605 ;
    END
  END i_dout0[5]
  PIN i_dout0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 626.150 0.000 626.430 4.000 ;
    END
  END i_dout0[6]
  PIN i_dout0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 817.885 282.920 821.885 283.520 ;
    END
  END i_dout0[7]
  PIN i_dout0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 817.885 318.960 821.885 319.560 ;
    END
  END i_dout0[8]
  PIN i_dout0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 817.885 330.520 821.885 331.120 ;
    END
  END i_dout0[9]
  PIN i_dout0_1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 556.690 0.000 556.970 4.000 ;
    END
  END i_dout0_1[0]
  PIN i_dout0_1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 817.885 367.240 821.885 367.840 ;
    END
  END i_dout0_1[10]
  PIN i_dout0_1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 817.885 403.280 821.885 403.880 ;
    END
  END i_dout0_1[11]
  PIN i_dout0_1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 817.885 439.320 821.885 439.920 ;
    END
  END i_dout0_1[12]
  PIN i_dout0_1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 690.550 0.000 690.830 4.000 ;
    END
  END i_dout0_1[13]
  PIN i_dout0_1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 817.885 463.800 821.885 464.400 ;
    END
  END i_dout0_1[14]
  PIN i_dout0_1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 700.210 0.000 700.490 4.000 ;
    END
  END i_dout0_1[15]
  PIN i_dout0_1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 459.040 4.000 459.640 ;
    END
  END i_dout0_1[16]
  PIN i_dout0_1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 503.240 4.000 503.840 ;
    END
  END i_dout0_1[17]
  PIN i_dout0_1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 733.790 828.605 734.070 832.605 ;
    END
  END i_dout0_1[18]
  PIN i_dout0_1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 590.280 4.000 590.880 ;
    END
  END i_dout0_1[19]
  PIN i_dout0_1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 817.885 53.080 821.885 53.680 ;
    END
  END i_dout0_1[1]
  PIN i_dout0_1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 817.885 571.920 821.885 572.520 ;
    END
  END i_dout0_1[20]
  PIN i_dout0_1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 744.830 0.000 745.110 4.000 ;
    END
  END i_dout0_1[21]
  PIN i_dout0_1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 817.885 596.400 821.885 597.000 ;
    END
  END i_dout0_1[22]
  PIN i_dout0_1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 757.710 828.605 757.990 832.605 ;
    END
  END i_dout0_1[23]
  PIN i_dout0_1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 722.200 4.000 722.800 ;
    END
  END i_dout0_1[24]
  PIN i_dout0_1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 771.970 828.605 772.250 832.605 ;
    END
  END i_dout0_1[25]
  PIN i_dout0_1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 784.390 0.000 784.670 4.000 ;
    END
  END i_dout0_1[26]
  PIN i_dout0_1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 817.885 729.000 821.885 729.600 ;
    END
  END i_dout0_1[27]
  PIN i_dout0_1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 817.885 765.040 821.885 765.640 ;
    END
  END i_dout0_1[28]
  PIN i_dout0_1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 780.680 4.000 781.280 ;
    END
  END i_dout0_1[29]
  PIN i_dout0_1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 591.190 828.605 591.470 832.605 ;
    END
  END i_dout0_1[2]
  PIN i_dout0_1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 817.885 801.080 821.885 801.680 ;
    END
  END i_dout0_1[30]
  PIN i_dout0_1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 814.750 828.605 815.030 832.605 ;
    END
  END i_dout0_1[31]
  PIN i_dout0_1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 79.600 4.000 80.200 ;
    END
  END i_dout0_1[3]
  PIN i_dout0_1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.430 0.000 611.710 4.000 ;
    END
  END i_dout0_1[4]
  PIN i_dout0_1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 196.560 4.000 197.160 ;
    END
  END i_dout0_1[5]
  PIN i_dout0_1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 225.800 4.000 226.400 ;
    END
  END i_dout0_1[6]
  PIN i_dout0_1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 635.810 0.000 636.090 4.000 ;
    END
  END i_dout0_1[7]
  PIN i_dout0_1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 284.280 4.000 284.880 ;
    END
  END i_dout0_1[8]
  PIN i_dout0_1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 327.800 4.000 328.400 ;
    END
  END i_dout0_1[9]
  PIN i_dout1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 558.070 828.605 558.350 832.605 ;
    END
  END i_dout1[0]
  PIN i_dout1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 817.885 391.040 821.885 391.640 ;
    END
  END i_dout1[10]
  PIN i_dout1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 691.010 828.605 691.290 832.605 ;
    END
  END i_dout1[11]
  PIN i_dout1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 386.280 4.000 386.880 ;
    END
  END i_dout1[12]
  PIN i_dout1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 429.800 4.000 430.400 ;
    END
  END i_dout1[13]
  PIN i_dout1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 817.885 475.360 821.885 475.960 ;
    END
  END i_dout1[14]
  PIN i_dout1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 710.330 0.000 710.610 4.000 ;
    END
  END i_dout1[15]
  PIN i_dout1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 474.000 4.000 474.600 ;
    END
  END i_dout1[16]
  PIN i_dout1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 817.885 523.640 821.885 524.240 ;
    END
  END i_dout1[17]
  PIN i_dout1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 546.760 4.000 547.360 ;
    END
  END i_dout1[18]
  PIN i_dout1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 725.050 0.000 725.330 4.000 ;
    END
  END i_dout1[19]
  PIN i_dout1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 817.885 77.560 821.885 78.160 ;
    END
  END i_dout1[1]
  PIN i_dout1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 619.520 4.000 620.120 ;
    END
  END i_dout1[20]
  PIN i_dout1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 817.885 584.160 821.885 584.760 ;
    END
  END i_dout1[21]
  PIN i_dout1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 817.885 607.960 821.885 608.560 ;
    END
  END i_dout1[22]
  PIN i_dout1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.010 0.000 760.290 4.000 ;
    END
  END i_dout1[23]
  PIN i_dout1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 817.885 644.680 821.885 645.280 ;
    END
  END i_dout1[24]
  PIN i_dout1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 774.730 0.000 775.010 4.000 ;
    END
  END i_dout1[25]
  PIN i_dout1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 817.885 692.960 821.885 693.560 ;
    END
  END i_dout1[26]
  PIN i_dout1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 817.885 752.800 821.885 753.400 ;
    END
  END i_dout1[27]
  PIN i_dout1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 795.890 828.605 796.170 832.605 ;
    END
  END i_dout1[28]
  PIN i_dout1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 805.090 828.605 805.370 832.605 ;
    END
  END i_dout1[29]
  PIN i_dout1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 817.885 113.600 821.885 114.200 ;
    END
  END i_dout1[2]
  PIN i_dout1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 810.150 828.605 810.430 832.605 ;
    END
  END i_dout1[30]
  PIN i_dout1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 824.200 4.000 824.800 ;
    END
  END i_dout1[31]
  PIN i_dout1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END i_dout1[3]
  PIN i_dout1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 152.360 4.000 152.960 ;
    END
  END i_dout1[4]
  PIN i_dout1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 817.885 210.160 821.885 210.760 ;
    END
  END i_dout1[5]
  PIN i_dout1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 631.210 0.000 631.490 4.000 ;
    END
  END i_dout1[6]
  PIN i_dout1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 817.885 294.480 821.885 295.080 ;
    END
  END i_dout1[7]
  PIN i_dout1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 298.560 4.000 299.160 ;
    END
  END i_dout1[8]
  PIN i_dout1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 817.885 342.760 821.885 343.360 ;
    END
  END i_dout1[9]
  PIN i_dout1_1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 817.885 5.480 821.885 6.080 ;
    END
  END i_dout1_1[0]
  PIN i_dout1_1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 686.410 828.605 686.690 832.605 ;
    END
  END i_dout1_1[10]
  PIN i_dout1_1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 357.040 4.000 357.640 ;
    END
  END i_dout1_1[11]
  PIN i_dout1_1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 680.430 0.000 680.710 4.000 ;
    END
  END i_dout1_1[12]
  PIN i_dout1_1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 415.520 4.000 416.120 ;
    END
  END i_dout1_1[13]
  PIN i_dout1_1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 705.270 828.605 705.550 832.605 ;
    END
  END i_dout1_1[14]
  PIN i_dout1_1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 719.530 828.605 719.810 832.605 ;
    END
  END i_dout1_1[15]
  PIN i_dout1_1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 724.590 828.605 724.870 832.605 ;
    END
  END i_dout1_1[16]
  PIN i_dout1_1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 817.885 512.080 821.885 512.680 ;
    END
  END i_dout1_1[17]
  PIN i_dout1_1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 532.480 4.000 533.080 ;
    END
  END i_dout1_1[18]
  PIN i_dout1_1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 817.885 560.360 821.885 560.960 ;
    END
  END i_dout1_1[19]
  PIN i_dout1_1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.930 828.605 577.210 832.605 ;
    END
  END i_dout1_1[1]
  PIN i_dout1_1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 605.240 4.000 605.840 ;
    END
  END i_dout1_1[20]
  PIN i_dout1_1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 634.480 4.000 635.080 ;
    END
  END i_dout1_1[21]
  PIN i_dout1_1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 754.950 0.000 755.230 4.000 ;
    END
  END i_dout1_1[22]
  PIN i_dout1_1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 762.310 828.605 762.590 832.605 ;
    END
  END i_dout1_1[23]
  PIN i_dout1_1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 764.610 0.000 764.890 4.000 ;
    END
  END i_dout1_1[24]
  PIN i_dout1_1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 776.570 828.605 776.850 832.605 ;
    END
  END i_dout1_1[25]
  PIN i_dout1_1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 789.450 0.000 789.730 4.000 ;
    END
  END i_dout1_1[26]
  PIN i_dout1_1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 786.230 828.605 786.510 832.605 ;
    END
  END i_dout1_1[27]
  PIN i_dout1_1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 751.440 4.000 752.040 ;
    END
  END i_dout1_1[28]
  PIN i_dout1_1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 817.885 777.280 821.885 777.880 ;
    END
  END i_dout1_1[29]
  PIN i_dout1_1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 591.650 0.000 591.930 4.000 ;
    END
  END i_dout1_1[2]
  PIN i_dout1_1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 804.170 0.000 804.450 4.000 ;
    END
  END i_dout1_1[30]
  PIN i_dout1_1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 817.885 825.560 821.885 826.160 ;
    END
  END i_dout1_1[31]
  PIN i_dout1_1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.880 4.000 94.480 ;
    END
  END i_dout1_1[3]
  PIN i_dout1_1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 817.885 174.120 821.885 174.720 ;
    END
  END i_dout1_1[4]
  PIN i_dout1_1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 621.090 0.000 621.370 4.000 ;
    END
  END i_dout1_1[5]
  PIN i_dout1_1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 653.290 828.605 653.570 832.605 ;
    END
  END i_dout1_1[6]
  PIN i_dout1_1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 657.890 828.605 658.170 832.605 ;
    END
  END i_dout1_1[7]
  PIN i_dout1_1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 672.150 828.605 672.430 832.605 ;
    END
  END i_dout1_1[8]
  PIN i_dout1_1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 665.710 0.000 665.990 4.000 ;
    END
  END i_dout1_1[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.390 828.605 2.670 832.605 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.530 828.605 144.810 832.605 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.790 828.605 159.070 832.605 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.050 828.605 173.330 832.605 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.310 828.605 187.590 832.605 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.570 828.605 201.850 832.605 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.830 828.605 216.110 832.605 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.090 828.605 230.370 832.605 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.350 828.605 244.630 832.605 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.610 828.605 258.890 832.605 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.870 828.605 273.150 832.605 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 828.605 16.470 832.605 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.130 828.605 287.410 832.605 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.390 828.605 301.670 832.605 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.650 828.605 315.930 832.605 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.910 828.605 330.190 832.605 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.170 828.605 344.450 832.605 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.430 828.605 358.710 832.605 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 372.690 828.605 372.970 832.605 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.950 828.605 387.230 832.605 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 401.210 828.605 401.490 832.605 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.470 828.605 415.750 832.605 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.450 828.605 30.730 832.605 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 429.730 828.605 430.010 832.605 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.990 828.605 444.270 832.605 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 458.250 828.605 458.530 832.605 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.510 828.605 472.790 832.605 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 486.770 828.605 487.050 832.605 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.030 828.605 501.310 832.605 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 515.290 828.605 515.570 832.605 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 529.550 828.605 529.830 832.605 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.710 828.605 44.990 832.605 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.970 828.605 59.250 832.605 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.230 828.605 73.510 832.605 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.490 828.605 87.770 832.605 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.750 828.605 102.030 832.605 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 828.605 116.290 832.605 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.270 828.605 130.550 832.605 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 828.605 7.270 832.605 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.590 828.605 149.870 832.605 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.850 828.605 164.130 832.605 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.110 828.605 178.390 832.605 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.370 828.605 192.650 832.605 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.630 828.605 206.910 832.605 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.890 828.605 221.170 832.605 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.150 828.605 235.430 832.605 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.410 828.605 249.690 832.605 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.670 828.605 263.950 832.605 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.930 828.605 278.210 832.605 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.250 828.605 21.530 832.605 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.190 828.605 292.470 832.605 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.450 828.605 306.730 832.605 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 320.710 828.605 320.990 832.605 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.970 828.605 335.250 832.605 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 349.230 828.605 349.510 832.605 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.490 828.605 363.770 832.605 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.750 828.605 378.030 832.605 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.010 828.605 392.290 832.605 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 406.270 828.605 406.550 832.605 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.070 828.605 420.350 832.605 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 828.605 35.790 832.605 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.330 828.605 434.610 832.605 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 448.590 828.605 448.870 832.605 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 462.850 828.605 463.130 832.605 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 477.110 828.605 477.390 832.605 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 491.370 828.605 491.650 832.605 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.630 828.605 505.910 832.605 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 519.890 828.605 520.170 832.605 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.150 828.605 534.430 832.605 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.770 828.605 50.050 832.605 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.030 828.605 64.310 832.605 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.290 828.605 78.570 832.605 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.550 828.605 92.830 832.605 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.810 828.605 107.090 832.605 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.070 828.605 121.350 832.605 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 828.605 135.610 832.605 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 828.605 11.870 832.605 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.190 828.605 154.470 832.605 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.450 828.605 168.730 832.605 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.710 828.605 182.990 832.605 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.970 828.605 197.250 832.605 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.230 828.605 211.510 832.605 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 828.605 225.770 832.605 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.750 828.605 240.030 832.605 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.010 828.605 254.290 832.605 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.270 828.605 268.550 832.605 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.530 828.605 282.810 832.605 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 828.605 26.130 832.605 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.790 828.605 297.070 832.605 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.050 828.605 311.330 832.605 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.310 828.605 325.590 832.605 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.570 828.605 339.850 832.605 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 353.830 828.605 354.110 832.605 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.090 828.605 368.370 832.605 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 382.350 828.605 382.630 832.605 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.610 828.605 396.890 832.605 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.870 828.605 411.150 832.605 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.130 828.605 425.410 832.605 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.110 828.605 40.390 832.605 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.390 828.605 439.670 832.605 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 453.650 828.605 453.930 832.605 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 467.910 828.605 468.190 832.605 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 482.170 828.605 482.450 832.605 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.430 828.605 496.710 832.605 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 510.690 828.605 510.970 832.605 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.950 828.605 525.230 832.605 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 539.210 828.605 539.490 832.605 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.370 828.605 54.650 832.605 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.630 828.605 68.910 832.605 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.890 828.605 83.170 832.605 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.150 828.605 97.430 832.605 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.410 828.605 111.690 832.605 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 828.605 125.950 832.605 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.930 828.605 140.210 832.605 ;
    END
  END io_out[9]
  PIN irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 527.250 0.000 527.530 4.000 ;
    END
  END irq[0]
  PIN irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.850 0.000 532.130 4.000 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 536.910 0.000 537.190 4.000 ;
    END
  END irq[2]
  PIN o_addr1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 562.670 828.605 562.950 832.605 ;
    END
  END o_addr1[0]
  PIN o_addr1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 817.885 89.800 821.885 90.400 ;
    END
  END o_addr1[1]
  PIN o_addr1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 50.360 4.000 50.960 ;
    END
  END o_addr1[2]
  PIN o_addr1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 615.110 828.605 615.390 832.605 ;
    END
  END o_addr1[3]
  PIN o_addr1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 167.320 4.000 167.920 ;
    END
  END o_addr1[4]
  PIN o_addr1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 639.030 828.605 639.310 832.605 ;
    END
  END o_addr1[5]
  PIN o_addr1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 240.080 4.000 240.680 ;
    END
  END o_addr1[6]
  PIN o_addr1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 662.490 828.605 662.770 832.605 ;
    END
  END o_addr1[7]
  PIN o_addr1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 655.590 0.000 655.870 4.000 ;
    END
  END o_addr1[8]
  PIN o_addr1_1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 817.885 17.040 821.885 17.640 ;
    END
  END o_addr1_1[0]
  PIN o_addr1_1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.990 828.605 582.270 832.605 ;
    END
  END o_addr1_1[1]
  PIN o_addr1_1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.400 4.000 36.000 ;
    END
  END o_addr1_1[2]
  PIN o_addr1_1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 610.510 828.605 610.790 832.605 ;
    END
  END o_addr1_1[3]
  PIN o_addr1_1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 624.770 828.605 625.050 832.605 ;
    END
  END o_addr1_1[4]
  PIN o_addr1_1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 633.970 828.605 634.250 832.605 ;
    END
  END o_addr1_1[5]
  PIN o_addr1_1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 817.885 234.640 821.885 235.240 ;
    END
  END o_addr1_1[6]
  PIN o_addr1_1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 640.870 0.000 641.150 4.000 ;
    END
  END o_addr1_1[7]
  PIN o_addr1_1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.990 0.000 651.270 4.000 ;
    END
  END o_addr1_1[8]
  PIN o_csb0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.970 0.000 542.250 4.000 ;
    END
  END o_csb0
  PIN o_csb0_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 543.810 828.605 544.090 832.605 ;
    END
  END o_csb0_1
  PIN o_csb1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 548.410 828.605 548.690 832.605 ;
    END
  END o_csb1
  PIN o_csb1_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.030 0.000 547.310 4.000 ;
    END
  END o_csb1_1
  PIN o_din0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 817.885 29.280 821.885 29.880 ;
    END
  END o_din0[0]
  PIN o_din0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 675.830 0.000 676.110 4.000 ;
    END
  END o_din0[10]
  PIN o_din0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 817.885 427.080 821.885 427.680 ;
    END
  END o_din0[11]
  PIN o_din0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 400.560 4.000 401.160 ;
    END
  END o_din0[12]
  PIN o_din0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.610 0.000 695.890 4.000 ;
    END
  END o_din0[13]
  PIN o_din0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 714.930 828.605 715.210 832.605 ;
    END
  END o_din0[14]
  PIN o_din0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 817.885 487.600 821.885 488.200 ;
    END
  END o_din0[15]
  PIN o_din0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 719.990 0.000 720.270 4.000 ;
    END
  END o_din0[16]
  PIN o_din0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 817.885 535.880 821.885 536.480 ;
    END
  END o_din0[17]
  PIN o_din0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 576.000 4.000 576.600 ;
    END
  END o_din0[18]
  PIN o_din0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 743.450 828.605 743.730 832.605 ;
    END
  END o_din0[19]
  PIN o_din0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.470 0.000 576.750 4.000 ;
    END
  END o_din0[1]
  PIN o_din0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 739.770 0.000 740.050 4.000 ;
    END
  END o_din0[20]
  PIN o_din0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 663.720 4.000 664.320 ;
    END
  END o_din0[21]
  PIN o_din0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 817.885 620.200 821.885 620.800 ;
    END
  END o_din0[22]
  PIN o_din0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 707.240 4.000 707.840 ;
    END
  END o_din0[23]
  PIN o_din0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 817.885 656.240 821.885 656.840 ;
    END
  END o_din0[24]
  PIN o_din0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 817.885 668.480 821.885 669.080 ;
    END
  END o_din0[25]
  PIN o_din0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 817.885 716.760 821.885 717.360 ;
    END
  END o_din0[26]
  PIN o_din0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 736.480 4.000 737.080 ;
    END
  END o_din0[27]
  PIN o_din0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 800.490 828.605 800.770 832.605 ;
    END
  END o_din0[28]
  PIN o_din0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 794.960 4.000 795.560 ;
    END
  END o_din0[29]
  PIN o_din0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END o_din0[2]
  PIN o_din0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 809.920 4.000 810.520 ;
    END
  END o_din0[30]
  PIN o_din0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 819.350 0.000 819.630 4.000 ;
    END
  END o_din0[31]
  PIN o_din0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 817.885 149.640 821.885 150.240 ;
    END
  END o_din0[3]
  PIN o_din0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 181.600 4.000 182.200 ;
    END
  END o_din0[4]
  PIN o_din0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 648.230 828.605 648.510 832.605 ;
    END
  END o_din0[5]
  PIN o_din0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 817.885 258.440 821.885 259.040 ;
    END
  END o_din0[6]
  PIN o_din0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 269.320 4.000 269.920 ;
    END
  END o_din0[7]
  PIN o_din0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 660.650 0.000 660.930 4.000 ;
    END
  END o_din0[8]
  PIN o_din0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 817.885 355.000 821.885 355.600 ;
    END
  END o_din0[9]
  PIN o_din0_1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 567.730 828.605 568.010 832.605 ;
    END
  END o_din0_1[0]
  PIN o_din0_1[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 670.770 0.000 671.050 4.000 ;
    END
  END o_din0_1[10]
  PIN o_din0_1[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 371.320 4.000 371.920 ;
    END
  END o_din0_1[11]
  PIN o_din0_1[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 696.070 828.605 696.350 832.605 ;
    END
  END o_din0_1[12]
  PIN o_din0_1[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 700.670 828.605 700.950 832.605 ;
    END
  END o_din0_1[13]
  PIN o_din0_1[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 444.760 4.000 445.360 ;
    END
  END o_din0_1[14]
  PIN o_din0_1[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 715.390 0.000 715.670 4.000 ;
    END
  END o_din0_1[15]
  PIN o_din0_1[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 488.280 4.000 488.880 ;
    END
  END o_din0_1[16]
  PIN o_din0_1[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 517.520 4.000 518.120 ;
    END
  END o_din0_1[17]
  PIN o_din0_1[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 561.720 4.000 562.320 ;
    END
  END o_din0_1[18]
  PIN o_din0_1[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 730.110 0.000 730.390 4.000 ;
    END
  END o_din0_1[19]
  PIN o_din0_1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 571.410 0.000 571.690 4.000 ;
    END
  END o_din0_1[1]
  PIN o_din0_1[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 735.170 0.000 735.450 4.000 ;
    END
  END o_din0_1[20]
  PIN o_din0_1[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 648.760 4.000 649.360 ;
    END
  END o_din0_1[21]
  PIN o_din0_1[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 678.000 4.000 678.600 ;
    END
  END o_din0_1[22]
  PIN o_din0_1[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 692.960 4.000 693.560 ;
    END
  END o_din0_1[23]
  PIN o_din0_1[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 769.670 0.000 769.950 4.000 ;
    END
  END o_din0_1[24]
  PIN o_din0_1[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 779.790 0.000 780.070 4.000 ;
    END
  END o_din0_1[25]
  PIN o_din0_1[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 817.885 704.520 821.885 705.120 ;
    END
  END o_din0_1[26]
  PIN o_din0_1[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 790.830 828.605 791.110 832.605 ;
    END
  END o_din0_1[27]
  PIN o_din0_1[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 765.720 4.000 766.320 ;
    END
  END o_din0_1[28]
  PIN o_din0_1[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 799.570 0.000 799.850 4.000 ;
    END
  END o_din0_1[29]
  PIN o_din0_1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 596.250 0.000 596.530 4.000 ;
    END
  END o_din0_1[2]
  PIN o_din0_1[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 817.885 813.320 821.885 813.920 ;
    END
  END o_din0_1[30]
  PIN o_din0_1[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 814.290 0.000 814.570 4.000 ;
    END
  END o_din0_1[31]
  PIN o_din0_1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.120 4.000 123.720 ;
    END
  END o_din0_1[3]
  PIN o_din0_1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 817.885 186.360 821.885 186.960 ;
    END
  END o_din0_1[4]
  PIN o_din0_1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 643.630 828.605 643.910 832.605 ;
    END
  END o_din0_1[5]
  PIN o_din0_1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 817.885 246.200 821.885 246.800 ;
    END
  END o_din0_1[6]
  PIN o_din0_1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 645.930 0.000 646.210 4.000 ;
    END
  END o_din0_1[7]
  PIN o_din0_1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.750 828.605 677.030 832.605 ;
    END
  END o_din0_1[8]
  PIN o_din0_1[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 342.080 4.000 342.680 ;
    END
  END o_din0_1[9]
  PIN o_waddr0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 572.330 828.605 572.610 832.605 ;
    END
  END o_waddr0[0]
  PIN o_waddr0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.590 828.605 586.870 832.605 ;
    END
  END o_waddr0[1]
  PIN o_waddr0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 817.885 125.840 821.885 126.440 ;
    END
  END o_waddr0[2]
  PIN o_waddr0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 601.310 0.000 601.590 4.000 ;
    END
  END o_waddr0[3]
  PIN o_waddr0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 616.030 0.000 616.310 4.000 ;
    END
  END o_waddr0[4]
  PIN o_waddr0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 817.885 222.400 821.885 223.000 ;
    END
  END o_waddr0[5]
  PIN o_waddr0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.040 4.000 255.640 ;
    END
  END o_waddr0[6]
  PIN o_waddr0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 817.885 306.720 821.885 307.320 ;
    END
  END o_waddr0[7]
  PIN o_waddr0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.840 4.000 313.440 ;
    END
  END o_waddr0[8]
  PIN o_waddr0_1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 817.885 41.520 821.885 42.120 ;
    END
  END o_waddr0_1[0]
  PIN o_waddr0_1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.120 4.000 21.720 ;
    END
  END o_waddr0_1[1]
  PIN o_waddr0_1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 596.250 828.605 596.530 832.605 ;
    END
  END o_waddr0_1[2]
  PIN o_waddr0_1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 817.885 161.880 821.885 162.480 ;
    END
  END o_waddr0_1[3]
  PIN o_waddr0_1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 817.885 197.920 821.885 198.520 ;
    END
  END o_waddr0_1[4]
  PIN o_waddr0_1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.840 4.000 211.440 ;
    END
  END o_waddr0_1[5]
  PIN o_waddr0_1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 817.885 270.680 821.885 271.280 ;
    END
  END o_waddr0_1[6]
  PIN o_waddr0_1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 667.550 828.605 667.830 832.605 ;
    END
  END o_waddr0_1[7]
  PIN o_waddr0_1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 681.810 828.605 682.090 832.605 ;
    END
  END o_waddr0_1[8]
  PIN o_web0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 551.630 0.000 551.910 4.000 ;
    END
  END o_web0
  PIN o_web0_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END o_web0_1
  PIN o_wmask0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 561.750 0.000 562.030 4.000 ;
    END
  END o_wmask0[0]
  PIN o_wmask0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.590 0.000 586.870 4.000 ;
    END
  END o_wmask0[1]
  PIN o_wmask0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 600.850 828.605 601.130 832.605 ;
    END
  END o_wmask0[2]
  PIN o_wmask0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 606.370 0.000 606.650 4.000 ;
    END
  END o_wmask0[3]
  PIN o_wmask0_1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 566.810 0.000 567.090 4.000 ;
    END
  END o_wmask0_1[0]
  PIN o_wmask0_1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.530 0.000 581.810 4.000 ;
    END
  END o_wmask0_1[1]
  PIN o_wmask0_1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 817.885 138.080 821.885 138.680 ;
    END
  END o_wmask0_1[2]
  PIN o_wmask0_1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 619.710 828.605 619.990 832.605 ;
    END
  END o_wmask0_1[3]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 821.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 821.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 821.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 821.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 821.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 821.680 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 821.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 821.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 821.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 821.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 821.680 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.390 0.000 2.670 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 0.000 7.270 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.050 0.000 12.330 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.830 0.000 32.110 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.190 0.000 200.470 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.910 0.000 215.190 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.090 0.000 230.370 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.810 0.000 245.090 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.530 0.000 259.810 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.710 0.000 274.990 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.430 0.000 289.710 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.150 0.000 304.430 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.870 0.000 319.150 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.050 0.000 334.330 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 348.770 0.000 349.050 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.490 0.000 363.770 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.670 0.000 378.950 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 393.390 0.000 393.670 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 408.110 0.000 408.390 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 423.290 0.000 423.570 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.010 0.000 438.290 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 452.730 0.000 453.010 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 467.450 0.000 467.730 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 482.630 0.000 482.910 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.390 0.000 71.670 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 497.350 0.000 497.630 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.070 0.000 512.350 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.170 0.000 91.450 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.950 0.000 111.230 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.130 0.000 126.410 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.850 0.000 141.130 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.570 0.000 155.850 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 0.000 171.030 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.470 0.000 185.750 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.110 0.000 17.390 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.890 0.000 37.170 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.250 0.000 205.530 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.970 0.000 220.250 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.690 0.000 234.970 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.870 0.000 250.150 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.590 0.000 264.870 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.310 0.000 279.590 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.490 0.000 294.770 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.210 0.000 309.490 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.930 0.000 324.210 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.110 0.000 339.390 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.670 0.000 56.950 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 353.830 0.000 354.110 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.550 0.000 368.830 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.270 0.000 383.550 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.450 0.000 398.730 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 413.170 0.000 413.450 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 427.890 0.000 428.170 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.070 0.000 443.350 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.790 0.000 458.070 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.510 0.000 472.790 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 487.230 0.000 487.510 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.450 0.000 76.730 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.410 0.000 502.690 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 517.130 0.000 517.410 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.230 0.000 96.510 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 0.000 116.290 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.730 0.000 131.010 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.910 0.000 146.190 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.630 0.000 160.910 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.350 0.000 175.630 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.530 0.000 190.810 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.310 0.000 210.590 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.030 0.000 225.310 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.750 0.000 240.030 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.930 0.000 255.210 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.650 0.000 269.930 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.370 0.000 284.650 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.090 0.000 299.370 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.270 0.000 314.550 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.990 0.000 329.270 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.710 0.000 343.990 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.730 0.000 62.010 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.890 0.000 359.170 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.610 0.000 373.890 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 388.330 0.000 388.610 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.050 0.000 403.330 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.230 0.000 418.510 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.950 0.000 433.230 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.670 0.000 447.950 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 462.850 0.000 463.130 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 477.570 0.000 477.850 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.290 0.000 492.570 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.510 0.000 81.790 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.470 0.000 507.750 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.190 0.000 522.470 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.290 0.000 101.570 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.070 0.000 121.350 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.790 0.000 136.070 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.510 0.000 150.790 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.690 0.000 165.970 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 0.000 180.690 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.130 0.000 195.410 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.550 0.000 46.830 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.330 0.000 66.610 4.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.570 0.000 86.850 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 0.000 106.630 4.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.170 0.000 22.450 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.770 0.000 27.050 4.000 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 816.815 821.525 ;
      LAYER met1 ;
        RECT 0.530 1.740 819.650 821.680 ;
      LAYER met2 ;
        RECT 0.560 828.325 2.110 829.330 ;
        RECT 2.950 828.325 6.710 829.330 ;
        RECT 7.550 828.325 11.310 829.330 ;
        RECT 12.150 828.325 15.910 829.330 ;
        RECT 16.750 828.325 20.970 829.330 ;
        RECT 21.810 828.325 25.570 829.330 ;
        RECT 26.410 828.325 30.170 829.330 ;
        RECT 31.010 828.325 35.230 829.330 ;
        RECT 36.070 828.325 39.830 829.330 ;
        RECT 40.670 828.325 44.430 829.330 ;
        RECT 45.270 828.325 49.490 829.330 ;
        RECT 50.330 828.325 54.090 829.330 ;
        RECT 54.930 828.325 58.690 829.330 ;
        RECT 59.530 828.325 63.750 829.330 ;
        RECT 64.590 828.325 68.350 829.330 ;
        RECT 69.190 828.325 72.950 829.330 ;
        RECT 73.790 828.325 78.010 829.330 ;
        RECT 78.850 828.325 82.610 829.330 ;
        RECT 83.450 828.325 87.210 829.330 ;
        RECT 88.050 828.325 92.270 829.330 ;
        RECT 93.110 828.325 96.870 829.330 ;
        RECT 97.710 828.325 101.470 829.330 ;
        RECT 102.310 828.325 106.530 829.330 ;
        RECT 107.370 828.325 111.130 829.330 ;
        RECT 111.970 828.325 115.730 829.330 ;
        RECT 116.570 828.325 120.790 829.330 ;
        RECT 121.630 828.325 125.390 829.330 ;
        RECT 126.230 828.325 129.990 829.330 ;
        RECT 130.830 828.325 135.050 829.330 ;
        RECT 135.890 828.325 139.650 829.330 ;
        RECT 140.490 828.325 144.250 829.330 ;
        RECT 145.090 828.325 149.310 829.330 ;
        RECT 150.150 828.325 153.910 829.330 ;
        RECT 154.750 828.325 158.510 829.330 ;
        RECT 159.350 828.325 163.570 829.330 ;
        RECT 164.410 828.325 168.170 829.330 ;
        RECT 169.010 828.325 172.770 829.330 ;
        RECT 173.610 828.325 177.830 829.330 ;
        RECT 178.670 828.325 182.430 829.330 ;
        RECT 183.270 828.325 187.030 829.330 ;
        RECT 187.870 828.325 192.090 829.330 ;
        RECT 192.930 828.325 196.690 829.330 ;
        RECT 197.530 828.325 201.290 829.330 ;
        RECT 202.130 828.325 206.350 829.330 ;
        RECT 207.190 828.325 210.950 829.330 ;
        RECT 211.790 828.325 215.550 829.330 ;
        RECT 216.390 828.325 220.610 829.330 ;
        RECT 221.450 828.325 225.210 829.330 ;
        RECT 226.050 828.325 229.810 829.330 ;
        RECT 230.650 828.325 234.870 829.330 ;
        RECT 235.710 828.325 239.470 829.330 ;
        RECT 240.310 828.325 244.070 829.330 ;
        RECT 244.910 828.325 249.130 829.330 ;
        RECT 249.970 828.325 253.730 829.330 ;
        RECT 254.570 828.325 258.330 829.330 ;
        RECT 259.170 828.325 263.390 829.330 ;
        RECT 264.230 828.325 267.990 829.330 ;
        RECT 268.830 828.325 272.590 829.330 ;
        RECT 273.430 828.325 277.650 829.330 ;
        RECT 278.490 828.325 282.250 829.330 ;
        RECT 283.090 828.325 286.850 829.330 ;
        RECT 287.690 828.325 291.910 829.330 ;
        RECT 292.750 828.325 296.510 829.330 ;
        RECT 297.350 828.325 301.110 829.330 ;
        RECT 301.950 828.325 306.170 829.330 ;
        RECT 307.010 828.325 310.770 829.330 ;
        RECT 311.610 828.325 315.370 829.330 ;
        RECT 316.210 828.325 320.430 829.330 ;
        RECT 321.270 828.325 325.030 829.330 ;
        RECT 325.870 828.325 329.630 829.330 ;
        RECT 330.470 828.325 334.690 829.330 ;
        RECT 335.530 828.325 339.290 829.330 ;
        RECT 340.130 828.325 343.890 829.330 ;
        RECT 344.730 828.325 348.950 829.330 ;
        RECT 349.790 828.325 353.550 829.330 ;
        RECT 354.390 828.325 358.150 829.330 ;
        RECT 358.990 828.325 363.210 829.330 ;
        RECT 364.050 828.325 367.810 829.330 ;
        RECT 368.650 828.325 372.410 829.330 ;
        RECT 373.250 828.325 377.470 829.330 ;
        RECT 378.310 828.325 382.070 829.330 ;
        RECT 382.910 828.325 386.670 829.330 ;
        RECT 387.510 828.325 391.730 829.330 ;
        RECT 392.570 828.325 396.330 829.330 ;
        RECT 397.170 828.325 400.930 829.330 ;
        RECT 401.770 828.325 405.990 829.330 ;
        RECT 406.830 828.325 410.590 829.330 ;
        RECT 411.430 828.325 415.190 829.330 ;
        RECT 416.030 828.325 419.790 829.330 ;
        RECT 420.630 828.325 424.850 829.330 ;
        RECT 425.690 828.325 429.450 829.330 ;
        RECT 430.290 828.325 434.050 829.330 ;
        RECT 434.890 828.325 439.110 829.330 ;
        RECT 439.950 828.325 443.710 829.330 ;
        RECT 444.550 828.325 448.310 829.330 ;
        RECT 449.150 828.325 453.370 829.330 ;
        RECT 454.210 828.325 457.970 829.330 ;
        RECT 458.810 828.325 462.570 829.330 ;
        RECT 463.410 828.325 467.630 829.330 ;
        RECT 468.470 828.325 472.230 829.330 ;
        RECT 473.070 828.325 476.830 829.330 ;
        RECT 477.670 828.325 481.890 829.330 ;
        RECT 482.730 828.325 486.490 829.330 ;
        RECT 487.330 828.325 491.090 829.330 ;
        RECT 491.930 828.325 496.150 829.330 ;
        RECT 496.990 828.325 500.750 829.330 ;
        RECT 501.590 828.325 505.350 829.330 ;
        RECT 506.190 828.325 510.410 829.330 ;
        RECT 511.250 828.325 515.010 829.330 ;
        RECT 515.850 828.325 519.610 829.330 ;
        RECT 520.450 828.325 524.670 829.330 ;
        RECT 525.510 828.325 529.270 829.330 ;
        RECT 530.110 828.325 533.870 829.330 ;
        RECT 534.710 828.325 538.930 829.330 ;
        RECT 539.770 828.325 543.530 829.330 ;
        RECT 544.370 828.325 548.130 829.330 ;
        RECT 548.970 828.325 553.190 829.330 ;
        RECT 554.030 828.325 557.790 829.330 ;
        RECT 558.630 828.325 562.390 829.330 ;
        RECT 563.230 828.325 567.450 829.330 ;
        RECT 568.290 828.325 572.050 829.330 ;
        RECT 572.890 828.325 576.650 829.330 ;
        RECT 577.490 828.325 581.710 829.330 ;
        RECT 582.550 828.325 586.310 829.330 ;
        RECT 587.150 828.325 590.910 829.330 ;
        RECT 591.750 828.325 595.970 829.330 ;
        RECT 596.810 828.325 600.570 829.330 ;
        RECT 601.410 828.325 605.170 829.330 ;
        RECT 606.010 828.325 610.230 829.330 ;
        RECT 611.070 828.325 614.830 829.330 ;
        RECT 615.670 828.325 619.430 829.330 ;
        RECT 620.270 828.325 624.490 829.330 ;
        RECT 625.330 828.325 629.090 829.330 ;
        RECT 629.930 828.325 633.690 829.330 ;
        RECT 634.530 828.325 638.750 829.330 ;
        RECT 639.590 828.325 643.350 829.330 ;
        RECT 644.190 828.325 647.950 829.330 ;
        RECT 648.790 828.325 653.010 829.330 ;
        RECT 653.850 828.325 657.610 829.330 ;
        RECT 658.450 828.325 662.210 829.330 ;
        RECT 663.050 828.325 667.270 829.330 ;
        RECT 668.110 828.325 671.870 829.330 ;
        RECT 672.710 828.325 676.470 829.330 ;
        RECT 677.310 828.325 681.530 829.330 ;
        RECT 682.370 828.325 686.130 829.330 ;
        RECT 686.970 828.325 690.730 829.330 ;
        RECT 691.570 828.325 695.790 829.330 ;
        RECT 696.630 828.325 700.390 829.330 ;
        RECT 701.230 828.325 704.990 829.330 ;
        RECT 705.830 828.325 710.050 829.330 ;
        RECT 710.890 828.325 714.650 829.330 ;
        RECT 715.490 828.325 719.250 829.330 ;
        RECT 720.090 828.325 724.310 829.330 ;
        RECT 725.150 828.325 728.910 829.330 ;
        RECT 729.750 828.325 733.510 829.330 ;
        RECT 734.350 828.325 738.570 829.330 ;
        RECT 739.410 828.325 743.170 829.330 ;
        RECT 744.010 828.325 747.770 829.330 ;
        RECT 748.610 828.325 752.830 829.330 ;
        RECT 753.670 828.325 757.430 829.330 ;
        RECT 758.270 828.325 762.030 829.330 ;
        RECT 762.870 828.325 767.090 829.330 ;
        RECT 767.930 828.325 771.690 829.330 ;
        RECT 772.530 828.325 776.290 829.330 ;
        RECT 777.130 828.325 781.350 829.330 ;
        RECT 782.190 828.325 785.950 829.330 ;
        RECT 786.790 828.325 790.550 829.330 ;
        RECT 791.390 828.325 795.610 829.330 ;
        RECT 796.450 828.325 800.210 829.330 ;
        RECT 801.050 828.325 804.810 829.330 ;
        RECT 805.650 828.325 809.870 829.330 ;
        RECT 810.710 828.325 814.470 829.330 ;
        RECT 815.310 828.325 819.070 829.330 ;
        RECT 0.560 4.280 819.620 828.325 ;
        RECT 0.560 1.710 2.110 4.280 ;
        RECT 2.950 1.710 6.710 4.280 ;
        RECT 7.550 1.710 11.770 4.280 ;
        RECT 12.610 1.710 16.830 4.280 ;
        RECT 17.670 1.710 21.890 4.280 ;
        RECT 22.730 1.710 26.490 4.280 ;
        RECT 27.330 1.710 31.550 4.280 ;
        RECT 32.390 1.710 36.610 4.280 ;
        RECT 37.450 1.710 41.670 4.280 ;
        RECT 42.510 1.710 46.270 4.280 ;
        RECT 47.110 1.710 51.330 4.280 ;
        RECT 52.170 1.710 56.390 4.280 ;
        RECT 57.230 1.710 61.450 4.280 ;
        RECT 62.290 1.710 66.050 4.280 ;
        RECT 66.890 1.710 71.110 4.280 ;
        RECT 71.950 1.710 76.170 4.280 ;
        RECT 77.010 1.710 81.230 4.280 ;
        RECT 82.070 1.710 86.290 4.280 ;
        RECT 87.130 1.710 90.890 4.280 ;
        RECT 91.730 1.710 95.950 4.280 ;
        RECT 96.790 1.710 101.010 4.280 ;
        RECT 101.850 1.710 106.070 4.280 ;
        RECT 106.910 1.710 110.670 4.280 ;
        RECT 111.510 1.710 115.730 4.280 ;
        RECT 116.570 1.710 120.790 4.280 ;
        RECT 121.630 1.710 125.850 4.280 ;
        RECT 126.690 1.710 130.450 4.280 ;
        RECT 131.290 1.710 135.510 4.280 ;
        RECT 136.350 1.710 140.570 4.280 ;
        RECT 141.410 1.710 145.630 4.280 ;
        RECT 146.470 1.710 150.230 4.280 ;
        RECT 151.070 1.710 155.290 4.280 ;
        RECT 156.130 1.710 160.350 4.280 ;
        RECT 161.190 1.710 165.410 4.280 ;
        RECT 166.250 1.710 170.470 4.280 ;
        RECT 171.310 1.710 175.070 4.280 ;
        RECT 175.910 1.710 180.130 4.280 ;
        RECT 180.970 1.710 185.190 4.280 ;
        RECT 186.030 1.710 190.250 4.280 ;
        RECT 191.090 1.710 194.850 4.280 ;
        RECT 195.690 1.710 199.910 4.280 ;
        RECT 200.750 1.710 204.970 4.280 ;
        RECT 205.810 1.710 210.030 4.280 ;
        RECT 210.870 1.710 214.630 4.280 ;
        RECT 215.470 1.710 219.690 4.280 ;
        RECT 220.530 1.710 224.750 4.280 ;
        RECT 225.590 1.710 229.810 4.280 ;
        RECT 230.650 1.710 234.410 4.280 ;
        RECT 235.250 1.710 239.470 4.280 ;
        RECT 240.310 1.710 244.530 4.280 ;
        RECT 245.370 1.710 249.590 4.280 ;
        RECT 250.430 1.710 254.650 4.280 ;
        RECT 255.490 1.710 259.250 4.280 ;
        RECT 260.090 1.710 264.310 4.280 ;
        RECT 265.150 1.710 269.370 4.280 ;
        RECT 270.210 1.710 274.430 4.280 ;
        RECT 275.270 1.710 279.030 4.280 ;
        RECT 279.870 1.710 284.090 4.280 ;
        RECT 284.930 1.710 289.150 4.280 ;
        RECT 289.990 1.710 294.210 4.280 ;
        RECT 295.050 1.710 298.810 4.280 ;
        RECT 299.650 1.710 303.870 4.280 ;
        RECT 304.710 1.710 308.930 4.280 ;
        RECT 309.770 1.710 313.990 4.280 ;
        RECT 314.830 1.710 318.590 4.280 ;
        RECT 319.430 1.710 323.650 4.280 ;
        RECT 324.490 1.710 328.710 4.280 ;
        RECT 329.550 1.710 333.770 4.280 ;
        RECT 334.610 1.710 338.830 4.280 ;
        RECT 339.670 1.710 343.430 4.280 ;
        RECT 344.270 1.710 348.490 4.280 ;
        RECT 349.330 1.710 353.550 4.280 ;
        RECT 354.390 1.710 358.610 4.280 ;
        RECT 359.450 1.710 363.210 4.280 ;
        RECT 364.050 1.710 368.270 4.280 ;
        RECT 369.110 1.710 373.330 4.280 ;
        RECT 374.170 1.710 378.390 4.280 ;
        RECT 379.230 1.710 382.990 4.280 ;
        RECT 383.830 1.710 388.050 4.280 ;
        RECT 388.890 1.710 393.110 4.280 ;
        RECT 393.950 1.710 398.170 4.280 ;
        RECT 399.010 1.710 402.770 4.280 ;
        RECT 403.610 1.710 407.830 4.280 ;
        RECT 408.670 1.710 412.890 4.280 ;
        RECT 413.730 1.710 417.950 4.280 ;
        RECT 418.790 1.710 423.010 4.280 ;
        RECT 423.850 1.710 427.610 4.280 ;
        RECT 428.450 1.710 432.670 4.280 ;
        RECT 433.510 1.710 437.730 4.280 ;
        RECT 438.570 1.710 442.790 4.280 ;
        RECT 443.630 1.710 447.390 4.280 ;
        RECT 448.230 1.710 452.450 4.280 ;
        RECT 453.290 1.710 457.510 4.280 ;
        RECT 458.350 1.710 462.570 4.280 ;
        RECT 463.410 1.710 467.170 4.280 ;
        RECT 468.010 1.710 472.230 4.280 ;
        RECT 473.070 1.710 477.290 4.280 ;
        RECT 478.130 1.710 482.350 4.280 ;
        RECT 483.190 1.710 486.950 4.280 ;
        RECT 487.790 1.710 492.010 4.280 ;
        RECT 492.850 1.710 497.070 4.280 ;
        RECT 497.910 1.710 502.130 4.280 ;
        RECT 502.970 1.710 507.190 4.280 ;
        RECT 508.030 1.710 511.790 4.280 ;
        RECT 512.630 1.710 516.850 4.280 ;
        RECT 517.690 1.710 521.910 4.280 ;
        RECT 522.750 1.710 526.970 4.280 ;
        RECT 527.810 1.710 531.570 4.280 ;
        RECT 532.410 1.710 536.630 4.280 ;
        RECT 537.470 1.710 541.690 4.280 ;
        RECT 542.530 1.710 546.750 4.280 ;
        RECT 547.590 1.710 551.350 4.280 ;
        RECT 552.190 1.710 556.410 4.280 ;
        RECT 557.250 1.710 561.470 4.280 ;
        RECT 562.310 1.710 566.530 4.280 ;
        RECT 567.370 1.710 571.130 4.280 ;
        RECT 571.970 1.710 576.190 4.280 ;
        RECT 577.030 1.710 581.250 4.280 ;
        RECT 582.090 1.710 586.310 4.280 ;
        RECT 587.150 1.710 591.370 4.280 ;
        RECT 592.210 1.710 595.970 4.280 ;
        RECT 596.810 1.710 601.030 4.280 ;
        RECT 601.870 1.710 606.090 4.280 ;
        RECT 606.930 1.710 611.150 4.280 ;
        RECT 611.990 1.710 615.750 4.280 ;
        RECT 616.590 1.710 620.810 4.280 ;
        RECT 621.650 1.710 625.870 4.280 ;
        RECT 626.710 1.710 630.930 4.280 ;
        RECT 631.770 1.710 635.530 4.280 ;
        RECT 636.370 1.710 640.590 4.280 ;
        RECT 641.430 1.710 645.650 4.280 ;
        RECT 646.490 1.710 650.710 4.280 ;
        RECT 651.550 1.710 655.310 4.280 ;
        RECT 656.150 1.710 660.370 4.280 ;
        RECT 661.210 1.710 665.430 4.280 ;
        RECT 666.270 1.710 670.490 4.280 ;
        RECT 671.330 1.710 675.550 4.280 ;
        RECT 676.390 1.710 680.150 4.280 ;
        RECT 680.990 1.710 685.210 4.280 ;
        RECT 686.050 1.710 690.270 4.280 ;
        RECT 691.110 1.710 695.330 4.280 ;
        RECT 696.170 1.710 699.930 4.280 ;
        RECT 700.770 1.710 704.990 4.280 ;
        RECT 705.830 1.710 710.050 4.280 ;
        RECT 710.890 1.710 715.110 4.280 ;
        RECT 715.950 1.710 719.710 4.280 ;
        RECT 720.550 1.710 724.770 4.280 ;
        RECT 725.610 1.710 729.830 4.280 ;
        RECT 730.670 1.710 734.890 4.280 ;
        RECT 735.730 1.710 739.490 4.280 ;
        RECT 740.330 1.710 744.550 4.280 ;
        RECT 745.390 1.710 749.610 4.280 ;
        RECT 750.450 1.710 754.670 4.280 ;
        RECT 755.510 1.710 759.730 4.280 ;
        RECT 760.570 1.710 764.330 4.280 ;
        RECT 765.170 1.710 769.390 4.280 ;
        RECT 770.230 1.710 774.450 4.280 ;
        RECT 775.290 1.710 779.510 4.280 ;
        RECT 780.350 1.710 784.110 4.280 ;
        RECT 784.950 1.710 789.170 4.280 ;
        RECT 790.010 1.710 794.230 4.280 ;
        RECT 795.070 1.710 799.290 4.280 ;
        RECT 800.130 1.710 803.890 4.280 ;
        RECT 804.730 1.710 808.950 4.280 ;
        RECT 809.790 1.710 814.010 4.280 ;
        RECT 814.850 1.710 819.070 4.280 ;
      LAYER met3 ;
        RECT 0.985 814.320 817.885 821.605 ;
        RECT 0.985 812.920 817.485 814.320 ;
        RECT 0.985 810.920 817.885 812.920 ;
        RECT 4.400 809.520 817.885 810.920 ;
        RECT 0.985 802.080 817.885 809.520 ;
        RECT 0.985 800.680 817.485 802.080 ;
        RECT 0.985 795.960 817.885 800.680 ;
        RECT 4.400 794.560 817.885 795.960 ;
        RECT 0.985 790.520 817.885 794.560 ;
        RECT 0.985 789.120 817.485 790.520 ;
        RECT 0.985 781.680 817.885 789.120 ;
        RECT 4.400 780.280 817.885 781.680 ;
        RECT 0.985 778.280 817.885 780.280 ;
        RECT 0.985 776.880 817.485 778.280 ;
        RECT 0.985 766.720 817.885 776.880 ;
        RECT 4.400 766.040 817.885 766.720 ;
        RECT 4.400 765.320 817.485 766.040 ;
        RECT 0.985 764.640 817.485 765.320 ;
        RECT 0.985 753.800 817.885 764.640 ;
        RECT 0.985 752.440 817.485 753.800 ;
        RECT 4.400 752.400 817.485 752.440 ;
        RECT 4.400 751.040 817.885 752.400 ;
        RECT 0.985 742.240 817.885 751.040 ;
        RECT 0.985 740.840 817.485 742.240 ;
        RECT 0.985 737.480 817.885 740.840 ;
        RECT 4.400 736.080 817.885 737.480 ;
        RECT 0.985 730.000 817.885 736.080 ;
        RECT 0.985 728.600 817.485 730.000 ;
        RECT 0.985 723.200 817.885 728.600 ;
        RECT 4.400 721.800 817.885 723.200 ;
        RECT 0.985 717.760 817.885 721.800 ;
        RECT 0.985 716.360 817.485 717.760 ;
        RECT 0.985 708.240 817.885 716.360 ;
        RECT 4.400 706.840 817.885 708.240 ;
        RECT 0.985 705.520 817.885 706.840 ;
        RECT 0.985 704.120 817.485 705.520 ;
        RECT 0.985 693.960 817.885 704.120 ;
        RECT 4.400 692.560 817.485 693.960 ;
        RECT 0.985 681.720 817.885 692.560 ;
        RECT 0.985 680.320 817.485 681.720 ;
        RECT 0.985 679.000 817.885 680.320 ;
        RECT 4.400 677.600 817.885 679.000 ;
        RECT 0.985 669.480 817.885 677.600 ;
        RECT 0.985 668.080 817.485 669.480 ;
        RECT 0.985 664.720 817.885 668.080 ;
        RECT 4.400 663.320 817.885 664.720 ;
        RECT 0.985 657.240 817.885 663.320 ;
        RECT 0.985 655.840 817.485 657.240 ;
        RECT 0.985 649.760 817.885 655.840 ;
        RECT 4.400 648.360 817.885 649.760 ;
        RECT 0.985 645.680 817.885 648.360 ;
        RECT 0.985 644.280 817.485 645.680 ;
        RECT 0.985 635.480 817.885 644.280 ;
        RECT 4.400 634.080 817.885 635.480 ;
        RECT 0.985 633.440 817.885 634.080 ;
        RECT 0.985 632.040 817.485 633.440 ;
        RECT 0.985 621.200 817.885 632.040 ;
        RECT 0.985 620.520 817.485 621.200 ;
        RECT 4.400 619.800 817.485 620.520 ;
        RECT 4.400 619.120 817.885 619.800 ;
        RECT 0.985 608.960 817.885 619.120 ;
        RECT 0.985 607.560 817.485 608.960 ;
        RECT 0.985 606.240 817.885 607.560 ;
        RECT 4.400 604.840 817.885 606.240 ;
        RECT 0.985 597.400 817.885 604.840 ;
        RECT 0.985 596.000 817.485 597.400 ;
        RECT 0.985 591.280 817.885 596.000 ;
        RECT 4.400 589.880 817.885 591.280 ;
        RECT 0.985 585.160 817.885 589.880 ;
        RECT 0.985 583.760 817.485 585.160 ;
        RECT 0.985 577.000 817.885 583.760 ;
        RECT 4.400 575.600 817.885 577.000 ;
        RECT 0.985 572.920 817.885 575.600 ;
        RECT 0.985 571.520 817.485 572.920 ;
        RECT 0.985 562.720 817.885 571.520 ;
        RECT 4.400 561.360 817.885 562.720 ;
        RECT 4.400 561.320 817.485 561.360 ;
        RECT 0.985 559.960 817.485 561.320 ;
        RECT 0.985 549.120 817.885 559.960 ;
        RECT 0.985 547.760 817.485 549.120 ;
        RECT 4.400 547.720 817.485 547.760 ;
        RECT 4.400 546.360 817.885 547.720 ;
        RECT 0.985 536.880 817.885 546.360 ;
        RECT 0.985 535.480 817.485 536.880 ;
        RECT 0.985 533.480 817.885 535.480 ;
        RECT 4.400 532.080 817.885 533.480 ;
        RECT 0.985 524.640 817.885 532.080 ;
        RECT 0.985 523.240 817.485 524.640 ;
        RECT 0.985 518.520 817.885 523.240 ;
        RECT 4.400 517.120 817.885 518.520 ;
        RECT 0.985 513.080 817.885 517.120 ;
        RECT 0.985 511.680 817.485 513.080 ;
        RECT 0.985 504.240 817.885 511.680 ;
        RECT 4.400 502.840 817.885 504.240 ;
        RECT 0.985 500.840 817.885 502.840 ;
        RECT 0.985 499.440 817.485 500.840 ;
        RECT 0.985 489.280 817.885 499.440 ;
        RECT 4.400 488.600 817.885 489.280 ;
        RECT 4.400 487.880 817.485 488.600 ;
        RECT 0.985 487.200 817.485 487.880 ;
        RECT 0.985 476.360 817.885 487.200 ;
        RECT 0.985 475.000 817.485 476.360 ;
        RECT 4.400 474.960 817.485 475.000 ;
        RECT 4.400 473.600 817.885 474.960 ;
        RECT 0.985 464.800 817.885 473.600 ;
        RECT 0.985 463.400 817.485 464.800 ;
        RECT 0.985 460.040 817.885 463.400 ;
        RECT 4.400 458.640 817.885 460.040 ;
        RECT 0.985 452.560 817.885 458.640 ;
        RECT 0.985 451.160 817.485 452.560 ;
        RECT 0.985 445.760 817.885 451.160 ;
        RECT 4.400 444.360 817.885 445.760 ;
        RECT 0.985 440.320 817.885 444.360 ;
        RECT 0.985 438.920 817.485 440.320 ;
        RECT 0.985 430.800 817.885 438.920 ;
        RECT 4.400 429.400 817.885 430.800 ;
        RECT 0.985 428.080 817.885 429.400 ;
        RECT 0.985 426.680 817.485 428.080 ;
        RECT 0.985 416.520 817.885 426.680 ;
        RECT 4.400 415.120 817.485 416.520 ;
        RECT 0.985 404.280 817.885 415.120 ;
        RECT 0.985 402.880 817.485 404.280 ;
        RECT 0.985 401.560 817.885 402.880 ;
        RECT 4.400 400.160 817.885 401.560 ;
        RECT 0.985 392.040 817.885 400.160 ;
        RECT 0.985 390.640 817.485 392.040 ;
        RECT 0.985 387.280 817.885 390.640 ;
        RECT 4.400 385.880 817.885 387.280 ;
        RECT 0.985 379.800 817.885 385.880 ;
        RECT 0.985 378.400 817.485 379.800 ;
        RECT 0.985 372.320 817.885 378.400 ;
        RECT 4.400 370.920 817.885 372.320 ;
        RECT 0.985 368.240 817.885 370.920 ;
        RECT 0.985 366.840 817.485 368.240 ;
        RECT 0.985 358.040 817.885 366.840 ;
        RECT 4.400 356.640 817.885 358.040 ;
        RECT 0.985 356.000 817.885 356.640 ;
        RECT 0.985 354.600 817.485 356.000 ;
        RECT 0.985 343.760 817.885 354.600 ;
        RECT 0.985 343.080 817.485 343.760 ;
        RECT 4.400 342.360 817.485 343.080 ;
        RECT 4.400 341.680 817.885 342.360 ;
        RECT 0.985 331.520 817.885 341.680 ;
        RECT 0.985 330.120 817.485 331.520 ;
        RECT 0.985 328.800 817.885 330.120 ;
        RECT 4.400 327.400 817.885 328.800 ;
        RECT 0.985 319.960 817.885 327.400 ;
        RECT 0.985 318.560 817.485 319.960 ;
        RECT 0.985 313.840 817.885 318.560 ;
        RECT 4.400 312.440 817.885 313.840 ;
        RECT 0.985 307.720 817.885 312.440 ;
        RECT 0.985 306.320 817.485 307.720 ;
        RECT 0.985 299.560 817.885 306.320 ;
        RECT 4.400 298.160 817.885 299.560 ;
        RECT 0.985 295.480 817.885 298.160 ;
        RECT 0.985 294.080 817.485 295.480 ;
        RECT 0.985 285.280 817.885 294.080 ;
        RECT 4.400 283.920 817.885 285.280 ;
        RECT 4.400 283.880 817.485 283.920 ;
        RECT 0.985 282.520 817.485 283.880 ;
        RECT 0.985 271.680 817.885 282.520 ;
        RECT 0.985 270.320 817.485 271.680 ;
        RECT 4.400 270.280 817.485 270.320 ;
        RECT 4.400 268.920 817.885 270.280 ;
        RECT 0.985 259.440 817.885 268.920 ;
        RECT 0.985 258.040 817.485 259.440 ;
        RECT 0.985 256.040 817.885 258.040 ;
        RECT 4.400 254.640 817.885 256.040 ;
        RECT 0.985 247.200 817.885 254.640 ;
        RECT 0.985 245.800 817.485 247.200 ;
        RECT 0.985 241.080 817.885 245.800 ;
        RECT 4.400 239.680 817.885 241.080 ;
        RECT 0.985 235.640 817.885 239.680 ;
        RECT 0.985 234.240 817.485 235.640 ;
        RECT 0.985 226.800 817.885 234.240 ;
        RECT 4.400 225.400 817.885 226.800 ;
        RECT 0.985 223.400 817.885 225.400 ;
        RECT 0.985 222.000 817.485 223.400 ;
        RECT 0.985 211.840 817.885 222.000 ;
        RECT 4.400 211.160 817.885 211.840 ;
        RECT 4.400 210.440 817.485 211.160 ;
        RECT 0.985 209.760 817.485 210.440 ;
        RECT 0.985 198.920 817.885 209.760 ;
        RECT 0.985 197.560 817.485 198.920 ;
        RECT 4.400 197.520 817.485 197.560 ;
        RECT 4.400 196.160 817.885 197.520 ;
        RECT 0.985 187.360 817.885 196.160 ;
        RECT 0.985 185.960 817.485 187.360 ;
        RECT 0.985 182.600 817.885 185.960 ;
        RECT 4.400 181.200 817.885 182.600 ;
        RECT 0.985 175.120 817.885 181.200 ;
        RECT 0.985 173.720 817.485 175.120 ;
        RECT 0.985 168.320 817.885 173.720 ;
        RECT 4.400 166.920 817.885 168.320 ;
        RECT 0.985 162.880 817.885 166.920 ;
        RECT 0.985 161.480 817.485 162.880 ;
        RECT 0.985 153.360 817.885 161.480 ;
        RECT 4.400 151.960 817.885 153.360 ;
        RECT 0.985 150.640 817.885 151.960 ;
        RECT 0.985 149.240 817.485 150.640 ;
        RECT 0.985 139.080 817.885 149.240 ;
        RECT 4.400 137.680 817.485 139.080 ;
        RECT 0.985 126.840 817.885 137.680 ;
        RECT 0.985 125.440 817.485 126.840 ;
        RECT 0.985 124.120 817.885 125.440 ;
        RECT 4.400 122.720 817.885 124.120 ;
        RECT 0.985 114.600 817.885 122.720 ;
        RECT 0.985 113.200 817.485 114.600 ;
        RECT 0.985 109.840 817.885 113.200 ;
        RECT 4.400 108.440 817.885 109.840 ;
        RECT 0.985 102.360 817.885 108.440 ;
        RECT 0.985 100.960 817.485 102.360 ;
        RECT 0.985 94.880 817.885 100.960 ;
        RECT 4.400 93.480 817.885 94.880 ;
        RECT 0.985 90.800 817.885 93.480 ;
        RECT 0.985 89.400 817.485 90.800 ;
        RECT 0.985 80.600 817.885 89.400 ;
        RECT 4.400 79.200 817.885 80.600 ;
        RECT 0.985 78.560 817.885 79.200 ;
        RECT 0.985 77.160 817.485 78.560 ;
        RECT 0.985 66.320 817.885 77.160 ;
        RECT 0.985 65.640 817.485 66.320 ;
        RECT 4.400 64.920 817.485 65.640 ;
        RECT 4.400 64.240 817.885 64.920 ;
        RECT 0.985 54.080 817.885 64.240 ;
        RECT 0.985 52.680 817.485 54.080 ;
        RECT 0.985 51.360 817.885 52.680 ;
        RECT 4.400 49.960 817.885 51.360 ;
        RECT 0.985 42.520 817.885 49.960 ;
        RECT 0.985 41.120 817.485 42.520 ;
        RECT 0.985 36.400 817.885 41.120 ;
        RECT 4.400 35.000 817.885 36.400 ;
        RECT 0.985 30.280 817.885 35.000 ;
        RECT 0.985 28.880 817.485 30.280 ;
        RECT 0.985 22.120 817.885 28.880 ;
        RECT 4.400 20.720 817.885 22.120 ;
        RECT 0.985 18.040 817.885 20.720 ;
        RECT 0.985 16.640 817.485 18.040 ;
        RECT 0.985 7.840 817.885 16.640 ;
        RECT 4.400 6.480 817.885 7.840 ;
        RECT 4.400 6.440 817.485 6.480 ;
        RECT 0.985 5.080 817.485 6.440 ;
        RECT 0.985 2.895 817.885 5.080 ;
      LAYER met4 ;
        RECT 1.215 10.240 20.640 820.585 ;
        RECT 23.040 10.240 97.440 820.585 ;
        RECT 99.840 10.240 174.240 820.585 ;
        RECT 176.640 10.240 251.040 820.585 ;
        RECT 253.440 10.240 327.840 820.585 ;
        RECT 330.240 10.240 404.640 820.585 ;
        RECT 407.040 10.240 481.440 820.585 ;
        RECT 483.840 10.240 558.240 820.585 ;
        RECT 560.640 10.240 635.040 820.585 ;
        RECT 637.440 10.240 711.840 820.585 ;
        RECT 714.240 10.240 788.145 820.585 ;
        RECT 1.215 2.895 788.145 10.240 ;
  END
END user_proj
END LIBRARY

