magic
tech sky130A
magscale 1 2
timestamp 1638672285
<< locali >>
rect 269221 700519 269255 700553
rect 269221 700485 269405 700519
rect 281365 700111 281399 700553
rect 36001 697595 36035 699329
rect 65625 698343 65659 699329
rect 70409 698411 70443 699329
rect 80161 698479 80195 699329
rect 85313 698547 85347 699329
rect 100033 698615 100067 699329
rect 109877 698683 109911 699329
rect 158821 698887 158855 699329
rect 168849 699091 168883 699329
rect 173725 699023 173759 699329
rect 188445 699227 188479 699329
rect 379529 699295 379563 699465
rect 367109 697527 367143 697833
rect 371893 697663 371927 697765
rect 386245 697731 386279 699465
rect 394157 699159 394191 699465
rect 408877 698955 408911 699465
rect 423689 698819 423723 699465
rect 438317 698751 438351 699465
rect 521853 697663 521887 699465
rect 367235 697561 367293 697595
rect 247969 663 248003 765
rect 340889 663 340923 765
rect 212123 561 212273 595
rect 6193 391 6227 561
rect 252385 323 252419 561
rect 254777 391 254811 561
rect 280721 255 280755 561
rect 310253 187 310287 561
rect 312645 323 312679 561
rect 335921 391 335955 561
rect 336105 119 336139 561
rect 355241 255 355275 561
rect 364809 391 364843 561
rect 365085 187 365119 561
rect 366097 527 366131 697
rect 370697 595 370731 697
rect 368213 119 368247 561
rect 370605 51 370639 561
rect 372077 323 372111 765
rect 372813 527 372847 697
rect 383117 595 383151 697
rect 404737 663 404771 901
rect 389465 459 389499 561
rect 404495 561 404829 595
rect 389373 119 389407 221
rect 390201 119 390235 357
rect 393789 119 393823 493
rect 396181 119 396215 357
rect 398021 255 398055 561
rect 404921 255 404955 629
rect 406485 323 406519 833
rect 406577 255 406611 765
rect 413753 663 413787 1309
rect 417157 663 417191 1037
rect 411453 459 411487 629
rect 418813 459 418847 765
rect 421665 595 421699 833
rect 422861 595 422895 697
rect 423781 595 423815 765
rect 424701 595 424735 765
rect 426357 527 426391 1309
rect 429025 527 429059 1037
rect 430405 459 430439 969
rect 432521 663 432555 833
rect 437949 663 437983 901
rect 435741 255 435775 493
rect 431785 221 431877 255
rect 431785 119 431819 221
rect 439881 51 439915 833
rect 442181 595 442215 1037
rect 443653 663 443687 765
rect 443837 595 443871 969
rect 448989 663 449023 969
rect 450001 595 450035 697
rect 451289 595 451323 697
rect 452393 595 452427 833
rect 453497 527 453531 765
rect 454693 663 454727 765
rect 454509 187 454543 561
rect 454785 459 454819 629
rect 455337 595 455371 1037
rect 455429 459 455463 901
rect 455889 119 455923 561
rect 456533 459 456567 1037
rect 458005 663 458039 1105
rect 458189 663 458223 765
rect 460213 663 460247 1173
rect 461811 901 461995 935
rect 461961 731 461995 901
rect 462237 663 462271 969
rect 469597 255 469631 697
rect 472265 663 472299 1105
rect 472817 663 472851 1037
rect 474565 663 474599 1173
rect 469781 323 469815 493
rect 474933 391 474967 629
rect 475117 595 475151 765
rect 476221 595 476255 1105
rect 476589 595 476623 969
rect 481465 663 481499 901
rect 481741 323 481775 561
rect 482845 323 482879 969
rect 483765 663 483799 1037
rect 486433 595 486467 833
rect 487721 663 487755 969
rect 489871 697 490021 731
rect 491125 663 491159 1105
rect 494437 663 494471 1241
rect 493275 629 493643 663
rect 493609 595 493643 629
rect 495357 595 495391 1173
rect 496737 595 496771 1105
rect 499405 595 499439 1037
rect 493459 493 493701 527
rect 492781 255 492815 357
rect 498209 51 498243 561
rect 502349 459 502383 1037
rect 505753 663 505787 901
rect 507317 527 507351 969
rect 509249 663 509283 969
rect 509709 663 509743 1037
rect 510261 391 510295 1241
rect 511273 663 511307 1173
rect 512469 663 512503 1105
rect 513297 663 513331 833
rect 515873 663 515907 765
rect 517069 663 517103 1037
rect 519369 663 519403 1105
rect 521853 663 521887 901
rect 524153 595 524187 765
rect 525073 459 525107 697
rect 525165 459 525199 969
rect 528845 459 528879 629
rect 530133 595 530167 833
rect 531881 595 531915 901
rect 533721 595 533755 1037
rect 535837 663 535871 1105
rect 536481 663 536515 833
rect 540805 663 540839 765
rect 543197 255 543231 629
rect 545497 391 545531 629
rect 548533 527 548567 697
rect 548901 527 548935 833
rect 549085 527 549119 901
rect 551201 595 551235 765
rect 555801 663 555835 1037
rect 558009 527 558043 1105
rect 558745 527 558779 969
rect 562241 867 562275 1173
rect 562609 459 562643 901
rect 561723 357 561965 391
<< viali >>
rect 269221 700553 269255 700587
rect 281365 700553 281399 700587
rect 269405 700485 269439 700519
rect 281365 700077 281399 700111
rect 379529 699465 379563 699499
rect 36001 699329 36035 699363
rect 65625 699329 65659 699363
rect 70409 699329 70443 699363
rect 80161 699329 80195 699363
rect 85313 699329 85347 699363
rect 100033 699329 100067 699363
rect 109877 699329 109911 699363
rect 158821 699329 158855 699363
rect 168849 699329 168883 699363
rect 168849 699057 168883 699091
rect 173725 699329 173759 699363
rect 188445 699329 188479 699363
rect 379529 699261 379563 699295
rect 386245 699465 386279 699499
rect 188445 699193 188479 699227
rect 173725 698989 173759 699023
rect 158821 698853 158855 698887
rect 109877 698649 109911 698683
rect 100033 698581 100067 698615
rect 85313 698513 85347 698547
rect 80161 698445 80195 698479
rect 70409 698377 70443 698411
rect 65625 698309 65659 698343
rect 36001 697561 36035 697595
rect 367109 697833 367143 697867
rect 371893 697765 371927 697799
rect 394157 699465 394191 699499
rect 394157 699125 394191 699159
rect 408877 699465 408911 699499
rect 408877 698921 408911 698955
rect 423689 699465 423723 699499
rect 423689 698785 423723 698819
rect 438317 699465 438351 699499
rect 438317 698717 438351 698751
rect 521853 699465 521887 699499
rect 386245 697697 386279 697731
rect 371893 697629 371927 697663
rect 521853 697629 521887 697663
rect 367201 697561 367235 697595
rect 367293 697561 367327 697595
rect 367109 697493 367143 697527
rect 413753 1309 413787 1343
rect 404737 901 404771 935
rect 247969 765 248003 799
rect 247969 629 248003 663
rect 340889 765 340923 799
rect 372077 765 372111 799
rect 340889 629 340923 663
rect 366097 697 366131 731
rect 6193 561 6227 595
rect 212089 561 212123 595
rect 212273 561 212307 595
rect 252385 561 252419 595
rect 6193 357 6227 391
rect 254777 561 254811 595
rect 254777 357 254811 391
rect 280721 561 280755 595
rect 252385 289 252419 323
rect 280721 221 280755 255
rect 310253 561 310287 595
rect 312645 561 312679 595
rect 335921 561 335955 595
rect 335921 357 335955 391
rect 336105 561 336139 595
rect 312645 289 312679 323
rect 310253 153 310287 187
rect 355241 561 355275 595
rect 364809 561 364843 595
rect 364809 357 364843 391
rect 365085 561 365119 595
rect 355241 221 355275 255
rect 370697 697 370731 731
rect 366097 493 366131 527
rect 368213 561 368247 595
rect 365085 153 365119 187
rect 336105 85 336139 119
rect 368213 85 368247 119
rect 370605 561 370639 595
rect 370697 561 370731 595
rect 372813 697 372847 731
rect 383117 697 383151 731
rect 406485 833 406519 867
rect 404737 629 404771 663
rect 404921 629 404955 663
rect 383117 561 383151 595
rect 389465 561 389499 595
rect 372813 493 372847 527
rect 398021 561 398055 595
rect 404461 561 404495 595
rect 404829 561 404863 595
rect 389465 425 389499 459
rect 393789 493 393823 527
rect 372077 289 372111 323
rect 390201 357 390235 391
rect 389373 221 389407 255
rect 389373 85 389407 119
rect 390201 85 390235 119
rect 393789 85 393823 119
rect 396181 357 396215 391
rect 398021 221 398055 255
rect 406485 289 406519 323
rect 406577 765 406611 799
rect 404921 221 404955 255
rect 426357 1309 426391 1343
rect 411453 629 411487 663
rect 413753 629 413787 663
rect 417157 1037 417191 1071
rect 421665 833 421699 867
rect 417157 629 417191 663
rect 418813 765 418847 799
rect 411453 425 411487 459
rect 423781 765 423815 799
rect 421665 561 421699 595
rect 422861 697 422895 731
rect 422861 561 422895 595
rect 423781 561 423815 595
rect 424701 765 424735 799
rect 424701 561 424735 595
rect 494437 1241 494471 1275
rect 460213 1173 460247 1207
rect 458005 1105 458039 1139
rect 426357 493 426391 527
rect 429025 1037 429059 1071
rect 442181 1037 442215 1071
rect 429025 493 429059 527
rect 430405 969 430439 1003
rect 418813 425 418847 459
rect 437949 901 437983 935
rect 432521 833 432555 867
rect 432521 629 432555 663
rect 437949 629 437983 663
rect 439881 833 439915 867
rect 430405 425 430439 459
rect 435741 493 435775 527
rect 406577 221 406611 255
rect 431877 221 431911 255
rect 435741 221 435775 255
rect 396181 85 396215 119
rect 431785 85 431819 119
rect 370605 17 370639 51
rect 455337 1037 455371 1071
rect 443837 969 443871 1003
rect 443653 765 443687 799
rect 443653 629 443687 663
rect 442181 561 442215 595
rect 448989 969 449023 1003
rect 452393 833 452427 867
rect 448989 629 449023 663
rect 450001 697 450035 731
rect 443837 561 443871 595
rect 450001 561 450035 595
rect 451289 697 451323 731
rect 451289 561 451323 595
rect 452393 561 452427 595
rect 453497 765 453531 799
rect 454693 765 454727 799
rect 454693 629 454727 663
rect 454785 629 454819 663
rect 453497 493 453531 527
rect 454509 561 454543 595
rect 456533 1037 456567 1071
rect 455337 561 455371 595
rect 455429 901 455463 935
rect 454785 425 454819 459
rect 455429 425 455463 459
rect 455889 561 455923 595
rect 454509 153 454543 187
rect 458005 629 458039 663
rect 458189 765 458223 799
rect 458189 629 458223 663
rect 474565 1173 474599 1207
rect 472265 1105 472299 1139
rect 462237 969 462271 1003
rect 461777 901 461811 935
rect 461961 697 461995 731
rect 460213 629 460247 663
rect 462237 629 462271 663
rect 469597 697 469631 731
rect 456533 425 456567 459
rect 472265 629 472299 663
rect 472817 1037 472851 1071
rect 472817 629 472851 663
rect 476221 1105 476255 1139
rect 475117 765 475151 799
rect 474565 629 474599 663
rect 474933 629 474967 663
rect 469781 493 469815 527
rect 475117 561 475151 595
rect 491125 1105 491159 1139
rect 483765 1037 483799 1071
rect 476221 561 476255 595
rect 476589 969 476623 1003
rect 482845 969 482879 1003
rect 481465 901 481499 935
rect 481465 629 481499 663
rect 476589 561 476623 595
rect 481741 561 481775 595
rect 474933 357 474967 391
rect 469781 289 469815 323
rect 481741 289 481775 323
rect 487721 969 487755 1003
rect 483765 629 483799 663
rect 486433 833 486467 867
rect 489837 697 489871 731
rect 490021 697 490055 731
rect 487721 629 487755 663
rect 510261 1241 510295 1275
rect 491125 629 491159 663
rect 493241 629 493275 663
rect 494437 629 494471 663
rect 495357 1173 495391 1207
rect 486433 561 486467 595
rect 493609 561 493643 595
rect 495357 561 495391 595
rect 496737 1105 496771 1139
rect 499405 1037 499439 1071
rect 496737 561 496771 595
rect 498209 561 498243 595
rect 499405 561 499439 595
rect 502349 1037 502383 1071
rect 493425 493 493459 527
rect 493701 493 493735 527
rect 482845 289 482879 323
rect 492781 357 492815 391
rect 469597 221 469631 255
rect 492781 221 492815 255
rect 455889 85 455923 119
rect 439881 17 439915 51
rect 509709 1037 509743 1071
rect 507317 969 507351 1003
rect 505753 901 505787 935
rect 505753 629 505787 663
rect 509249 969 509283 1003
rect 509249 629 509283 663
rect 509709 629 509743 663
rect 507317 493 507351 527
rect 502349 425 502383 459
rect 511273 1173 511307 1207
rect 562241 1173 562275 1207
rect 511273 629 511307 663
rect 512469 1105 512503 1139
rect 519369 1105 519403 1139
rect 517069 1037 517103 1071
rect 512469 629 512503 663
rect 513297 833 513331 867
rect 513297 629 513331 663
rect 515873 765 515907 799
rect 515873 629 515907 663
rect 517069 629 517103 663
rect 535837 1105 535871 1139
rect 533721 1037 533755 1071
rect 525165 969 525199 1003
rect 519369 629 519403 663
rect 521853 901 521887 935
rect 521853 629 521887 663
rect 524153 765 524187 799
rect 524153 561 524187 595
rect 525073 697 525107 731
rect 525073 425 525107 459
rect 531881 901 531915 935
rect 530133 833 530167 867
rect 525165 425 525199 459
rect 528845 629 528879 663
rect 530133 561 530167 595
rect 531881 561 531915 595
rect 558009 1105 558043 1139
rect 555801 1037 555835 1071
rect 549085 901 549119 935
rect 535837 629 535871 663
rect 536481 833 536515 867
rect 548901 833 548935 867
rect 536481 629 536515 663
rect 540805 765 540839 799
rect 548533 697 548567 731
rect 540805 629 540839 663
rect 543197 629 543231 663
rect 533721 561 533755 595
rect 528845 425 528879 459
rect 510261 357 510295 391
rect 545497 629 545531 663
rect 548533 493 548567 527
rect 548901 493 548935 527
rect 551201 765 551235 799
rect 555801 629 555835 663
rect 551201 561 551235 595
rect 549085 493 549119 527
rect 558009 493 558043 527
rect 558745 969 558779 1003
rect 562241 833 562275 867
rect 562609 901 562643 935
rect 558745 493 558779 527
rect 562609 425 562643 459
rect 545497 357 545531 391
rect 561689 357 561723 391
rect 561965 357 561999 391
rect 543197 221 543231 255
rect 498209 17 498243 51
<< metal1 >>
rect 235442 703808 235448 703860
rect 235500 703848 235506 703860
rect 300854 703848 300860 703860
rect 235500 703820 300860 703848
rect 235500 703808 235506 703820
rect 300854 703808 300860 703820
rect 300912 703808 300918 703860
rect 271782 703740 271788 703792
rect 271840 703780 271846 703792
rect 364702 703780 364708 703792
rect 271840 703752 364708 703780
rect 271840 703740 271846 703752
rect 364702 703740 364708 703752
rect 364760 703740 364766 703792
rect 170490 703672 170496 703724
rect 170548 703712 170554 703724
rect 315482 703712 315488 703724
rect 170548 703684 315488 703712
rect 170548 703672 170554 703684
rect 315482 703672 315488 703684
rect 315540 703672 315546 703724
rect 257246 703604 257252 703656
rect 257304 703644 257310 703656
rect 429654 703644 429660 703656
rect 257304 703616 429660 703644
rect 257304 703604 257310 703616
rect 429654 703604 429660 703616
rect 429712 703604 429718 703656
rect 242434 703536 242440 703588
rect 242492 703576 242498 703588
rect 494422 703576 494428 703588
rect 242492 703548 494428 703576
rect 242492 703536 242498 703548
rect 494422 703536 494428 703548
rect 494480 703536 494486 703588
rect 227622 703468 227628 703520
rect 227680 703508 227686 703520
rect 503898 703508 503904 703520
rect 227680 703480 503904 703508
rect 227680 703468 227686 703480
rect 503898 703468 503904 703480
rect 503956 703468 503962 703520
rect 105446 703400 105452 703452
rect 105504 703440 105510 703452
rect 330294 703440 330300 703452
rect 105504 703412 330300 703440
rect 105504 703400 105510 703412
rect 330294 703400 330300 703412
rect 330352 703400 330358 703452
rect 40494 703332 40500 703384
rect 40552 703372 40558 703384
rect 345014 703372 345020 703384
rect 40552 703344 345020 703372
rect 40552 703332 40558 703344
rect 345014 703332 345020 703344
rect 345072 703332 345078 703384
rect 1578 703264 1584 703316
rect 1636 703304 1642 703316
rect 359734 703304 359740 703316
rect 1636 703276 359740 703304
rect 1636 703264 1642 703276
rect 359734 703264 359740 703276
rect 359792 703264 359798 703316
rect 212994 703196 213000 703248
rect 213052 703236 213058 703248
rect 576394 703236 576400 703248
rect 213052 703208 576400 703236
rect 213052 703196 213058 703208
rect 576394 703196 576400 703208
rect 576452 703196 576458 703248
rect 1670 703128 1676 703180
rect 1728 703168 1734 703180
rect 374454 703168 374460 703180
rect 1728 703140 374460 703168
rect 1728 703128 1734 703140
rect 374454 703128 374460 703140
rect 374512 703128 374518 703180
rect 198274 703060 198280 703112
rect 198332 703100 198338 703112
rect 575014 703100 575020 703112
rect 198332 703072 575020 703100
rect 198332 703060 198338 703072
rect 575014 703060 575020 703072
rect 575072 703060 575078 703112
rect 1762 702992 1768 703044
rect 1820 703032 1826 703044
rect 389174 703032 389180 703044
rect 1820 703004 389180 703032
rect 1820 702992 1826 703004
rect 389174 702992 389180 703004
rect 389232 702992 389238 703044
rect 183370 702924 183376 702976
rect 183428 702964 183434 702976
rect 573634 702964 573640 702976
rect 183428 702936 573640 702964
rect 183428 702924 183434 702936
rect 573634 702924 573640 702936
rect 573692 702924 573698 702976
rect 1854 702856 1860 702908
rect 1912 702896 1918 702908
rect 403894 702896 403900 702908
rect 1912 702868 403900 702896
rect 1912 702856 1918 702868
rect 403894 702856 403900 702868
rect 403952 702856 403958 702908
rect 139302 702788 139308 702840
rect 139360 702828 139366 702840
rect 572162 702828 572168 702840
rect 139360 702800 572168 702828
rect 139360 702788 139366 702800
rect 572162 702788 572168 702800
rect 572220 702788 572226 702840
rect 2498 702720 2504 702772
rect 2556 702760 2562 702772
rect 448146 702760 448152 702772
rect 2556 702732 448152 702760
rect 2556 702720 2562 702732
rect 448146 702720 448152 702732
rect 448204 702720 448210 702772
rect 474 702652 480 702704
rect 532 702692 538 702704
rect 477586 702692 477592 702704
rect 532 702664 477592 702692
rect 532 702652 538 702664
rect 477586 702652 477592 702664
rect 477644 702652 477650 702704
rect 290 702584 296 702636
rect 348 702624 354 702636
rect 507118 702624 507124 702636
rect 348 702596 507124 702624
rect 348 702584 354 702596
rect 507118 702584 507124 702596
rect 507176 702584 507182 702636
rect 14 702516 20 702568
rect 72 702556 78 702568
rect 536834 702556 536840 702568
rect 72 702528 536840 702556
rect 72 702516 78 702528
rect 536834 702516 536840 702528
rect 536892 702516 536898 702568
rect 21450 702448 21456 702500
rect 21508 702488 21514 702500
rect 576118 702488 576124 702500
rect 21508 702460 576124 702488
rect 21508 702448 21514 702460
rect 576118 702448 576124 702460
rect 576176 702448 576182 702500
rect 276014 702380 276020 702432
rect 276072 702420 276078 702432
rect 305730 702420 305736 702432
rect 276072 702392 305736 702420
rect 276072 702380 276078 702392
rect 305730 702380 305736 702392
rect 305788 702380 305794 702432
rect 4338 702312 4344 702364
rect 4396 702352 4402 702364
rect 472710 702352 472716 702364
rect 4396 702324 472716 702352
rect 4396 702312 4402 702324
rect 472710 702312 472716 702324
rect 472768 702312 472774 702364
rect 247402 702244 247408 702296
rect 247460 702284 247466 702296
rect 313274 702284 313280 702296
rect 247460 702256 313280 702284
rect 247460 702244 247466 702256
rect 313274 702244 313280 702256
rect 313332 702244 313338 702296
rect 280982 702176 280988 702228
rect 281040 702216 281046 702228
rect 384298 702216 384304 702228
rect 281040 702188 384304 702216
rect 281040 702176 281046 702188
rect 384298 702176 384304 702188
rect 384356 702176 384362 702228
rect 232682 702108 232688 702160
rect 232740 702148 232746 702160
rect 349798 702148 349804 702160
rect 232740 702120 349804 702148
rect 232740 702108 232746 702120
rect 349798 702108 349804 702120
rect 349856 702108 349862 702160
rect 154022 702040 154028 702092
rect 154080 702080 154086 702092
rect 291838 702080 291844 702092
rect 154080 702052 291844 702080
rect 154080 702040 154086 702052
rect 291838 702040 291844 702052
rect 291896 702040 291902 702092
rect 178586 701972 178592 702024
rect 178644 702012 178650 702024
rect 325602 702012 325608 702024
rect 178644 701984 325608 702012
rect 178644 701972 178650 701984
rect 325602 701972 325608 701984
rect 325660 701972 325666 702024
rect 75454 701904 75460 701956
rect 75512 701944 75518 701956
rect 232866 701944 232872 701956
rect 75512 701916 232872 701944
rect 75512 701904 75518 701916
rect 232866 701904 232872 701916
rect 232924 701904 232930 701956
rect 260834 701904 260840 701956
rect 260892 701944 260898 701956
rect 399018 701944 399024 701956
rect 260892 701916 399024 701944
rect 260892 701904 260898 701916
rect 399018 701904 399024 701916
rect 399076 701904 399082 701956
rect 114278 701836 114284 701888
rect 114336 701876 114342 701888
rect 277486 701876 277492 701888
rect 114336 701848 277492 701876
rect 114336 701836 114342 701848
rect 277486 701836 277492 701848
rect 277544 701836 277550 701888
rect 282914 701836 282920 701888
rect 282972 701876 282978 701888
rect 320450 701876 320456 701888
rect 282972 701848 320456 701876
rect 282972 701836 282978 701848
rect 320450 701836 320456 701848
rect 320508 701836 320514 701888
rect 320910 701836 320916 701888
rect 320968 701876 320974 701888
rect 482554 701876 482560 701888
rect 320968 701848 482560 701876
rect 320968 701836 320974 701848
rect 482554 701836 482560 701848
rect 482612 701836 482618 701888
rect 224954 701768 224960 701820
rect 225012 701808 225018 701820
rect 414198 701808 414204 701820
rect 225012 701780 414204 701808
rect 225012 701768 225018 701780
rect 414198 701768 414204 701780
rect 414256 701768 414262 701820
rect 104802 701700 104808 701752
rect 104860 701740 104866 701752
rect 340874 701740 340880 701752
rect 104860 701712 340880 701740
rect 104860 701700 104866 701712
rect 340874 701700 340880 701712
rect 340932 701700 340938 701752
rect 6638 701632 6644 701684
rect 6696 701672 6702 701684
rect 252278 701672 252284 701684
rect 6696 701644 252284 701672
rect 6696 701632 6702 701644
rect 252278 701632 252284 701644
rect 252336 701632 252342 701684
rect 253198 701632 253204 701684
rect 253256 701672 253262 701684
rect 453022 701672 453028 701684
rect 253256 701644 453028 701672
rect 253256 701632 253262 701644
rect 453022 701632 453028 701644
rect 453080 701632 453086 701684
rect 148962 701564 148968 701616
rect 149020 701604 149026 701616
rect 567838 701604 567844 701616
rect 149020 701576 567844 701604
rect 149020 701564 149026 701576
rect 567838 701564 567844 701576
rect 567896 701564 567902 701616
rect 4246 701496 4252 701548
rect 4304 701536 4310 701548
rect 428458 701536 428464 701548
rect 4304 701508 428464 701536
rect 4304 701496 4310 701508
rect 428458 701496 428464 701508
rect 428516 701496 428522 701548
rect 144270 701428 144276 701480
rect 144328 701468 144334 701480
rect 574922 701468 574928 701480
rect 144328 701440 574928 701468
rect 144328 701428 144334 701440
rect 574922 701428 574928 701440
rect 574980 701428 574986 701480
rect 134426 701360 134432 701412
rect 134484 701400 134490 701412
rect 576210 701400 576216 701412
rect 134484 701372 576216 701400
rect 134484 701360 134490 701372
rect 576210 701360 576216 701372
rect 576268 701360 576274 701412
rect 129458 701292 129464 701344
rect 129516 701332 129522 701344
rect 573450 701332 573456 701344
rect 129516 701304 573456 701332
rect 129516 701292 129522 701304
rect 573450 701292 573456 701304
rect 573508 701292 573514 701344
rect 2406 701224 2412 701276
rect 2464 701264 2470 701276
rect 458174 701264 458180 701276
rect 2464 701236 458180 701264
rect 2464 701224 2470 701236
rect 458174 701224 458180 701236
rect 458232 701224 458238 701276
rect 119706 701156 119712 701208
rect 119764 701196 119770 701208
rect 574830 701196 574836 701208
rect 119764 701168 574836 701196
rect 119764 701156 119770 701168
rect 574830 701156 574836 701168
rect 574888 701156 574894 701208
rect 566 701088 572 701140
rect 624 701128 630 701140
rect 467834 701128 467840 701140
rect 624 701100 467840 701128
rect 624 701088 630 701100
rect 467834 701088 467840 701100
rect 467892 701088 467898 701140
rect 335354 701060 335360 701072
rect 313292 701032 335360 701060
rect 72970 700952 72976 701004
rect 73028 700992 73034 701004
rect 313292 700992 313320 701032
rect 335354 701020 335360 701032
rect 335412 701020 335418 701072
rect 340966 701020 340972 701072
rect 341024 701060 341030 701072
rect 511994 701060 512000 701072
rect 341024 701032 512000 701060
rect 341024 701020 341030 701032
rect 511994 701020 512000 701032
rect 512052 701020 512058 701072
rect 556890 701020 556896 701072
rect 556948 701060 556954 701072
rect 564434 701060 564440 701072
rect 556948 701032 564440 701060
rect 556948 701020 556954 701032
rect 564434 701020 564440 701032
rect 564492 701020 564498 701072
rect 73028 700964 313320 700992
rect 316006 700964 321554 700992
rect 73028 700952 73034 700964
rect 137830 700884 137836 700936
rect 137888 700924 137894 700936
rect 282914 700924 282920 700936
rect 137888 700896 282920 700924
rect 137888 700884 137894 700896
rect 282914 700884 282920 700896
rect 282972 700884 282978 700936
rect 284110 700884 284116 700936
rect 284168 700924 284174 700936
rect 295886 700924 295892 700936
rect 284168 700896 295892 700924
rect 284168 700884 284174 700896
rect 295886 700884 295892 700896
rect 295944 700884 295950 700936
rect 298002 700884 298008 700936
rect 298060 700924 298066 700936
rect 300118 700924 300124 700936
rect 298060 700896 300124 700924
rect 298060 700884 298066 700896
rect 300118 700884 300124 700896
rect 300176 700884 300182 700936
rect 313274 700884 313280 700936
rect 313332 700924 313338 700936
rect 316006 700924 316034 700964
rect 313332 700896 316034 700924
rect 321526 700924 321554 700964
rect 462314 700924 462320 700936
rect 321526 700896 462320 700924
rect 313332 700884 313338 700896
rect 462314 700884 462320 700896
rect 462372 700884 462378 700936
rect 503898 700884 503904 700936
rect 503956 700924 503962 700936
rect 559650 700924 559656 700936
rect 503956 700896 559656 700924
rect 503956 700884 503962 700896
rect 559650 700884 559656 700896
rect 559708 700884 559714 700936
rect 154114 700816 154120 700868
rect 154172 700856 154178 700868
rect 325326 700856 325332 700868
rect 154172 700828 325332 700856
rect 154172 700816 154178 700828
rect 325326 700816 325332 700828
rect 325384 700816 325390 700868
rect 325602 700816 325608 700868
rect 325660 700856 325666 700868
rect 580718 700856 580724 700868
rect 325660 700828 580724 700856
rect 325660 700816 325666 700828
rect 580718 700816 580724 700828
rect 580776 700816 580782 700868
rect 3786 700748 3792 700800
rect 3844 700788 3850 700800
rect 207014 700788 207020 700800
rect 3844 700760 207020 700788
rect 3844 700748 3850 700760
rect 207014 700748 207020 700760
rect 207072 700748 207078 700800
rect 252278 700748 252284 700800
rect 252336 700788 252342 700800
rect 478506 700788 478512 700800
rect 252336 700760 478512 700788
rect 252336 700748 252342 700760
rect 478506 700748 478512 700760
rect 478564 700748 478570 700800
rect 3326 700680 3332 700732
rect 3384 700720 3390 700732
rect 253198 700720 253204 700732
rect 3384 700692 253204 700720
rect 3384 700680 3390 700692
rect 253198 700680 253204 700692
rect 253256 700680 253262 700732
rect 266998 700680 267004 700732
rect 267056 700720 267062 700732
rect 413646 700720 413652 700732
rect 267056 700692 413652 700720
rect 267056 700680 267062 700692
rect 413646 700680 413652 700692
rect 413704 700680 413710 700732
rect 89162 700612 89168 700664
rect 89220 700652 89226 700664
rect 340046 700652 340052 700664
rect 89220 700624 340052 700652
rect 89220 700612 89226 700624
rect 340046 700612 340052 700624
rect 340104 700612 340110 700664
rect 340874 700612 340880 700664
rect 340932 700652 340938 700664
rect 580442 700652 580448 700664
rect 340932 700624 580448 700652
rect 340932 700612 340938 700624
rect 580442 700612 580448 700624
rect 580500 700612 580506 700664
rect 3142 700544 3148 700596
rect 3200 700584 3206 700596
rect 260834 700584 260840 700596
rect 3200 700556 260840 700584
rect 3200 700544 3206 700556
rect 260834 700544 260840 700556
rect 260892 700544 260898 700596
rect 267642 700544 267648 700596
rect 267700 700584 267706 700596
rect 269209 700587 269267 700593
rect 269209 700584 269221 700587
rect 267700 700556 269221 700584
rect 267700 700544 267706 700556
rect 269209 700553 269221 700556
rect 269255 700553 269267 700587
rect 280982 700584 280988 700596
rect 269209 700547 269267 700553
rect 269316 700556 280988 700584
rect 2958 700476 2964 700528
rect 3016 700516 3022 700528
rect 269316 700516 269344 700556
rect 280982 700544 280988 700556
rect 281040 700544 281046 700596
rect 281353 700587 281411 700593
rect 281353 700553 281365 700587
rect 281399 700584 281411 700587
rect 332502 700584 332508 700596
rect 281399 700556 332508 700584
rect 281399 700553 281411 700556
rect 281353 700547 281411 700553
rect 332502 700544 332508 700556
rect 332560 700544 332566 700596
rect 349798 700544 349804 700596
rect 349856 700584 349862 700596
rect 527174 700584 527180 700596
rect 349856 700556 527180 700584
rect 349856 700544 349862 700556
rect 527174 700544 527180 700556
rect 527232 700544 527238 700596
rect 3016 700488 269344 700516
rect 269393 700519 269451 700525
rect 3016 700476 3022 700488
rect 269393 700485 269405 700519
rect 269439 700516 269451 700519
rect 291378 700516 291384 700528
rect 269439 700488 291384 700516
rect 269439 700485 269451 700488
rect 269393 700479 269451 700485
rect 291378 700476 291384 700488
rect 291436 700476 291442 700528
rect 291838 700476 291844 700528
rect 291896 700516 291902 700528
rect 580626 700516 580632 700528
rect 291896 700488 580632 700516
rect 291896 700476 291902 700488
rect 580626 700476 580632 700488
rect 580684 700476 580690 700528
rect 4062 700408 4068 700460
rect 4120 700448 4126 700460
rect 224954 700448 224960 700460
rect 4120 700420 224960 700448
rect 4120 700408 4126 700420
rect 224954 700408 224960 700420
rect 225012 700408 225018 700460
rect 237098 700408 237104 700460
rect 237156 700448 237162 700460
rect 543458 700448 543464 700460
rect 237156 700420 543464 700448
rect 237156 700408 237162 700420
rect 543458 700408 543464 700420
rect 543516 700408 543522 700460
rect 24302 700340 24308 700392
rect 24360 700380 24366 700392
rect 354950 700380 354956 700392
rect 24360 700352 354956 700380
rect 24360 700340 24366 700352
rect 354950 700340 354956 700352
rect 355008 700340 355014 700392
rect 8110 700272 8116 700324
rect 8168 700312 8174 700324
rect 349890 700312 349896 700324
rect 8168 700284 349896 700312
rect 8168 700272 8174 700284
rect 349890 700272 349896 700284
rect 349948 700272 349954 700324
rect 262122 700204 262128 700256
rect 262180 700244 262186 700256
rect 397454 700244 397460 700256
rect 262180 700216 397460 700244
rect 262180 700204 262186 700216
rect 397454 700204 397460 700216
rect 397512 700204 397518 700256
rect 218974 700136 218980 700188
rect 219032 700176 219038 700188
rect 310928 700176 310934 700188
rect 219032 700148 310934 700176
rect 219032 700136 219038 700148
rect 310928 700136 310934 700148
rect 310986 700136 310992 700188
rect 202782 700068 202788 700120
rect 202840 700108 202846 700120
rect 276014 700108 276020 700120
rect 202840 700080 276020 700108
rect 202840 700068 202846 700080
rect 276014 700068 276020 700080
rect 276072 700068 276078 700120
rect 276520 700068 276526 700120
rect 276578 700108 276584 700120
rect 281353 700111 281411 700117
rect 281353 700108 281365 700111
rect 276578 700080 281365 700108
rect 276578 700068 276584 700080
rect 281353 700077 281365 700080
rect 281399 700077 281411 700111
rect 281353 700071 281411 700077
rect 281488 700068 281494 700120
rect 281546 700108 281552 700120
rect 348786 700108 348792 700120
rect 281546 700080 348792 700108
rect 281546 700068 281552 700080
rect 348786 700068 348792 700080
rect 348844 700068 348850 700120
rect 217870 700000 217876 700052
rect 217928 700040 217934 700052
rect 563514 700040 563520 700052
rect 217928 700012 563520 700040
rect 217928 700000 217934 700012
rect 563514 700000 563520 700012
rect 563572 700000 563578 700052
rect 222838 699932 222844 699984
rect 222896 699972 222902 699984
rect 579062 699972 579068 699984
rect 222896 699944 579068 699972
rect 222896 699932 222902 699944
rect 579062 699932 579068 699944
rect 579120 699932 579126 699984
rect 1026 699864 1032 699916
rect 1084 699904 1090 699916
rect 364610 699904 364616 699916
rect 1084 699876 364616 699904
rect 1084 699864 1090 699876
rect 364610 699864 364616 699876
rect 364668 699864 364674 699916
rect 208118 699796 208124 699848
rect 208176 699836 208182 699848
rect 570874 699836 570880 699848
rect 208176 699808 570880 699836
rect 208176 699796 208182 699808
rect 570874 699796 570880 699808
rect 570932 699796 570938 699848
rect 3050 699728 3056 699780
rect 3108 699768 3114 699780
rect 369762 699768 369768 699780
rect 3108 699740 369768 699768
rect 3108 699728 3114 699740
rect 369762 699728 369768 699740
rect 369820 699728 369826 699780
rect 193214 699660 193220 699712
rect 193272 699700 193278 699712
rect 578970 699700 578976 699712
rect 193272 699672 578976 699700
rect 193272 699660 193278 699672
rect 578970 699660 578976 699672
rect 579028 699660 579034 699712
rect 277486 699592 277492 699644
rect 277544 699632 277550 699644
rect 580534 699632 580540 699644
rect 277544 699604 580540 699632
rect 277544 699592 277550 699604
rect 580534 699592 580540 699604
rect 580592 699592 580598 699644
rect 3970 699524 3976 699576
rect 4028 699564 4034 699576
rect 320910 699564 320916 699576
rect 4028 699536 320916 699564
rect 4028 699524 4034 699536
rect 320910 699524 320916 699536
rect 320968 699524 320974 699576
rect 3694 699456 3700 699508
rect 3752 699496 3758 699508
rect 340966 699496 340972 699508
rect 3752 699468 340972 699496
rect 3752 699456 3758 699468
rect 340966 699456 340972 699468
rect 341024 699456 341030 699508
rect 379514 699496 379520 699508
rect 379475 699468 379520 699496
rect 379514 699456 379520 699468
rect 379572 699456 379578 699508
rect 386230 699496 386236 699508
rect 386191 699468 386236 699496
rect 386230 699456 386236 699468
rect 386288 699456 386294 699508
rect 394142 699496 394148 699508
rect 394103 699468 394148 699496
rect 394142 699456 394148 699468
rect 394200 699456 394206 699508
rect 408862 699496 408868 699508
rect 408823 699468 408868 699496
rect 408862 699456 408868 699468
rect 408920 699456 408926 699508
rect 423674 699496 423680 699508
rect 423635 699468 423680 699496
rect 423674 699456 423680 699468
rect 423732 699456 423738 699508
rect 438302 699496 438308 699508
rect 438263 699468 438308 699496
rect 438302 699456 438308 699468
rect 438360 699456 438366 699508
rect 521838 699496 521844 699508
rect 521799 699468 521844 699496
rect 521838 699456 521844 699468
rect 521896 699456 521902 699508
rect 232866 699388 232872 699440
rect 232924 699428 232930 699440
rect 580350 699428 580356 699440
rect 232924 699400 580356 699428
rect 232924 699388 232930 699400
rect 580350 699388 580356 699400
rect 580408 699388 580414 699440
rect 35986 699360 35992 699372
rect 35947 699332 35992 699360
rect 35986 699320 35992 699332
rect 36044 699320 36050 699372
rect 65610 699360 65616 699372
rect 65571 699332 65616 699360
rect 65610 699320 65616 699332
rect 65668 699320 65674 699372
rect 70394 699360 70400 699372
rect 70355 699332 70400 699360
rect 70394 699320 70400 699332
rect 70452 699320 70458 699372
rect 80146 699360 80152 699372
rect 80107 699332 80152 699360
rect 80146 699320 80152 699332
rect 80204 699320 80210 699372
rect 85298 699360 85304 699372
rect 85259 699332 85304 699360
rect 85298 699320 85304 699332
rect 85356 699320 85362 699372
rect 100018 699360 100024 699372
rect 99979 699332 100024 699360
rect 100018 699320 100024 699332
rect 100076 699320 100082 699372
rect 109862 699360 109868 699372
rect 109823 699332 109868 699360
rect 109862 699320 109868 699332
rect 109920 699320 109926 699372
rect 158806 699360 158812 699372
rect 158767 699332 158812 699360
rect 158806 699320 158812 699332
rect 158864 699320 158870 699372
rect 168834 699360 168840 699372
rect 168795 699332 168840 699360
rect 168834 699320 168840 699332
rect 168892 699320 168898 699372
rect 173710 699360 173716 699372
rect 173671 699332 173716 699360
rect 173710 699320 173716 699332
rect 173768 699320 173774 699372
rect 188430 699360 188436 699372
rect 188391 699332 188436 699360
rect 188430 699320 188436 699332
rect 188488 699320 188494 699372
rect 202966 699320 202972 699372
rect 203024 699360 203030 699372
rect 573726 699360 573732 699372
rect 203024 699332 573732 699360
rect 203024 699320 203030 699332
rect 573726 699320 573732 699332
rect 573784 699320 573790 699372
rect 934 699252 940 699304
rect 992 699292 998 699304
rect 379517 699295 379575 699301
rect 379517 699292 379529 699295
rect 992 699264 379529 699292
rect 992 699252 998 699264
rect 379517 699261 379529 699264
rect 379563 699261 379575 699295
rect 379517 699255 379575 699261
rect 188433 699227 188491 699233
rect 188433 699193 188445 699227
rect 188479 699224 188491 699227
rect 569586 699224 569592 699236
rect 188479 699196 569592 699224
rect 188479 699193 188491 699196
rect 188433 699187 188491 699193
rect 569586 699184 569592 699196
rect 569644 699184 569650 699236
rect 842 699116 848 699168
rect 900 699156 906 699168
rect 394145 699159 394203 699165
rect 394145 699156 394157 699159
rect 900 699128 394157 699156
rect 900 699116 906 699128
rect 394145 699125 394157 699128
rect 394191 699125 394203 699159
rect 394145 699119 394203 699125
rect 168837 699091 168895 699097
rect 168837 699057 168849 699091
rect 168883 699088 168895 699091
rect 565354 699088 565360 699100
rect 168883 699060 565360 699088
rect 168883 699057 168895 699060
rect 168837 699051 168895 699057
rect 565354 699048 565360 699060
rect 565412 699048 565418 699100
rect 173713 699023 173771 699029
rect 173713 698989 173725 699023
rect 173759 699020 173771 699023
rect 573542 699020 573548 699032
rect 173759 698992 573548 699020
rect 173759 698989 173771 698992
rect 173713 698983 173771 698989
rect 573542 698980 573548 698992
rect 573600 698980 573606 699032
rect 750 698912 756 698964
rect 808 698952 814 698964
rect 408865 698955 408923 698961
rect 408865 698952 408877 698955
rect 808 698924 408877 698952
rect 808 698912 814 698924
rect 408865 698921 408877 698924
rect 408911 698921 408923 698955
rect 408865 698915 408923 698921
rect 158809 698887 158867 698893
rect 158809 698853 158821 698887
rect 158855 698884 158867 698887
rect 578878 698884 578884 698896
rect 158855 698856 578884 698884
rect 158855 698853 158867 698856
rect 158809 698847 158867 698853
rect 578878 698844 578884 698856
rect 578936 698844 578942 698896
rect 658 698776 664 698828
rect 716 698816 722 698828
rect 423677 698819 423735 698825
rect 423677 698816 423689 698819
rect 716 698788 423689 698816
rect 716 698776 722 698788
rect 423677 698785 423689 698788
rect 423723 698785 423735 698819
rect 423677 698779 423735 698785
rect 2590 698708 2596 698760
rect 2648 698748 2654 698760
rect 438305 698751 438363 698757
rect 438305 698748 438317 698751
rect 2648 698720 438317 698748
rect 2648 698708 2654 698720
rect 438305 698717 438317 698720
rect 438351 698717 438363 698751
rect 438305 698711 438363 698717
rect 109865 698683 109923 698689
rect 109865 698649 109877 698683
rect 109911 698680 109923 698683
rect 569494 698680 569500 698692
rect 109911 698652 569500 698680
rect 109911 698649 109923 698652
rect 109865 698643 109923 698649
rect 569494 698640 569500 698652
rect 569552 698640 569558 698692
rect 100021 698615 100079 698621
rect 100021 698581 100033 698615
rect 100067 698612 100079 698615
rect 572070 698612 572076 698624
rect 100067 698584 572076 698612
rect 100067 698581 100079 698584
rect 100021 698575 100079 698581
rect 572070 698572 572076 698584
rect 572128 698572 572134 698624
rect 85301 698547 85359 698553
rect 85301 698513 85313 698547
rect 85347 698544 85359 698547
rect 571978 698544 571984 698556
rect 85347 698516 571984 698544
rect 85347 698513 85359 698516
rect 85301 698507 85359 698513
rect 571978 698504 571984 698516
rect 572036 698504 572042 698556
rect 80149 698479 80207 698485
rect 80149 698445 80161 698479
rect 80195 698476 80207 698479
rect 566734 698476 566740 698488
rect 80195 698448 566740 698476
rect 80195 698445 80207 698448
rect 80149 698439 80207 698445
rect 566734 698436 566740 698448
rect 566792 698436 566798 698488
rect 70397 698411 70455 698417
rect 70397 698377 70409 698411
rect 70443 698408 70455 698411
rect 569402 698408 569408 698420
rect 70443 698380 569408 698408
rect 70443 698377 70455 698380
rect 70397 698371 70455 698377
rect 569402 698368 569408 698380
rect 569460 698368 569466 698420
rect 65613 698343 65671 698349
rect 65613 698309 65625 698343
rect 65659 698340 65671 698343
rect 566550 698340 566556 698352
rect 65659 698312 566556 698340
rect 65659 698309 65671 698312
rect 65613 698303 65671 698309
rect 566550 698300 566556 698312
rect 566608 698300 566614 698352
rect 563514 698232 563520 698284
rect 563572 698272 563578 698284
rect 580166 698272 580172 698284
rect 563572 698244 580172 698272
rect 563572 698232 563578 698244
rect 580166 698232 580172 698244
rect 580224 698232 580230 698284
rect 367097 697867 367155 697873
rect 367097 697833 367109 697867
rect 367143 697864 367155 697867
rect 367143 697836 376754 697864
rect 367143 697833 367155 697836
rect 367097 697827 367155 697833
rect 371881 697799 371939 697805
rect 371881 697796 371893 697799
rect 367204 697768 371893 697796
rect 367204 697728 367232 697768
rect 371881 697765 371893 697768
rect 371927 697765 371939 697799
rect 371881 697759 371939 697765
rect 367066 697700 367232 697728
rect 376726 697728 376754 697836
rect 386233 697731 386291 697737
rect 386233 697728 386245 697731
rect 376726 697700 386245 697728
rect 198 697620 204 697672
rect 256 697660 262 697672
rect 367066 697660 367094 697700
rect 386233 697697 386245 697700
rect 386279 697697 386291 697731
rect 386233 697691 386291 697697
rect 256 697632 367094 697660
rect 371881 697663 371939 697669
rect 256 697620 262 697632
rect 371881 697629 371893 697663
rect 371927 697660 371939 697663
rect 521841 697663 521899 697669
rect 521841 697660 521853 697663
rect 371927 697632 521853 697660
rect 371927 697629 371939 697632
rect 371881 697623 371939 697629
rect 521841 697629 521853 697632
rect 521887 697629 521899 697663
rect 521841 697623 521899 697629
rect 35989 697595 36047 697601
rect 35989 697561 36001 697595
rect 36035 697592 36047 697595
rect 367189 697595 367247 697601
rect 367189 697592 367201 697595
rect 36035 697564 367201 697592
rect 36035 697561 36047 697564
rect 35989 697555 36047 697561
rect 367189 697561 367201 697564
rect 367235 697561 367247 697595
rect 367189 697555 367247 697561
rect 367281 697595 367339 697601
rect 367281 697561 367293 697595
rect 367327 697561 367339 697595
rect 574738 697592 574744 697604
rect 367281 697555 367339 697561
rect 376726 697564 574744 697592
rect 3418 697484 3424 697536
rect 3476 697524 3482 697536
rect 367097 697527 367155 697533
rect 367097 697524 367109 697527
rect 3476 697496 367109 697524
rect 3476 697484 3482 697496
rect 367097 697493 367109 697496
rect 367143 697493 367155 697527
rect 367296 697524 367324 697555
rect 376726 697524 376754 697564
rect 574738 697552 574744 697564
rect 574796 697552 574802 697604
rect 367296 697496 376754 697524
rect 367097 697487 367155 697493
rect 576394 671984 576400 672036
rect 576452 672024 576458 672036
rect 579614 672024 579620 672036
rect 576452 671996 579620 672024
rect 576452 671984 576458 671996
rect 579614 671984 579620 671996
rect 579672 671984 579678 672036
rect 573726 644376 573732 644428
rect 573784 644416 573790 644428
rect 580166 644416 580172 644428
rect 573784 644388 580172 644416
rect 573784 644376 573790 644388
rect 580166 644376 580172 644388
rect 580224 644376 580230 644428
rect 570874 632000 570880 632052
rect 570932 632040 570938 632052
rect 580166 632040 580172 632052
rect 570932 632012 580172 632040
rect 570932 632000 570938 632012
rect 580166 632000 580172 632012
rect 580224 632000 580230 632052
rect 3050 619080 3056 619132
rect 3108 619120 3114 619132
rect 4246 619120 4252 619132
rect 3108 619092 4252 619120
rect 3108 619080 3114 619092
rect 4246 619080 4252 619092
rect 4304 619080 4310 619132
rect 575014 618196 575020 618248
rect 575072 618236 575078 618248
rect 580166 618236 580172 618248
rect 575072 618208 580172 618236
rect 575072 618196 575078 618208
rect 580166 618196 580172 618208
rect 580224 618196 580230 618248
rect 569586 591948 569592 592000
rect 569644 591988 569650 592000
rect 580166 591988 580172 592000
rect 569644 591960 580172 591988
rect 569644 591948 569650 591960
rect 580166 591948 580172 591960
rect 580224 591948 580230 592000
rect 573634 564340 573640 564392
rect 573692 564380 573698 564392
rect 580166 564380 580172 564392
rect 573692 564352 580172 564380
rect 573692 564340 573698 564352
rect 580166 564340 580172 564352
rect 580224 564340 580230 564392
rect 573542 538160 573548 538212
rect 573600 538200 573606 538212
rect 580166 538200 580172 538212
rect 573600 538172 580172 538200
rect 573600 538160 573606 538172
rect 580166 538160 580172 538172
rect 580224 538160 580230 538212
rect 3142 514768 3148 514820
rect 3200 514808 3206 514820
rect 4338 514808 4344 514820
rect 3200 514780 4344 514808
rect 3200 514768 3206 514780
rect 4338 514768 4344 514780
rect 4396 514768 4402 514820
rect 565354 511912 565360 511964
rect 565412 511952 565418 511964
rect 580166 511952 580172 511964
rect 565412 511924 580172 511952
rect 565412 511912 565418 511924
rect 580166 511912 580172 511924
rect 580224 511912 580230 511964
rect 576302 471928 576308 471980
rect 576360 471968 576366 471980
rect 579798 471968 579804 471980
rect 576360 471940 579804 471968
rect 576360 471928 576366 471940
rect 579798 471928 579804 471940
rect 579856 471928 579862 471980
rect 574922 431876 574928 431928
rect 574980 431916 574986 431928
rect 579706 431916 579712 431928
rect 574980 431888 579712 431916
rect 574980 431876 574986 431888
rect 579706 431876 579712 431888
rect 579764 431876 579770 431928
rect 567838 419432 567844 419484
rect 567896 419472 567902 419484
rect 580166 419472 580172 419484
rect 567896 419444 580172 419472
rect 567896 419432 567902 419444
rect 580166 419432 580172 419444
rect 580224 419432 580230 419484
rect 572162 405628 572168 405680
rect 572220 405668 572226 405680
rect 580166 405668 580172 405680
rect 572220 405640 580172 405668
rect 572220 405628 572226 405640
rect 580166 405628 580172 405640
rect 580224 405628 580230 405680
rect 573450 379448 573456 379500
rect 573508 379488 573514 379500
rect 579614 379488 579620 379500
rect 573508 379460 579620 379488
rect 573508 379448 573514 379460
rect 579614 379448 579620 379460
rect 579672 379448 579678 379500
rect 576210 365644 576216 365696
rect 576268 365684 576274 365696
rect 580166 365684 580172 365696
rect 576268 365656 580172 365684
rect 576268 365644 576274 365656
rect 580166 365644 580172 365656
rect 580224 365644 580230 365696
rect 570782 353200 570788 353252
rect 570840 353240 570846 353252
rect 580166 353240 580172 353252
rect 570840 353212 580172 353240
rect 570840 353200 570846 353212
rect 580166 353200 580172 353212
rect 580224 353200 580230 353252
rect 574830 313216 574836 313268
rect 574888 313256 574894 313268
rect 579706 313256 579712 313268
rect 574888 313228 579712 313256
rect 574888 313216 574894 313228
rect 579706 313216 579712 313228
rect 579764 313216 579770 313268
rect 569494 299412 569500 299464
rect 569552 299452 569558 299464
rect 579798 299452 579804 299464
rect 569552 299424 579804 299452
rect 569552 299412 569558 299424
rect 579798 299412 579804 299424
rect 579856 299412 579862 299464
rect 572070 273164 572076 273216
rect 572128 273204 572134 273216
rect 580166 273204 580172 273216
rect 572128 273176 580172 273204
rect 572128 273164 572134 273176
rect 580166 273164 580172 273176
rect 580224 273164 580230 273216
rect 565262 245556 565268 245608
rect 565320 245596 565326 245608
rect 580166 245596 580172 245608
rect 565320 245568 580172 245596
rect 565320 245556 565326 245568
rect 580166 245556 580172 245568
rect 580224 245556 580230 245608
rect 571978 233180 571984 233232
rect 572036 233220 572042 233232
rect 580166 233220 580172 233232
rect 572036 233192 580172 233220
rect 572036 233180 572042 233192
rect 580166 233180 580172 233192
rect 580224 233180 580230 233232
rect 573358 219376 573364 219428
rect 573416 219416 573422 219428
rect 580166 219416 580172 219428
rect 573416 219388 580172 219416
rect 573416 219376 573422 219388
rect 580166 219376 580172 219388
rect 580224 219376 580230 219428
rect 566734 206932 566740 206984
rect 566792 206972 566798 206984
rect 579890 206972 579896 206984
rect 566792 206944 579896 206972
rect 566792 206932 566798 206944
rect 579890 206932 579896 206944
rect 579948 206932 579954 206984
rect 569402 193128 569408 193180
rect 569460 193168 569466 193180
rect 580166 193168 580172 193180
rect 569460 193140 580172 193168
rect 569460 193128 569466 193140
rect 580166 193128 580172 193140
rect 580224 193128 580230 193180
rect 566550 166948 566556 167000
rect 566608 166988 566614 167000
rect 580166 166988 580172 167000
rect 566608 166960 580172 166988
rect 566608 166948 566614 166960
rect 580166 166948 580172 166960
rect 580224 166948 580230 167000
rect 569310 153144 569316 153196
rect 569368 153184 569374 153196
rect 579798 153184 579804 153196
rect 569368 153156 579804 153184
rect 569368 153144 569374 153156
rect 579798 153144 579804 153156
rect 579856 153144 579862 153196
rect 570690 139340 570696 139392
rect 570748 139380 570754 139392
rect 580166 139380 580172 139392
rect 570748 139352 580172 139380
rect 570748 139340 570754 139352
rect 580166 139340 580172 139352
rect 580224 139340 580230 139392
rect 565170 126896 565176 126948
rect 565228 126936 565234 126948
rect 580166 126936 580172 126948
rect 565228 126908 580172 126936
rect 565228 126896 565234 126908
rect 580166 126896 580172 126908
rect 580224 126896 580230 126948
rect 566642 113092 566648 113144
rect 566700 113132 566706 113144
rect 580166 113132 580172 113144
rect 566700 113104 580172 113132
rect 566700 113092 566706 113104
rect 580166 113092 580172 113104
rect 580224 113092 580230 113144
rect 570598 100648 570604 100700
rect 570656 100688 570662 100700
rect 580166 100688 580172 100700
rect 570656 100660 580172 100688
rect 570656 100648 570662 100660
rect 580166 100648 580172 100660
rect 580224 100648 580230 100700
rect 574738 86912 574744 86964
rect 574796 86952 574802 86964
rect 580166 86952 580172 86964
rect 574796 86924 580172 86952
rect 574796 86912 574802 86924
rect 580166 86912 580172 86924
rect 580224 86912 580230 86964
rect 565078 73108 565084 73160
rect 565136 73148 565142 73160
rect 579982 73148 579988 73160
rect 565136 73120 579988 73148
rect 565136 73108 565142 73120
rect 579982 73108 579988 73120
rect 580040 73108 580046 73160
rect 569218 60664 569224 60716
rect 569276 60704 569282 60716
rect 580166 60704 580172 60716
rect 569276 60676 580172 60704
rect 569276 60664 569282 60676
rect 580166 60664 580172 60676
rect 580224 60664 580230 60716
rect 576118 46860 576124 46912
rect 576176 46900 576182 46912
rect 580166 46900 580172 46912
rect 576176 46872 580172 46900
rect 576176 46860 576182 46872
rect 580166 46860 580172 46872
rect 580224 46860 580230 46912
rect 566458 33056 566464 33108
rect 566516 33096 566522 33108
rect 580166 33096 580172 33108
rect 566516 33068 580172 33096
rect 566516 33056 566522 33068
rect 580166 33056 580172 33068
rect 580224 33056 580230 33108
rect 577498 20612 577504 20664
rect 577556 20652 577562 20664
rect 579706 20652 579712 20664
rect 577556 20624 579712 20652
rect 577556 20612 577562 20624
rect 579706 20612 579712 20624
rect 579764 20612 579770 20664
rect 569862 3068 569868 3120
rect 569920 3108 569926 3120
rect 577406 3108 577412 3120
rect 569920 3080 577412 3108
rect 569920 3068 569926 3080
rect 577406 3068 577412 3080
rect 577464 3068 577470 3120
rect 563698 3000 563704 3052
rect 563756 3040 563762 3052
rect 583386 3040 583392 3052
rect 563756 3012 583392 3040
rect 563756 3000 563762 3012
rect 583386 3000 583392 3012
rect 583444 3000 583450 3052
rect 563514 2932 563520 2984
rect 563572 2972 563578 2984
rect 573910 2972 573916 2984
rect 563572 2944 573916 2972
rect 563572 2932 563578 2944
rect 573910 2932 573916 2944
rect 573968 2932 573974 2984
rect 563606 2864 563612 2916
rect 563664 2904 563670 2916
rect 563664 2876 567194 2904
rect 563664 2864 563670 2876
rect 567166 2836 567194 2876
rect 575474 2864 575480 2916
rect 575532 2904 575538 2916
rect 582190 2904 582196 2916
rect 575532 2876 582196 2904
rect 575532 2864 575538 2876
rect 582190 2864 582196 2876
rect 582248 2864 582254 2916
rect 576302 2836 576308 2848
rect 567166 2808 576308 2836
rect 576302 2796 576308 2808
rect 576360 2796 576366 2848
rect 2958 2048 2964 2100
rect 3016 2088 3022 2100
rect 564434 2088 564440 2100
rect 3016 2060 564440 2088
rect 3016 2048 3022 2060
rect 564434 2048 564440 2060
rect 564492 2048 564498 2100
rect 565906 1368 565912 1420
rect 565964 1408 565970 1420
rect 569126 1408 569132 1420
rect 565964 1380 569132 1408
rect 565964 1368 565970 1380
rect 569126 1368 569132 1380
rect 569184 1368 569190 1420
rect 413741 1343 413799 1349
rect 413741 1309 413753 1343
rect 413787 1340 413799 1343
rect 426345 1343 426403 1349
rect 426345 1340 426357 1343
rect 413787 1312 426357 1340
rect 413787 1309 413799 1312
rect 413741 1303 413799 1309
rect 426345 1309 426357 1312
rect 426391 1309 426403 1343
rect 426345 1303 426403 1309
rect 494425 1275 494483 1281
rect 494425 1241 494437 1275
rect 494471 1272 494483 1275
rect 510249 1275 510307 1281
rect 510249 1272 510261 1275
rect 494471 1244 510261 1272
rect 494471 1241 494483 1244
rect 494425 1235 494483 1241
rect 510249 1241 510261 1244
rect 510295 1241 510307 1275
rect 510249 1235 510307 1241
rect 460201 1207 460259 1213
rect 460201 1173 460213 1207
rect 460247 1204 460259 1207
rect 474553 1207 474611 1213
rect 474553 1204 474565 1207
rect 460247 1176 474565 1204
rect 460247 1173 460259 1176
rect 460201 1167 460259 1173
rect 474553 1173 474565 1176
rect 474599 1173 474611 1207
rect 474553 1167 474611 1173
rect 495345 1207 495403 1213
rect 495345 1173 495357 1207
rect 495391 1204 495403 1207
rect 511261 1207 511319 1213
rect 511261 1204 511273 1207
rect 495391 1176 511273 1204
rect 495391 1173 495403 1176
rect 495345 1167 495403 1173
rect 511261 1173 511273 1176
rect 511307 1173 511319 1207
rect 511261 1167 511319 1173
rect 562229 1207 562287 1213
rect 562229 1173 562241 1207
rect 562275 1204 562287 1207
rect 566826 1204 566832 1216
rect 562275 1176 566832 1204
rect 562275 1173 562287 1176
rect 562229 1167 562287 1173
rect 566826 1164 566832 1176
rect 566884 1164 566890 1216
rect 457993 1139 458051 1145
rect 457993 1105 458005 1139
rect 458039 1136 458051 1139
rect 472253 1139 472311 1145
rect 472253 1136 472265 1139
rect 458039 1108 472265 1136
rect 458039 1105 458051 1108
rect 457993 1099 458051 1105
rect 472253 1105 472265 1108
rect 472299 1105 472311 1139
rect 472253 1099 472311 1105
rect 476209 1139 476267 1145
rect 476209 1105 476221 1139
rect 476255 1136 476267 1139
rect 491113 1139 491171 1145
rect 491113 1136 491125 1139
rect 476255 1108 491125 1136
rect 476255 1105 476267 1108
rect 476209 1099 476267 1105
rect 491113 1105 491125 1108
rect 491159 1105 491171 1139
rect 491113 1099 491171 1105
rect 496725 1139 496783 1145
rect 496725 1105 496737 1139
rect 496771 1136 496783 1139
rect 512457 1139 512515 1145
rect 512457 1136 512469 1139
rect 496771 1108 512469 1136
rect 496771 1105 496783 1108
rect 496725 1099 496783 1105
rect 512457 1105 512469 1108
rect 512503 1105 512515 1139
rect 512457 1099 512515 1105
rect 519357 1139 519415 1145
rect 519357 1105 519369 1139
rect 519403 1136 519415 1139
rect 535825 1139 535883 1145
rect 535825 1136 535837 1139
rect 519403 1108 535837 1136
rect 519403 1105 519415 1108
rect 519357 1099 519415 1105
rect 535825 1105 535837 1108
rect 535871 1105 535883 1139
rect 535825 1099 535883 1105
rect 557997 1139 558055 1145
rect 557997 1105 558009 1139
rect 558043 1136 558055 1139
rect 563606 1136 563612 1148
rect 558043 1108 563612 1136
rect 558043 1105 558055 1108
rect 557997 1099 558055 1105
rect 563606 1096 563612 1108
rect 563664 1096 563670 1148
rect 417145 1071 417203 1077
rect 417145 1037 417157 1071
rect 417191 1068 417203 1071
rect 429013 1071 429071 1077
rect 429013 1068 429025 1071
rect 417191 1040 429025 1068
rect 417191 1037 417203 1040
rect 417145 1031 417203 1037
rect 429013 1037 429025 1040
rect 429059 1037 429071 1071
rect 429013 1031 429071 1037
rect 442169 1071 442227 1077
rect 442169 1037 442181 1071
rect 442215 1068 442227 1071
rect 455325 1071 455383 1077
rect 455325 1068 455337 1071
rect 442215 1040 455337 1068
rect 442215 1037 442227 1040
rect 442169 1031 442227 1037
rect 455325 1037 455337 1040
rect 455371 1037 455383 1071
rect 455325 1031 455383 1037
rect 456521 1071 456579 1077
rect 456521 1037 456533 1071
rect 456567 1068 456579 1071
rect 472805 1071 472863 1077
rect 456567 1040 465764 1068
rect 456567 1037 456579 1040
rect 456521 1031 456579 1037
rect 430393 1003 430451 1009
rect 430393 969 430405 1003
rect 430439 1000 430451 1003
rect 443825 1003 443883 1009
rect 443825 1000 443837 1003
rect 430439 972 443837 1000
rect 430439 969 430451 972
rect 430393 963 430451 969
rect 443825 969 443837 972
rect 443871 969 443883 1003
rect 443825 963 443883 969
rect 448977 1003 449035 1009
rect 448977 969 448989 1003
rect 449023 1000 449035 1003
rect 462225 1003 462283 1009
rect 462225 1000 462237 1003
rect 449023 972 462237 1000
rect 449023 969 449035 972
rect 448977 963 449035 969
rect 462225 969 462237 972
rect 462271 969 462283 1003
rect 462225 963 462283 969
rect 404725 935 404783 941
rect 370792 904 377168 932
rect 247957 799 248015 805
rect 247957 765 247969 799
rect 248003 796 248015 799
rect 340877 799 340935 805
rect 248003 768 253520 796
rect 248003 765 248015 768
rect 247957 759 248015 765
rect 4062 688 4068 740
rect 4120 728 4126 740
rect 4120 700 5534 728
rect 4120 688 4126 700
rect 1670 620 1676 672
rect 1728 660 1734 672
rect 5350 660 5356 672
rect 1728 632 5356 660
rect 1728 620 1734 632
rect 5350 620 5356 632
rect 5408 620 5414 672
rect 5506 660 5534 700
rect 245764 700 251220 728
rect 245764 672 245792 700
rect 7742 660 7748 672
rect 5506 632 7748 660
rect 7742 620 7748 632
rect 7800 620 7806 672
rect 11054 620 11060 672
rect 11112 660 11118 672
rect 14458 660 14464 672
rect 11112 632 14464 660
rect 11112 620 11118 632
rect 14458 620 14464 632
rect 14516 620 14522 672
rect 19426 620 19432 672
rect 19484 660 19490 672
rect 22370 660 22376 672
rect 19484 632 22376 660
rect 19484 620 19490 632
rect 22370 620 22376 632
rect 22428 620 22434 672
rect 23014 620 23020 672
rect 23072 660 23078 672
rect 25774 660 25780 672
rect 23072 632 25780 660
rect 23072 620 23078 632
rect 25774 620 25780 632
rect 25832 620 25838 672
rect 28810 620 28816 672
rect 28868 660 28874 672
rect 31662 660 31668 672
rect 28868 632 31668 660
rect 28868 620 28874 632
rect 31662 620 31668 632
rect 31720 620 31726 672
rect 32398 620 32404 672
rect 32456 660 32462 672
rect 34882 660 34888 672
rect 32456 632 34888 660
rect 32456 620 32462 632
rect 34882 620 34888 632
rect 34940 620 34946 672
rect 38378 620 38384 672
rect 38436 660 38442 672
rect 38436 632 39804 660
rect 38436 620 38442 632
rect 566 552 572 604
rect 624 592 630 604
rect 4246 592 4252 604
rect 624 564 4252 592
rect 624 552 630 564
rect 4246 552 4252 564
rect 4304 552 4310 604
rect 5258 552 5264 604
rect 5316 592 5322 604
rect 6181 595 6239 601
rect 6181 592 6193 595
rect 5316 564 6193 592
rect 5316 552 5322 564
rect 6181 561 6193 564
rect 6227 561 6239 595
rect 6181 555 6239 561
rect 6454 552 6460 604
rect 6512 552 6518 604
rect 7650 552 7656 604
rect 7708 592 7714 604
rect 7708 564 10456 592
rect 7708 552 7714 564
rect 6472 524 6500 552
rect 10318 524 10324 536
rect 6472 496 10324 524
rect 10318 484 10324 496
rect 10376 484 10382 536
rect 10428 524 10456 564
rect 12342 552 12348 604
rect 12400 592 12406 604
rect 15562 592 15568 604
rect 12400 564 15568 592
rect 12400 552 12406 564
rect 15562 552 15568 564
rect 15620 552 15626 604
rect 18506 552 18512 604
rect 18564 592 18570 604
rect 21266 592 21272 604
rect 18564 564 21272 592
rect 18564 552 18570 564
rect 21266 552 21272 564
rect 21324 552 21330 604
rect 21818 552 21824 604
rect 21876 592 21882 604
rect 24854 592 24860 604
rect 21876 564 24860 592
rect 21876 552 21882 564
rect 24854 552 24860 564
rect 24912 552 24918 604
rect 25314 552 25320 604
rect 25372 592 25378 604
rect 28074 592 28080 604
rect 25372 564 28080 592
rect 25372 552 25378 564
rect 28074 552 28080 564
rect 28132 552 28138 604
rect 28718 552 28724 604
rect 28776 592 28782 604
rect 29178 592 29184 604
rect 28776 564 29184 592
rect 28776 552 28782 564
rect 29178 552 29184 564
rect 29236 552 29242 604
rect 30098 552 30104 604
rect 30156 592 30162 604
rect 32582 592 32588 604
rect 30156 564 32588 592
rect 30156 552 30162 564
rect 32582 552 32588 564
rect 32640 552 32646 604
rect 33594 552 33600 604
rect 33652 592 33658 604
rect 36078 592 36084 604
rect 33652 564 36084 592
rect 33652 552 33658 564
rect 36078 552 36084 564
rect 36136 552 36142 604
rect 37182 552 37188 604
rect 37240 592 37246 604
rect 37240 564 38654 592
rect 37240 552 37246 564
rect 11514 524 11520 536
rect 10428 496 11520 524
rect 11514 484 11520 496
rect 11572 484 11578 536
rect 13354 484 13360 536
rect 13412 524 13418 536
rect 16666 524 16672 536
rect 13412 496 16672 524
rect 13412 484 13418 496
rect 16666 484 16672 496
rect 16724 484 16730 536
rect 31478 484 31484 536
rect 31536 524 31542 536
rect 33778 524 33784 536
rect 31536 496 33784 524
rect 31536 484 31542 496
rect 33778 484 33784 496
rect 33836 484 33842 536
rect 3234 416 3240 468
rect 3292 456 3298 468
rect 6638 456 6644 468
rect 3292 428 6644 456
rect 3292 416 3298 428
rect 6638 416 6644 428
rect 6696 416 6702 468
rect 24854 416 24860 468
rect 24912 456 24918 468
rect 26878 456 26884 468
rect 24912 428 26884 456
rect 24912 416 24918 428
rect 26878 416 26884 428
rect 26936 416 26942 468
rect 6181 391 6239 397
rect 6181 357 6193 391
rect 6227 388 6239 391
rect 8938 388 8944 400
rect 6227 360 8944 388
rect 6227 357 6239 360
rect 6181 351 6239 357
rect 8938 348 8944 360
rect 8996 348 9002 400
rect 14550 348 14556 400
rect 14608 388 14614 400
rect 17862 388 17868 400
rect 14608 360 17868 388
rect 14608 348 14614 360
rect 17862 348 17868 360
rect 17920 348 17926 400
rect 38626 388 38654 564
rect 39574 552 39580 604
rect 39632 552 39638 604
rect 39776 592 39804 632
rect 40678 620 40684 672
rect 40736 660 40742 672
rect 42794 660 42800 672
rect 40736 632 42800 660
rect 40736 620 40742 632
rect 42794 620 42800 632
rect 42852 620 42858 672
rect 46658 620 46664 672
rect 46716 660 46722 672
rect 48498 660 48504 672
rect 46716 632 48504 660
rect 46716 620 46722 632
rect 48498 620 48504 632
rect 48556 620 48562 672
rect 48958 620 48964 672
rect 49016 660 49022 672
rect 50798 660 50804 672
rect 49016 632 50804 660
rect 49016 620 49022 632
rect 50798 620 50804 632
rect 50856 620 50862 672
rect 63218 620 63224 672
rect 63276 660 63282 672
rect 63276 632 63494 660
rect 63276 620 63282 632
rect 40770 592 40776 604
rect 39776 564 40776 592
rect 40770 552 40776 564
rect 40828 552 40834 604
rect 41874 552 41880 604
rect 41932 592 41938 604
rect 43990 592 43996 604
rect 41932 564 43996 592
rect 41932 552 41938 564
rect 43990 552 43996 564
rect 44048 552 44054 604
rect 47854 552 47860 604
rect 47912 592 47918 604
rect 49602 592 49608 604
rect 47912 564 49608 592
rect 47912 552 47918 564
rect 49602 552 49608 564
rect 49660 552 49666 604
rect 50154 552 50160 604
rect 50212 552 50218 604
rect 51350 552 51356 604
rect 51408 592 51414 604
rect 53006 592 53012 604
rect 51408 564 53012 592
rect 51408 552 51414 564
rect 53006 552 53012 564
rect 53064 552 53070 604
rect 54938 552 54944 604
rect 54996 592 55002 604
rect 56410 592 56416 604
rect 54996 564 56416 592
rect 54996 552 55002 564
rect 56410 552 56416 564
rect 56468 552 56474 604
rect 62022 552 62028 604
rect 62080 592 62086 604
rect 63310 592 63316 604
rect 62080 564 63316 592
rect 62080 552 62086 564
rect 63310 552 63316 564
rect 63368 552 63374 604
rect 63466 592 63494 632
rect 64322 620 64328 672
rect 64380 660 64386 672
rect 65610 660 65616 672
rect 64380 632 65616 660
rect 64380 620 64386 632
rect 65610 620 65616 632
rect 65668 620 65674 672
rect 66714 620 66720 672
rect 66772 660 66778 672
rect 68002 660 68008 672
rect 66772 632 68008 660
rect 66772 620 66778 632
rect 68002 620 68008 632
rect 68060 620 68066 672
rect 69106 620 69112 672
rect 69164 660 69170 672
rect 70578 660 70584 672
rect 69164 632 70584 660
rect 69164 620 69170 632
rect 70578 620 70584 632
rect 70636 620 70642 672
rect 133230 620 133236 672
rect 133288 660 133294 672
rect 134150 660 134156 672
rect 133288 632 134156 660
rect 133288 620 133294 632
rect 134150 620 134156 632
rect 134208 620 134214 672
rect 136174 620 136180 672
rect 136232 660 136238 672
rect 137646 660 137652 672
rect 136232 632 137652 660
rect 136232 620 136238 632
rect 137646 620 137652 632
rect 137704 620 137710 672
rect 138750 620 138756 672
rect 138808 660 138814 672
rect 140038 660 140044 672
rect 138808 632 140044 660
rect 138808 620 138814 632
rect 140038 620 140044 632
rect 140096 620 140102 672
rect 151354 620 151360 672
rect 151412 660 151418 672
rect 153010 660 153016 672
rect 151412 632 153016 660
rect 151412 620 151418 632
rect 153010 620 153016 632
rect 153068 620 153074 672
rect 153654 620 153660 672
rect 153712 660 153718 672
rect 155402 660 155408 672
rect 153712 632 155408 660
rect 153712 620 153718 632
rect 155402 620 155408 632
rect 155460 620 155466 672
rect 162762 620 162768 672
rect 162820 660 162826 672
rect 164878 660 164884 672
rect 162820 632 164884 660
rect 162820 620 162826 632
rect 164878 620 164884 632
rect 164936 620 164942 672
rect 166074 660 166080 672
rect 165908 632 166080 660
rect 64414 592 64420 604
rect 63466 564 64420 592
rect 64414 552 64420 564
rect 64472 552 64478 604
rect 65518 552 65524 604
rect 65576 592 65582 604
rect 66806 592 66812 604
rect 65576 564 66812 592
rect 65576 552 65582 564
rect 66806 552 66812 564
rect 66864 552 66870 604
rect 70302 552 70308 604
rect 70360 592 70366 604
rect 71222 592 71228 604
rect 70360 564 71228 592
rect 70360 552 70366 564
rect 71222 552 71228 564
rect 71280 552 71286 604
rect 76190 552 76196 604
rect 76248 592 76254 604
rect 76926 592 76932 604
rect 76248 564 76932 592
rect 76248 552 76254 564
rect 76926 552 76932 564
rect 76984 552 76990 604
rect 77386 552 77392 604
rect 77444 592 77450 604
rect 78030 592 78036 604
rect 77444 564 78036 592
rect 77444 552 77450 564
rect 78030 552 78036 564
rect 78088 552 78094 604
rect 78582 552 78588 604
rect 78640 592 78646 604
rect 79134 592 79140 604
rect 78640 564 79140 592
rect 78640 552 78646 564
rect 79134 552 79140 564
rect 79192 552 79198 604
rect 79686 552 79692 604
rect 79744 592 79750 604
rect 80330 592 80336 604
rect 79744 564 80336 592
rect 79744 552 79750 564
rect 80330 552 80336 564
rect 80388 552 80394 604
rect 80882 552 80888 604
rect 80940 592 80946 604
rect 81434 592 81440 604
rect 80940 564 81440 592
rect 80940 552 80946 564
rect 81434 552 81440 564
rect 81492 552 81498 604
rect 82078 552 82084 604
rect 82136 592 82142 604
rect 82722 592 82728 604
rect 82136 564 82728 592
rect 82136 552 82142 564
rect 82722 552 82728 564
rect 82780 552 82786 604
rect 121822 552 121828 604
rect 121880 592 121886 604
rect 122282 592 122288 604
rect 121880 564 122288 592
rect 121880 552 121886 564
rect 122282 552 122288 564
rect 122340 552 122346 604
rect 124122 552 124128 604
rect 124180 592 124186 604
rect 124674 592 124680 604
rect 124180 564 124680 592
rect 124180 552 124186 564
rect 124674 552 124680 564
rect 124732 552 124738 604
rect 125226 552 125232 604
rect 125284 592 125290 604
rect 125870 592 125876 604
rect 125284 564 125876 592
rect 125284 552 125290 564
rect 125870 552 125876 564
rect 125928 552 125934 604
rect 126422 552 126428 604
rect 126480 592 126486 604
rect 126974 592 126980 604
rect 126480 564 126980 592
rect 126480 552 126486 564
rect 126974 552 126980 564
rect 127032 552 127038 604
rect 127526 552 127532 604
rect 127584 592 127590 604
rect 128170 592 128176 604
rect 127584 564 128176 592
rect 127584 552 127590 564
rect 128170 552 128176 564
rect 128228 552 128234 604
rect 128630 552 128636 604
rect 128688 592 128694 604
rect 129366 592 129372 604
rect 128688 564 129372 592
rect 128688 552 128694 564
rect 129366 552 129372 564
rect 129424 552 129430 604
rect 133874 552 133880 604
rect 133932 592 133938 604
rect 135254 592 135260 604
rect 133932 564 135260 592
rect 133932 552 133938 564
rect 135254 552 135260 564
rect 135312 552 135318 604
rect 136450 552 136456 604
rect 136508 552 136514 604
rect 137554 552 137560 604
rect 137612 592 137618 604
rect 138842 592 138848 604
rect 137612 564 138848 592
rect 137612 552 137618 564
rect 138842 552 138848 564
rect 138900 552 138906 604
rect 139946 552 139952 604
rect 140004 592 140010 604
rect 141234 592 141240 604
rect 140004 564 141240 592
rect 140004 552 140010 564
rect 141234 552 141240 564
rect 141292 552 141298 604
rect 144546 552 144552 604
rect 144604 592 144610 604
rect 145926 592 145932 604
rect 144604 564 145932 592
rect 144604 552 144610 564
rect 145926 552 145932 564
rect 145984 552 145990 604
rect 146846 552 146852 604
rect 146904 592 146910 604
rect 148318 592 148324 604
rect 146904 564 148324 592
rect 146904 552 146910 564
rect 148318 552 148324 564
rect 148376 552 148382 604
rect 152550 552 152556 604
rect 152608 592 152614 604
rect 154206 592 154212 604
rect 152608 564 154212 592
rect 152608 552 152614 564
rect 154206 552 154212 564
rect 154264 552 154270 604
rect 154758 552 154764 604
rect 154816 592 154822 604
rect 156598 592 156604 604
rect 154816 564 156604 592
rect 154816 552 154822 564
rect 156598 552 156604 564
rect 156656 552 156662 604
rect 157058 552 157064 604
rect 157116 592 157122 604
rect 158898 592 158904 604
rect 157116 564 158904 592
rect 157116 552 157122 564
rect 158898 552 158904 564
rect 158956 552 158962 604
rect 161566 552 161572 604
rect 161624 592 161630 604
rect 163682 592 163688 604
rect 161624 564 163688 592
rect 161624 552 161630 564
rect 163682 552 163688 564
rect 163740 552 163746 604
rect 39592 456 39620 552
rect 50172 524 50200 552
rect 51902 524 51908 536
rect 50172 496 51908 524
rect 51902 484 51908 496
rect 51960 484 51966 536
rect 67726 484 67732 536
rect 67784 524 67790 536
rect 69382 524 69388 536
rect 67784 496 69388 524
rect 67784 484 67790 496
rect 69382 484 69388 496
rect 69440 484 69446 536
rect 134978 484 134984 536
rect 135036 524 135042 536
rect 136468 524 136496 552
rect 135036 496 136496 524
rect 135036 484 135042 496
rect 141050 484 141056 536
rect 141108 524 141114 536
rect 142062 524 142068 536
rect 141108 496 142068 524
rect 141108 484 141114 496
rect 142062 484 142068 496
rect 142120 484 142126 536
rect 158162 484 158168 536
rect 158220 524 158226 536
rect 159726 524 159732 536
rect 158220 496 159732 524
rect 158220 484 158226 496
rect 159726 484 159732 496
rect 159784 484 159790 536
rect 42150 456 42156 468
rect 39592 428 42156 456
rect 42150 416 42156 428
rect 42208 416 42214 468
rect 163406 416 163412 468
rect 163464 456 163470 468
rect 165908 456 165936 632
rect 166074 620 166080 632
rect 166132 620 166138 672
rect 167086 620 167092 672
rect 167144 660 167150 672
rect 169570 660 169576 672
rect 167144 632 169576 660
rect 167144 620 167150 632
rect 169570 620 169576 632
rect 169628 620 169634 672
rect 180886 620 180892 672
rect 180944 660 180950 672
rect 183738 660 183744 672
rect 180944 632 183744 660
rect 180944 620 180950 632
rect 183738 620 183744 632
rect 183796 620 183802 672
rect 186130 660 186136 672
rect 184216 632 186136 660
rect 165982 552 165988 604
rect 166040 592 166046 604
rect 168374 592 168380 604
rect 166040 564 168380 592
rect 166040 552 166046 564
rect 168374 552 168380 564
rect 168432 552 168438 604
rect 170674 552 170680 604
rect 170732 592 170738 604
rect 173158 592 173164 604
rect 170732 564 173164 592
rect 170732 552 170738 564
rect 173158 552 173164 564
rect 173216 552 173222 604
rect 179782 552 179788 604
rect 179840 592 179846 604
rect 182542 592 182548 604
rect 179840 564 182548 592
rect 179840 552 179846 564
rect 182542 552 182548 564
rect 182600 552 182606 604
rect 183186 552 183192 604
rect 183244 592 183250 604
rect 184216 592 184244 632
rect 186130 620 186136 632
rect 186188 620 186194 672
rect 191098 620 191104 672
rect 191156 660 191162 672
rect 194410 660 194416 672
rect 191156 632 194416 660
rect 191156 620 191162 632
rect 194410 620 194416 632
rect 194468 620 194474 672
rect 211614 620 211620 672
rect 211672 660 211678 672
rect 215662 660 215668 672
rect 211672 632 215668 660
rect 211672 620 211678 632
rect 215662 620 215668 632
rect 215720 620 215726 672
rect 220170 620 220176 672
rect 220228 660 220234 672
rect 225322 660 225328 672
rect 220228 632 225328 660
rect 220228 620 220234 632
rect 225322 620 225328 632
rect 225380 620 225386 672
rect 226150 620 226156 672
rect 226208 660 226214 672
rect 231026 660 231032 672
rect 226208 632 231032 660
rect 226208 620 226214 632
rect 231026 620 231032 632
rect 231084 620 231090 672
rect 234614 660 234620 672
rect 231780 632 234620 660
rect 183244 564 184244 592
rect 183244 552 183250 564
rect 189994 552 190000 604
rect 190052 592 190058 604
rect 193214 592 193220 604
rect 190052 564 193220 592
rect 190052 552 190058 564
rect 193214 552 193220 564
rect 193272 552 193278 604
rect 196802 552 196808 604
rect 196860 552 196866 604
rect 199102 592 199108 604
rect 198706 564 199108 592
rect 187694 484 187700 536
rect 187752 524 187758 536
rect 191006 524 191012 536
rect 187752 496 191012 524
rect 187752 484 187758 496
rect 191006 484 191012 496
rect 191064 484 191070 536
rect 192938 484 192944 536
rect 192996 524 193002 536
rect 196820 524 196848 552
rect 192996 496 196848 524
rect 192996 484 193002 496
rect 163464 428 165936 456
rect 163464 416 163470 428
rect 39850 388 39856 400
rect 38626 360 39856 388
rect 39850 348 39856 360
rect 39908 348 39914 400
rect 42886 348 42892 400
rect 42944 388 42950 400
rect 45094 388 45100 400
rect 42944 360 45100 388
rect 42944 348 42950 360
rect 45094 348 45100 360
rect 45152 348 45158 400
rect 71314 348 71320 400
rect 71372 388 71378 400
rect 72326 388 72332 400
rect 71372 360 72332 388
rect 71372 348 71378 360
rect 72326 348 72332 360
rect 72384 348 72390 400
rect 72418 348 72424 400
rect 72476 388 72482 400
rect 73522 388 73528 400
rect 72476 360 73528 388
rect 72476 348 72482 360
rect 73522 348 73528 360
rect 73580 348 73586 400
rect 73614 348 73620 400
rect 73672 388 73678 400
rect 74626 388 74632 400
rect 73672 360 74632 388
rect 73672 348 73678 360
rect 74626 348 74632 360
rect 74684 348 74690 400
rect 130930 348 130936 400
rect 130988 388 130994 400
rect 131942 388 131948 400
rect 130988 360 131948 388
rect 130988 348 130994 360
rect 131942 348 131948 360
rect 132000 348 132006 400
rect 132034 348 132040 400
rect 132092 388 132098 400
rect 133138 388 133144 400
rect 132092 360 133144 388
rect 132092 348 132098 360
rect 133138 348 133144 360
rect 133196 348 133202 400
rect 160462 348 160468 400
rect 160520 388 160526 400
rect 162670 388 162676 400
rect 160520 360 162676 388
rect 160520 348 160526 360
rect 162670 348 162676 360
rect 162728 348 162734 400
rect 188798 348 188804 400
rect 188856 388 188862 400
rect 192202 388 192208 400
rect 188856 360 192208 388
rect 188856 348 188862 360
rect 192202 348 192208 360
rect 192260 348 192266 400
rect 195238 348 195244 400
rect 195296 388 195302 400
rect 198706 388 198734 564
rect 199102 552 199108 564
rect 199160 552 199166 604
rect 203610 552 203616 604
rect 203668 592 203674 604
rect 204162 592 204168 604
rect 203668 564 204168 592
rect 203668 552 203674 564
rect 204162 552 204168 564
rect 204220 552 204226 604
rect 205726 552 205732 604
rect 205784 592 205790 604
rect 209774 592 209780 604
rect 205784 564 209780 592
rect 205784 552 205790 564
rect 209774 552 209780 564
rect 209832 552 209838 604
rect 210418 552 210424 604
rect 210476 592 210482 604
rect 212077 595 212135 601
rect 212077 592 212089 595
rect 210476 564 212089 592
rect 210476 552 210482 564
rect 212077 561 212089 564
rect 212123 561 212135 595
rect 212077 555 212135 561
rect 212166 552 212172 604
rect 212224 552 212230 604
rect 212261 595 212319 601
rect 212261 561 212273 595
rect 212307 592 212319 595
rect 214466 592 214472 604
rect 212307 564 214472 592
rect 212307 561 212319 564
rect 212261 555 212319 561
rect 214466 552 214472 564
rect 214524 552 214530 604
rect 219526 552 219532 604
rect 219584 592 219590 604
rect 223942 592 223948 604
rect 219584 564 223948 592
rect 219584 552 219590 564
rect 223942 552 223948 564
rect 224000 552 224006 604
rect 225046 552 225052 604
rect 225104 592 225110 604
rect 229830 592 229836 604
rect 225104 564 227714 592
rect 225104 552 225110 564
rect 208394 484 208400 536
rect 208452 524 208458 536
rect 212184 524 212212 552
rect 208452 496 212212 524
rect 208452 484 208458 496
rect 218422 484 218428 536
rect 218480 524 218486 536
rect 222930 524 222936 536
rect 218480 496 222936 524
rect 218480 484 218486 496
rect 222930 484 222936 496
rect 222988 484 222994 536
rect 227346 484 227352 536
rect 227404 484 227410 536
rect 227686 524 227714 564
rect 229066 564 229836 592
rect 229066 524 229094 564
rect 229830 552 229836 564
rect 229888 552 229894 604
rect 227686 496 229094 524
rect 229646 484 229652 536
rect 229704 524 229710 536
rect 231780 524 231808 632
rect 234614 620 234620 632
rect 234672 620 234678 672
rect 235442 620 235448 672
rect 235500 660 235506 672
rect 240502 660 240508 672
rect 235500 632 240508 660
rect 235500 620 235506 632
rect 240502 620 240508 632
rect 240560 620 240566 672
rect 241146 620 241152 672
rect 241204 660 241210 672
rect 241204 632 245700 660
rect 241204 620 241210 632
rect 231854 552 231860 604
rect 231912 592 231918 604
rect 237006 592 237012 604
rect 231912 564 237012 592
rect 231912 552 231918 564
rect 237006 552 237012 564
rect 237064 552 237070 604
rect 238110 552 238116 604
rect 238168 552 238174 604
rect 238846 552 238852 604
rect 238904 592 238910 604
rect 244090 592 244096 604
rect 238904 564 244096 592
rect 238904 552 238910 564
rect 244090 552 244096 564
rect 244148 552 244154 604
rect 245194 592 245200 604
rect 244476 564 245200 592
rect 229704 496 231808 524
rect 229704 484 229710 496
rect 233142 484 233148 536
rect 233200 524 233206 536
rect 238128 524 238156 552
rect 233200 496 238156 524
rect 233200 484 233206 496
rect 239950 484 239956 536
rect 240008 524 240014 536
rect 244476 524 244504 564
rect 245194 552 245200 564
rect 245252 552 245258 604
rect 245672 592 245700 632
rect 245746 620 245752 672
rect 245804 620 245810 672
rect 247954 660 247960 672
rect 247915 632 247960 660
rect 247954 620 247960 632
rect 248012 620 248018 672
rect 251192 604 251220 700
rect 253492 672 253520 768
rect 309980 768 315528 796
rect 284404 700 288388 728
rect 253474 620 253480 672
rect 253532 620 253538 672
rect 254578 620 254584 672
rect 254636 660 254642 672
rect 254636 632 257200 660
rect 254636 620 254642 632
rect 246022 592 246028 604
rect 245672 564 246028 592
rect 246022 552 246028 564
rect 246080 552 246086 604
rect 249978 592 249984 604
rect 247006 564 249984 592
rect 240008 496 244504 524
rect 240008 484 240014 496
rect 244550 484 244556 536
rect 244608 524 244614 536
rect 247006 524 247034 564
rect 249978 552 249984 564
rect 250036 552 250042 604
rect 251174 552 251180 604
rect 251232 552 251238 604
rect 252370 592 252376 604
rect 252331 564 252376 592
rect 252370 552 252376 564
rect 252428 552 252434 604
rect 254670 552 254676 604
rect 254728 552 254734 604
rect 254765 595 254823 601
rect 254765 561 254777 595
rect 254811 592 254823 595
rect 257062 592 257068 604
rect 254811 564 257068 592
rect 254811 561 254823 564
rect 254765 555 254823 561
rect 257062 552 257068 564
rect 257120 552 257126 604
rect 257172 592 257200 632
rect 257246 620 257252 672
rect 257304 660 257310 672
rect 258258 660 258264 672
rect 257304 632 258264 660
rect 257304 620 257310 632
rect 258258 620 258264 632
rect 258316 620 258322 672
rect 260466 620 260472 672
rect 260524 660 260530 672
rect 266538 660 266544 672
rect 260524 632 266544 660
rect 260524 620 260530 632
rect 266538 620 266544 632
rect 266596 620 266602 672
rect 268838 660 268844 672
rect 267660 632 268844 660
rect 260650 592 260656 604
rect 257172 564 260656 592
rect 260650 552 260656 564
rect 260708 552 260714 604
rect 262674 552 262680 604
rect 262732 592 262738 604
rect 267660 592 267688 632
rect 268838 620 268844 632
rect 268896 620 268902 672
rect 272886 620 272892 672
rect 272944 660 272950 672
rect 272944 632 277440 660
rect 272944 620 272950 632
rect 262732 564 267688 592
rect 262732 552 262738 564
rect 267734 552 267740 604
rect 267792 552 267798 604
rect 270034 592 270040 604
rect 268212 564 270040 592
rect 244608 496 247034 524
rect 244608 484 244614 496
rect 249058 484 249064 536
rect 249116 524 249122 536
rect 254688 524 254716 552
rect 249116 496 254716 524
rect 249116 484 249122 496
rect 261570 484 261576 536
rect 261628 524 261634 536
rect 267752 524 267780 552
rect 261628 496 267780 524
rect 261628 484 261634 496
rect 212534 416 212540 468
rect 212592 456 212598 468
rect 216582 456 216588 468
rect 212592 428 216588 456
rect 212592 416 212598 428
rect 216582 416 216588 428
rect 216640 416 216646 468
rect 222470 416 222476 468
rect 222528 456 222534 468
rect 227364 456 227392 484
rect 222528 428 227392 456
rect 222528 416 222534 428
rect 234338 416 234344 468
rect 234396 456 234402 468
rect 239030 456 239036 468
rect 234396 428 239036 456
rect 234396 416 234402 428
rect 239030 416 239036 428
rect 239088 416 239094 468
rect 253106 416 253112 468
rect 253164 456 253170 468
rect 259086 456 259092 468
rect 253164 428 259092 456
rect 253164 416 253170 428
rect 259086 416 259092 428
rect 259144 416 259150 468
rect 263686 416 263692 468
rect 263744 456 263750 468
rect 268212 456 268240 564
rect 270034 552 270040 564
rect 270092 552 270098 604
rect 270678 552 270684 604
rect 270736 592 270742 604
rect 276750 592 276756 604
rect 270736 564 276756 592
rect 270736 552 270742 564
rect 276750 552 276756 564
rect 276808 552 276814 604
rect 277412 592 277440 632
rect 277486 620 277492 672
rect 277544 660 277550 672
rect 284294 660 284300 672
rect 277544 632 284300 660
rect 277544 620 277550 632
rect 284294 620 284300 632
rect 284352 620 284358 672
rect 279510 592 279516 604
rect 277412 564 279516 592
rect 279510 552 279516 564
rect 279568 552 279574 604
rect 280706 592 280712 604
rect 280667 564 280712 592
rect 280706 552 280712 564
rect 280764 552 280770 604
rect 281810 552 281816 604
rect 281868 592 281874 604
rect 284404 592 284432 700
rect 286594 660 286600 672
rect 285646 632 286600 660
rect 281868 564 284432 592
rect 281868 552 281874 564
rect 285398 552 285404 604
rect 285456 552 285462 604
rect 268378 484 268384 536
rect 268436 524 268442 536
rect 274542 524 274548 536
rect 268436 496 274548 524
rect 268436 484 268442 496
rect 274542 484 274548 496
rect 274600 484 274606 536
rect 278590 484 278596 536
rect 278648 524 278654 536
rect 285416 524 285444 552
rect 278648 496 285444 524
rect 278648 484 278654 496
rect 263744 428 268240 456
rect 263744 416 263750 428
rect 269482 416 269488 468
rect 269540 456 269546 468
rect 276198 456 276204 468
rect 269540 428 276204 456
rect 269540 416 269546 428
rect 276198 416 276204 428
rect 276256 416 276262 468
rect 279234 416 279240 468
rect 279292 456 279298 468
rect 285646 456 285674 632
rect 286594 620 286600 632
rect 286652 620 286658 672
rect 288360 660 288388 700
rect 292546 700 298508 728
rect 288986 660 288992 672
rect 288360 632 288992 660
rect 288986 620 288992 632
rect 289044 620 289050 672
rect 291102 620 291108 672
rect 291160 660 291166 672
rect 292546 660 292574 700
rect 298480 672 298508 700
rect 309980 672 310008 768
rect 310118 700 315436 728
rect 291160 632 292574 660
rect 291160 620 291166 632
rect 293402 620 293408 672
rect 293460 660 293466 672
rect 293460 632 295564 660
rect 293460 620 293466 632
rect 287606 552 287612 604
rect 287664 592 287670 604
rect 294874 592 294880 604
rect 287664 564 294880 592
rect 287664 552 287670 564
rect 294874 552 294880 564
rect 294932 552 294938 604
rect 294506 484 294512 536
rect 294564 524 294570 536
rect 295536 524 295564 632
rect 298462 620 298468 672
rect 298520 620 298526 672
rect 300210 620 300216 672
rect 300268 660 300274 672
rect 300268 632 304304 660
rect 300268 620 300274 632
rect 295610 552 295616 604
rect 295668 592 295674 604
rect 303154 592 303160 604
rect 295668 564 303160 592
rect 295668 552 295674 564
rect 303154 552 303160 564
rect 303212 552 303218 604
rect 304276 592 304304 632
rect 307662 620 307668 672
rect 307720 660 307726 672
rect 307720 632 309916 660
rect 307720 620 307726 632
rect 307938 592 307944 604
rect 304276 564 307944 592
rect 307938 552 307944 564
rect 307996 552 308002 604
rect 309042 552 309048 604
rect 309100 552 309106 604
rect 309888 592 309916 632
rect 309962 620 309968 672
rect 310020 620 310026 672
rect 310118 592 310146 700
rect 310238 592 310244 604
rect 309888 564 310146 592
rect 310199 564 310244 592
rect 310238 552 310244 564
rect 310296 552 310302 604
rect 311434 552 311440 604
rect 311492 552 311498 604
rect 312630 592 312636 604
rect 312591 564 312636 592
rect 312630 552 312636 564
rect 312688 552 312694 604
rect 300578 524 300584 536
rect 294564 496 295334 524
rect 295536 496 300584 524
rect 294564 484 294570 496
rect 279292 428 285674 456
rect 279292 416 279298 428
rect 288802 416 288808 468
rect 288860 456 288866 468
rect 294598 456 294604 468
rect 288860 428 294604 456
rect 288860 416 288866 428
rect 294598 416 294604 428
rect 294656 416 294662 468
rect 295306 456 295334 496
rect 300578 484 300584 496
rect 300636 484 300642 536
rect 301314 484 301320 536
rect 301372 524 301378 536
rect 309060 524 309088 552
rect 301372 496 309088 524
rect 301372 484 301378 496
rect 301774 456 301780 468
rect 295306 428 301780 456
rect 301774 416 301780 428
rect 301832 416 301838 468
rect 303614 416 303620 468
rect 303672 456 303678 468
rect 311452 456 311480 552
rect 315408 524 315436 700
rect 315500 592 315528 768
rect 340877 765 340889 799
rect 340923 796 340935 799
rect 340923 768 347728 796
rect 340923 765 340935 768
rect 340877 759 340935 765
rect 316006 700 321554 728
rect 316006 672 316034 700
rect 315942 620 315948 672
rect 316000 632 316034 672
rect 318518 660 318524 672
rect 316144 632 318524 660
rect 316000 620 316006 632
rect 316144 592 316172 632
rect 318518 620 318524 632
rect 318576 620 318582 672
rect 321526 660 321554 700
rect 335372 700 343634 728
rect 335372 672 335400 700
rect 324406 660 324412 672
rect 321526 632 324412 660
rect 324406 620 324412 632
rect 324464 620 324470 672
rect 325142 620 325148 672
rect 325200 660 325206 672
rect 333606 660 333612 672
rect 325200 632 333612 660
rect 325200 620 325206 632
rect 333606 620 333612 632
rect 333664 620 333670 672
rect 335354 620 335360 672
rect 335412 620 335418 672
rect 338666 660 338672 672
rect 336016 632 338672 660
rect 315500 564 316172 592
rect 316218 552 316224 604
rect 316276 552 316282 604
rect 317138 552 317144 604
rect 317196 592 317202 604
rect 325602 592 325608 604
rect 317196 564 325608 592
rect 317196 552 317202 564
rect 325602 552 325608 564
rect 325660 552 325666 604
rect 327442 552 327448 604
rect 327500 592 327506 604
rect 335909 595 335967 601
rect 335909 592 335921 595
rect 327500 564 335921 592
rect 327500 552 327506 564
rect 335909 561 335921 564
rect 335955 561 335967 595
rect 335909 555 335967 561
rect 316236 524 316264 552
rect 315408 496 316264 524
rect 319346 484 319352 536
rect 319404 524 319410 536
rect 327810 524 327816 536
rect 319404 496 327816 524
rect 319404 484 319410 496
rect 327810 484 327816 496
rect 327868 484 327874 536
rect 329742 484 329748 536
rect 329800 524 329806 536
rect 336016 524 336044 632
rect 338666 620 338672 632
rect 338724 620 338730 672
rect 340874 660 340880 672
rect 340835 632 340880 660
rect 340874 620 340880 632
rect 340932 620 340938 672
rect 343606 660 343634 700
rect 344554 660 344560 672
rect 343606 632 344560 660
rect 344554 620 344560 632
rect 344612 620 344618 672
rect 336093 595 336151 601
rect 336093 561 336105 595
rect 336139 592 336151 595
rect 339862 592 339868 604
rect 336139 564 339868 592
rect 336139 561 336151 564
rect 336093 555 336151 561
rect 339862 552 339868 564
rect 339920 552 339926 604
rect 342070 552 342076 604
rect 342128 592 342134 604
rect 347700 592 347728 768
rect 366085 731 366143 737
rect 366085 697 366097 731
rect 366131 728 366143 731
rect 370685 731 370743 737
rect 370685 728 370697 731
rect 366131 700 370697 728
rect 366131 697 366143 700
rect 366085 691 366143 697
rect 370685 697 370697 700
rect 370731 697 370743 731
rect 370685 691 370743 697
rect 347774 620 347780 672
rect 347832 660 347838 672
rect 349246 660 349252 672
rect 347832 632 349252 660
rect 347832 620 347838 632
rect 349246 620 349252 632
rect 349304 620 349310 672
rect 360838 660 360844 672
rect 351886 632 360844 660
rect 349062 592 349068 604
rect 342128 564 343634 592
rect 347700 564 349068 592
rect 342128 552 342134 564
rect 329800 496 336044 524
rect 343606 524 343634 564
rect 349062 552 349068 564
rect 349120 552 349126 604
rect 351270 552 351276 604
rect 351328 592 351334 604
rect 351886 592 351914 632
rect 360838 620 360844 632
rect 360896 620 360902 672
rect 364996 632 368336 660
rect 355226 592 355232 604
rect 351328 564 351914 592
rect 355187 564 355232 592
rect 351328 552 351334 564
rect 355226 552 355232 564
rect 355284 552 355290 604
rect 355870 552 355876 604
rect 355928 592 355934 604
rect 364797 595 364855 601
rect 364797 592 364809 595
rect 355928 564 364809 592
rect 355928 552 355934 564
rect 364797 561 364809 564
rect 364843 561 364855 595
rect 364797 555 364855 561
rect 351178 524 351184 536
rect 343606 496 351184 524
rect 329800 484 329806 496
rect 351178 484 351184 496
rect 351236 484 351242 536
rect 352466 484 352472 536
rect 352524 524 352530 536
rect 361942 524 361948 536
rect 352524 496 361948 524
rect 352524 484 352530 496
rect 361942 484 361948 496
rect 362000 484 362006 536
rect 303672 428 311480 456
rect 303672 416 303678 428
rect 312446 416 312452 468
rect 312504 456 312510 468
rect 320726 456 320732 468
rect 312504 428 320732 456
rect 312504 416 312510 428
rect 320726 416 320732 428
rect 320784 416 320790 468
rect 322842 416 322848 468
rect 322900 456 322906 468
rect 331214 456 331220 468
rect 322900 428 331220 456
rect 322900 416 322906 428
rect 331214 416 331220 428
rect 331272 416 331278 468
rect 331950 416 331956 468
rect 332008 456 332014 468
rect 341150 456 341156 468
rect 332008 428 341156 456
rect 332008 416 332014 428
rect 341150 416 341156 428
rect 341208 416 341214 468
rect 343174 416 343180 468
rect 343232 456 343238 468
rect 350626 456 350632 468
rect 343232 428 350632 456
rect 343232 416 343238 428
rect 350626 416 350632 428
rect 350684 416 350690 468
rect 353570 416 353576 468
rect 353628 456 353634 468
rect 353628 428 358814 456
rect 353628 416 353634 428
rect 195296 360 198734 388
rect 195296 348 195302 360
rect 217226 348 217232 400
rect 217284 388 217290 400
rect 221734 388 221740 400
rect 217284 360 221740 388
rect 217284 348 217290 360
rect 221734 348 221740 360
rect 221792 348 221798 400
rect 243354 348 243360 400
rect 243412 388 243418 400
rect 248966 388 248972 400
rect 243412 360 248972 388
rect 243412 348 243418 360
rect 248966 348 248972 360
rect 249024 348 249030 400
rect 250898 348 250904 400
rect 250956 388 250962 400
rect 254765 391 254823 397
rect 254765 388 254777 391
rect 250956 360 254777 388
rect 250956 348 250962 360
rect 254765 357 254777 360
rect 254811 357 254823 391
rect 254765 351 254823 357
rect 259270 348 259276 400
rect 259328 388 259334 400
rect 264974 388 264980 400
rect 259328 360 264980 388
rect 259328 348 259334 360
rect 264974 348 264980 360
rect 265032 348 265038 400
rect 271782 348 271788 400
rect 271840 388 271846 400
rect 278498 388 278504 400
rect 271840 360 278504 388
rect 271840 348 271846 360
rect 278498 348 278504 360
rect 278556 348 278562 400
rect 280430 348 280436 400
rect 280488 388 280494 400
rect 285674 388 285680 400
rect 280488 360 285680 388
rect 280488 348 280494 360
rect 285674 348 285680 360
rect 285732 348 285738 400
rect 299014 348 299020 400
rect 299072 388 299078 400
rect 306926 388 306932 400
rect 299072 360 306932 388
rect 299072 348 299078 360
rect 306926 348 306932 360
rect 306984 348 306990 400
rect 311066 348 311072 400
rect 311124 388 311130 400
rect 319530 388 319536 400
rect 311124 360 319536 388
rect 311124 348 311130 360
rect 319530 348 319536 360
rect 319588 348 319594 400
rect 321554 348 321560 400
rect 321612 388 321618 400
rect 330110 388 330116 400
rect 321612 360 330116 388
rect 321612 348 321618 360
rect 330110 348 330116 360
rect 330168 348 330174 400
rect 335909 391 335967 397
rect 335909 357 335921 391
rect 335955 388 335967 391
rect 336458 388 336464 400
rect 335955 360 336464 388
rect 335955 357 335967 360
rect 335909 351 335967 357
rect 336458 348 336464 360
rect 336516 348 336522 400
rect 336550 348 336556 400
rect 336608 388 336614 400
rect 345474 388 345480 400
rect 336608 360 345480 388
rect 336608 348 336614 360
rect 345474 348 345480 360
rect 345532 348 345538 400
rect 349062 348 349068 400
rect 349120 388 349126 400
rect 358446 388 358452 400
rect 349120 360 358452 388
rect 349120 348 349126 360
rect 358446 348 358452 360
rect 358504 348 358510 400
rect 246758 280 246764 332
rect 246816 320 246822 332
rect 252373 323 252431 329
rect 252373 320 252385 323
rect 246816 292 252385 320
rect 246816 280 246822 292
rect 252373 289 252385 292
rect 252419 289 252431 323
rect 252373 283 252431 289
rect 256878 280 256884 332
rect 256936 320 256942 332
rect 262766 320 262772 332
rect 256936 292 262772 320
rect 256936 280 256942 292
rect 262766 280 262772 292
rect 262824 280 262830 332
rect 275830 280 275836 332
rect 275888 320 275894 332
rect 283282 320 283288 332
rect 275888 292 283288 320
rect 275888 280 275894 292
rect 283282 280 283288 292
rect 283340 280 283346 332
rect 284110 280 284116 332
rect 284168 320 284174 332
rect 291194 320 291200 332
rect 284168 292 291200 320
rect 284168 280 284174 292
rect 291194 280 291200 292
rect 291252 280 291258 332
rect 296806 280 296812 332
rect 296864 320 296870 332
rect 303982 320 303988 332
rect 296864 292 303988 320
rect 296864 280 296870 292
rect 303982 280 303988 292
rect 304040 280 304046 332
rect 304718 280 304724 332
rect 304776 320 304782 332
rect 312633 323 312691 329
rect 312633 320 312645 323
rect 304776 292 312645 320
rect 304776 280 304782 292
rect 312633 289 312645 292
rect 312679 289 312691 323
rect 312633 283 312691 289
rect 318334 280 318340 332
rect 318392 320 318398 332
rect 326614 320 326620 332
rect 318392 292 326620 320
rect 318392 280 318398 292
rect 326614 280 326620 292
rect 326672 280 326678 332
rect 344370 280 344376 332
rect 344428 320 344434 332
rect 353846 320 353852 332
rect 344428 292 353852 320
rect 344428 280 344434 292
rect 353846 280 353852 292
rect 353904 280 353910 332
rect 354674 280 354680 332
rect 354732 320 354738 332
rect 358786 320 358814 428
rect 359274 416 359280 468
rect 359332 456 359338 468
rect 364996 456 365024 632
rect 365073 595 365131 601
rect 365073 561 365085 595
rect 365119 592 365131 595
rect 367002 592 367008 604
rect 365119 564 367008 592
rect 365119 561 365131 564
rect 365073 555 365131 561
rect 367002 552 367008 564
rect 367060 552 367066 604
rect 368198 592 368204 604
rect 368159 564 368204 592
rect 368198 552 368204 564
rect 368256 552 368262 604
rect 368308 592 368336 632
rect 369302 620 369308 672
rect 369360 660 369366 672
rect 370792 660 370820 904
rect 371988 836 377076 864
rect 369360 632 370820 660
rect 369360 620 369366 632
rect 371602 620 371608 672
rect 371660 660 371666 672
rect 371988 660 372016 836
rect 372065 799 372123 805
rect 372065 765 372077 799
rect 372111 796 372123 799
rect 372111 768 375328 796
rect 372111 765 372123 768
rect 372065 759 372123 765
rect 372801 731 372859 737
rect 372801 697 372813 731
rect 372847 728 372859 731
rect 372847 700 374316 728
rect 372847 697 372859 700
rect 372801 691 372859 697
rect 374288 672 374316 700
rect 375300 672 375328 768
rect 371660 632 372016 660
rect 371660 620 371666 632
rect 374270 620 374276 672
rect 374328 620 374334 672
rect 375282 620 375288 672
rect 375340 620 375346 672
rect 369394 592 369400 604
rect 368308 564 369400 592
rect 369394 552 369400 564
rect 369452 552 369458 604
rect 370590 592 370596 604
rect 370551 564 370596 592
rect 370590 552 370596 564
rect 370648 552 370654 604
rect 370685 595 370743 601
rect 370685 561 370697 595
rect 370731 592 370743 595
rect 376478 592 376484 604
rect 370731 564 376484 592
rect 370731 561 370743 564
rect 370685 555 370743 561
rect 376478 552 376484 564
rect 376536 552 376542 604
rect 377048 592 377076 836
rect 377140 660 377168 904
rect 404725 901 404737 935
rect 404771 932 404783 935
rect 437937 935 437995 941
rect 437937 932 437949 935
rect 404771 904 416728 932
rect 404771 901 404783 904
rect 404725 895 404783 901
rect 406473 867 406531 873
rect 406473 833 406485 867
rect 406519 864 406531 867
rect 406519 836 415440 864
rect 406519 833 406531 836
rect 406473 827 406531 833
rect 406565 799 406623 805
rect 406565 765 406577 799
rect 406611 796 406623 799
rect 406611 768 414336 796
rect 406611 765 406623 768
rect 406565 759 406623 765
rect 383105 731 383163 737
rect 383105 697 383117 731
rect 383151 728 383163 731
rect 383151 700 394280 728
rect 383151 697 383163 700
rect 383105 691 383163 697
rect 394252 672 394280 700
rect 400186 700 405734 728
rect 377950 660 377956 672
rect 377140 632 377956 660
rect 377950 620 377956 632
rect 378008 620 378014 672
rect 379514 620 379520 672
rect 379572 660 379578 672
rect 390278 660 390284 672
rect 379572 632 390284 660
rect 379572 620 379578 632
rect 390278 620 390284 632
rect 390336 620 390342 672
rect 394234 620 394240 672
rect 394292 620 394298 672
rect 395614 620 395620 672
rect 395672 660 395678 672
rect 400186 660 400214 700
rect 395672 632 400214 660
rect 395672 620 395678 632
rect 401134 620 401140 672
rect 401192 660 401198 672
rect 401192 632 404676 660
rect 401192 620 401198 632
rect 380158 592 380164 604
rect 377048 564 380164 592
rect 380158 552 380164 564
rect 380216 552 380222 604
rect 380802 552 380808 604
rect 380860 592 380866 604
rect 383102 592 383108 604
rect 380860 564 382274 592
rect 383063 564 383108 592
rect 380860 552 380866 564
rect 366082 524 366088 536
rect 366043 496 366088 524
rect 366082 484 366088 496
rect 366140 484 366146 536
rect 372801 527 372859 533
rect 372801 524 372813 527
rect 367066 496 372813 524
rect 359332 428 365024 456
rect 359332 416 359338 428
rect 366726 416 366732 468
rect 366784 456 366790 468
rect 367066 456 367094 496
rect 372801 493 372813 496
rect 372847 493 372859 527
rect 372801 487 372859 493
rect 373810 484 373816 536
rect 373868 524 373874 536
rect 380894 524 380900 536
rect 373868 496 380900 524
rect 373868 484 373874 496
rect 380894 484 380900 496
rect 380952 484 380958 536
rect 382246 524 382274 564
rect 383102 552 383108 564
rect 383160 552 383166 604
rect 389450 592 389456 604
rect 389411 564 389456 592
rect 389450 552 389456 564
rect 389508 552 389514 604
rect 389910 552 389916 604
rect 389968 592 389974 604
rect 392394 592 392400 604
rect 389968 564 392400 592
rect 389968 552 389974 564
rect 392394 552 392400 564
rect 392452 552 392458 604
rect 393314 552 393320 604
rect 393372 592 393378 604
rect 398009 595 398067 601
rect 398009 592 398021 595
rect 393372 564 398021 592
rect 393372 552 393378 564
rect 398009 561 398021 564
rect 398055 561 398067 595
rect 398009 555 398067 561
rect 398834 552 398840 604
rect 398892 592 398898 604
rect 404449 595 404507 601
rect 404449 592 404461 595
rect 398892 564 404461 592
rect 398892 552 398898 564
rect 404449 561 404461 564
rect 404495 561 404507 595
rect 404449 555 404507 561
rect 391566 524 391572 536
rect 382246 496 391572 524
rect 391566 484 391572 496
rect 391624 484 391630 536
rect 393777 527 393835 533
rect 393777 493 393789 527
rect 393823 524 393835 527
rect 399938 524 399944 536
rect 393823 496 399944 524
rect 393823 493 393835 496
rect 393777 487 393835 493
rect 399938 484 399944 496
rect 399996 484 400002 536
rect 400306 484 400312 536
rect 400364 524 400370 536
rect 403434 524 403440 536
rect 400364 496 403440 524
rect 400364 484 400370 496
rect 403434 484 403440 496
rect 403492 484 403498 536
rect 404648 524 404676 632
rect 404722 620 404728 672
rect 404780 660 404786 672
rect 404780 632 404825 660
rect 404780 620 404786 632
rect 404906 620 404912 672
rect 404964 660 404970 672
rect 405706 660 405734 700
rect 414308 672 414336 768
rect 407206 660 407212 672
rect 404964 632 405009 660
rect 405706 632 407212 660
rect 404964 620 404970 632
rect 407206 620 407212 632
rect 407264 620 407270 672
rect 411441 663 411499 669
rect 411441 629 411453 663
rect 411487 660 411499 663
rect 413738 660 413744 672
rect 411487 632 413232 660
rect 413699 632 413744 660
rect 411487 629 411499 632
rect 411441 623 411499 629
rect 404817 595 404875 601
rect 404817 561 404829 595
rect 404863 592 404875 595
rect 410794 592 410800 604
rect 404863 564 410800 592
rect 404863 561 404875 564
rect 404817 555 404875 561
rect 410794 552 410800 564
rect 410852 552 410858 604
rect 413094 552 413100 604
rect 413152 552 413158 604
rect 413204 592 413232 632
rect 413738 620 413744 632
rect 413796 620 413802 672
rect 414290 620 414296 672
rect 414348 620 414354 672
rect 415412 660 415440 836
rect 416700 672 416728 904
rect 437446 904 437949 932
rect 421653 867 421711 873
rect 421653 833 421665 867
rect 421699 864 421711 867
rect 432509 867 432567 873
rect 432509 864 432521 867
rect 421699 836 432521 864
rect 421699 833 421711 836
rect 421653 827 421711 833
rect 432509 833 432521 836
rect 432555 833 432567 867
rect 437446 864 437474 904
rect 437937 901 437949 904
rect 437983 901 437995 935
rect 437937 895 437995 901
rect 455417 935 455475 941
rect 455417 901 455429 935
rect 455463 932 455475 935
rect 461765 935 461823 941
rect 461765 932 461777 935
rect 455463 904 461777 932
rect 455463 901 455475 904
rect 455417 895 455475 901
rect 461765 901 461777 904
rect 461811 901 461823 935
rect 465736 932 465764 1040
rect 472805 1037 472817 1071
rect 472851 1068 472863 1071
rect 483753 1071 483811 1077
rect 472851 1040 483704 1068
rect 472851 1037 472863 1040
rect 472805 1031 472863 1037
rect 476577 1003 476635 1009
rect 476577 969 476589 1003
rect 476623 1000 476635 1003
rect 482833 1003 482891 1009
rect 482833 1000 482845 1003
rect 476623 972 482845 1000
rect 476623 969 476635 972
rect 476577 963 476635 969
rect 482833 969 482845 972
rect 482879 969 482891 1003
rect 483676 1000 483704 1040
rect 483753 1037 483765 1071
rect 483799 1068 483811 1071
rect 499393 1071 499451 1077
rect 499393 1068 499405 1071
rect 483799 1040 499405 1068
rect 483799 1037 483811 1040
rect 483753 1031 483811 1037
rect 499393 1037 499405 1040
rect 499439 1037 499451 1071
rect 499393 1031 499451 1037
rect 502337 1071 502395 1077
rect 502337 1037 502349 1071
rect 502383 1068 502395 1071
rect 509697 1071 509755 1077
rect 509697 1068 509709 1071
rect 502383 1040 509709 1068
rect 502383 1037 502395 1040
rect 502337 1031 502395 1037
rect 509697 1037 509709 1040
rect 509743 1037 509755 1071
rect 509697 1031 509755 1037
rect 517057 1071 517115 1077
rect 517057 1037 517069 1071
rect 517103 1068 517115 1071
rect 533709 1071 533767 1077
rect 533709 1068 533721 1071
rect 517103 1040 533721 1068
rect 517103 1037 517115 1040
rect 517057 1031 517115 1037
rect 533709 1037 533721 1040
rect 533755 1037 533767 1071
rect 533709 1031 533767 1037
rect 555789 1071 555847 1077
rect 555789 1037 555801 1071
rect 555835 1068 555847 1071
rect 563514 1068 563520 1080
rect 555835 1040 563520 1068
rect 555835 1037 555847 1040
rect 555789 1031 555847 1037
rect 563514 1028 563520 1040
rect 563572 1028 563578 1080
rect 487709 1003 487767 1009
rect 487709 1000 487721 1003
rect 483676 972 487721 1000
rect 482833 963 482891 969
rect 487709 969 487721 972
rect 487755 969 487767 1003
rect 507305 1003 507363 1009
rect 507305 1000 507317 1003
rect 487709 963 487767 969
rect 493428 972 507317 1000
rect 481453 935 481511 941
rect 465736 904 466454 932
rect 461765 895 461823 901
rect 432509 827 432567 833
rect 432616 836 437474 864
rect 439869 867 439927 873
rect 418801 799 418859 805
rect 418801 765 418813 799
rect 418847 796 418859 799
rect 423769 799 423827 805
rect 423769 796 423781 799
rect 418847 768 423781 796
rect 418847 765 418859 768
rect 418801 759 418859 765
rect 423769 765 423781 768
rect 423815 765 423827 799
rect 423769 759 423827 765
rect 424689 799 424747 805
rect 424689 765 424701 799
rect 424735 796 424747 799
rect 432616 796 432644 836
rect 439869 833 439881 867
rect 439915 864 439927 867
rect 452381 867 452439 873
rect 439915 836 444374 864
rect 439915 833 439927 836
rect 439869 827 439927 833
rect 443641 799 443699 805
rect 443641 796 443653 799
rect 424735 768 432644 796
rect 435192 768 443653 796
rect 424735 765 424747 768
rect 424689 759 424747 765
rect 422849 731 422907 737
rect 422849 697 422861 731
rect 422895 728 422907 731
rect 422895 700 435128 728
rect 422895 697 422907 700
rect 422849 691 422907 697
rect 415486 660 415492 672
rect 415412 632 415492 660
rect 415486 620 415492 632
rect 415544 620 415550 672
rect 416682 620 416688 672
rect 416740 620 416746 672
rect 417142 660 417148 672
rect 417103 632 417148 660
rect 417142 620 417148 632
rect 417200 620 417206 672
rect 418338 620 418344 672
rect 418396 660 418402 672
rect 430850 660 430856 672
rect 418396 632 430856 660
rect 418396 620 418402 632
rect 430850 620 430856 632
rect 430908 620 430914 672
rect 432509 663 432567 669
rect 432509 629 432521 663
rect 432555 660 432567 663
rect 434438 660 434444 672
rect 432555 632 434444 660
rect 432555 629 432567 632
rect 432509 623 432567 629
rect 434438 620 434444 632
rect 434496 620 434502 672
rect 419902 592 419908 604
rect 413204 564 419908 592
rect 419902 552 419908 564
rect 419960 552 419966 604
rect 421650 592 421656 604
rect 421611 564 421656 592
rect 421650 552 421656 564
rect 421708 552 421714 604
rect 422846 592 422852 604
rect 422807 564 422852 592
rect 422846 552 422852 564
rect 422904 552 422910 604
rect 423766 592 423772 604
rect 423727 564 423772 592
rect 423766 552 423772 564
rect 423824 552 423830 604
rect 424686 592 424692 604
rect 424647 564 424692 592
rect 424686 552 424692 564
rect 424744 552 424750 604
rect 424962 552 424968 604
rect 425020 552 425026 604
rect 433242 592 433248 604
rect 429166 564 433248 592
rect 413112 524 413140 552
rect 404648 496 413140 524
rect 414934 484 414940 536
rect 414992 524 414998 536
rect 421742 524 421748 536
rect 414992 496 421748 524
rect 414992 484 414998 496
rect 421742 484 421748 496
rect 421800 484 421806 536
rect 424502 484 424508 536
rect 424560 524 424566 536
rect 424980 524 425008 552
rect 426342 524 426348 536
rect 424560 496 425008 524
rect 426303 496 426348 524
rect 424560 484 424566 496
rect 426342 484 426348 496
rect 426400 484 426406 536
rect 429010 524 429016 536
rect 428971 496 429016 524
rect 429010 484 429016 496
rect 429068 484 429074 536
rect 366784 428 367094 456
rect 366784 416 366790 428
rect 367830 416 367836 468
rect 367888 456 367894 468
rect 375650 456 375656 468
rect 367888 428 375656 456
rect 367888 416 367894 428
rect 375650 416 375656 428
rect 375708 416 375714 468
rect 378410 416 378416 468
rect 378468 456 378474 468
rect 389453 459 389511 465
rect 389453 456 389465 459
rect 378468 428 389465 456
rect 378468 416 378474 428
rect 389453 425 389465 428
rect 389499 425 389511 459
rect 406194 456 406200 468
rect 389453 419 389511 425
rect 397840 428 406200 456
rect 364797 391 364855 397
rect 364797 357 364809 391
rect 364843 388 364855 391
rect 365990 388 365996 400
rect 364843 360 365996 388
rect 364843 357 364855 360
rect 364797 351 364855 357
rect 365990 348 365996 360
rect 366048 348 366054 400
rect 376294 348 376300 400
rect 376352 388 376358 400
rect 386966 388 386972 400
rect 376352 360 386972 388
rect 376352 348 376358 360
rect 386966 348 386972 360
rect 387024 348 387030 400
rect 388806 348 388812 400
rect 388864 388 388870 400
rect 390189 391 390247 397
rect 390189 388 390201 391
rect 388864 360 390201 388
rect 388864 348 388870 360
rect 390189 357 390201 360
rect 390235 357 390247 391
rect 390189 351 390247 357
rect 391014 348 391020 400
rect 391072 388 391078 400
rect 396169 391 396227 397
rect 391072 360 396074 388
rect 391072 348 391078 360
rect 363690 320 363696 332
rect 354732 292 356054 320
rect 358786 292 363696 320
rect 354732 280 354738 292
rect 255682 212 255688 264
rect 255740 252 255746 264
rect 261938 252 261944 264
rect 255740 224 261944 252
rect 255740 212 255746 224
rect 261938 212 261944 224
rect 261996 212 262002 264
rect 264882 212 264888 264
rect 264940 252 264946 264
rect 271046 252 271052 264
rect 264940 224 271052 252
rect 264940 212 264946 224
rect 271046 212 271052 224
rect 271104 212 271110 264
rect 274082 212 274088 264
rect 274140 252 274146 264
rect 280709 255 280767 261
rect 280709 252 280721 255
rect 274140 224 280721 252
rect 274140 212 274146 224
rect 280709 221 280721 224
rect 280755 221 280767 255
rect 280709 215 280767 221
rect 289814 212 289820 264
rect 289872 252 289878 264
rect 296990 252 296996 264
rect 289872 224 296996 252
rect 289872 212 289878 224
rect 296990 212 296996 224
rect 297048 212 297054 264
rect 297910 212 297916 264
rect 297968 252 297974 264
rect 305730 252 305736 264
rect 297968 224 305736 252
rect 297968 212 297974 224
rect 305730 212 305736 224
rect 305788 212 305794 264
rect 308766 212 308772 264
rect 308824 252 308830 264
rect 316586 252 316592 264
rect 308824 224 316592 252
rect 308824 212 308830 224
rect 316586 212 316592 224
rect 316644 212 316650 264
rect 326338 212 326344 264
rect 326396 252 326402 264
rect 335354 252 335360 264
rect 326396 224 335360 252
rect 326396 212 326402 224
rect 335354 212 335360 224
rect 335412 212 335418 264
rect 345566 212 345572 264
rect 345624 252 345630 264
rect 355229 255 355287 261
rect 355229 252 355241 255
rect 345624 224 355241 252
rect 345624 212 345630 224
rect 355229 221 355241 224
rect 355275 221 355287 255
rect 356026 252 356054 292
rect 363690 280 363696 292
rect 363748 280 363754 332
rect 364886 280 364892 332
rect 364944 320 364950 332
rect 372065 323 372123 329
rect 372065 320 372077 323
rect 364944 292 372077 320
rect 364944 280 364950 292
rect 372065 289 372077 292
rect 372111 289 372123 323
rect 372065 283 372123 289
rect 381998 280 382004 332
rect 382056 320 382062 332
rect 393222 320 393228 332
rect 382056 292 393228 320
rect 382056 280 382062 292
rect 393222 280 393228 292
rect 393280 280 393286 332
rect 396046 320 396074 360
rect 396169 357 396181 391
rect 396215 388 396227 391
rect 397840 388 397868 428
rect 406194 416 406200 428
rect 406252 416 406258 468
rect 408126 416 408132 468
rect 408184 456 408190 468
rect 411441 459 411499 465
rect 411441 456 411453 459
rect 408184 428 411453 456
rect 408184 416 408190 428
rect 411441 425 411453 428
rect 411487 425 411499 459
rect 411441 419 411499 425
rect 411530 416 411536 468
rect 411588 456 411594 468
rect 418801 459 418859 465
rect 418801 456 418813 459
rect 411588 428 418813 456
rect 411588 416 411594 428
rect 418801 425 418813 428
rect 418847 425 418859 459
rect 418801 419 418859 425
rect 420546 416 420552 468
rect 420604 456 420610 468
rect 429166 456 429194 564
rect 433242 552 433248 564
rect 433300 552 433306 604
rect 435100 592 435128 700
rect 435192 672 435220 768
rect 443641 765 443653 768
rect 443687 765 443699 799
rect 444346 796 444374 836
rect 452381 833 452393 867
rect 452427 864 452439 867
rect 452427 836 466224 864
rect 452427 833 452439 836
rect 452381 827 452439 833
rect 453485 799 453543 805
rect 453485 796 453497 799
rect 444346 768 453497 796
rect 443641 759 443699 765
rect 453485 765 453497 768
rect 453531 765 453543 799
rect 453485 759 453543 765
rect 454681 799 454739 805
rect 454681 765 454693 799
rect 454727 796 454739 799
rect 458177 799 458235 805
rect 458177 796 458189 799
rect 454727 768 458189 796
rect 454727 765 454739 768
rect 454681 759 454739 765
rect 458177 765 458189 768
rect 458223 765 458235 799
rect 458177 759 458235 765
rect 459526 768 460934 796
rect 449989 731 450047 737
rect 449989 728 450001 731
rect 437446 700 450001 728
rect 435174 620 435180 672
rect 435232 620 435238 672
rect 436462 620 436468 672
rect 436520 660 436526 672
rect 437446 660 437474 700
rect 449989 697 450001 700
rect 450035 697 450047 731
rect 449989 691 450047 697
rect 451277 731 451335 737
rect 451277 697 451289 731
rect 451323 728 451335 731
rect 459526 728 459554 768
rect 451323 700 459554 728
rect 451323 697 451335 700
rect 451277 691 451335 697
rect 437934 660 437940 672
rect 436520 632 437474 660
rect 437895 632 437940 660
rect 436520 620 436526 632
rect 437934 620 437940 632
rect 437992 620 437998 672
rect 442626 660 442632 672
rect 439056 632 442632 660
rect 435542 592 435548 604
rect 435100 564 435548 592
rect 435542 552 435548 564
rect 435600 552 435606 604
rect 439056 592 439084 632
rect 442626 620 442632 632
rect 442684 620 442690 672
rect 443641 663 443699 669
rect 443641 629 443653 663
rect 443687 660 443699 663
rect 448238 660 448244 672
rect 443687 632 448244 660
rect 443687 629 443699 632
rect 443641 623 443699 629
rect 448238 620 448244 632
rect 448296 620 448302 672
rect 448974 660 448980 672
rect 448935 632 448980 660
rect 448974 620 448980 632
rect 449032 620 449038 672
rect 454681 663 454739 669
rect 454681 660 454693 663
rect 449866 632 454693 660
rect 441522 592 441528 604
rect 435652 564 439084 592
rect 439148 564 441528 592
rect 429470 484 429476 536
rect 429528 524 429534 536
rect 435652 524 435680 564
rect 429528 496 435680 524
rect 435729 527 435787 533
rect 429528 484 429534 496
rect 435729 493 435741 527
rect 435775 524 435787 527
rect 439148 524 439176 564
rect 441522 552 441528 564
rect 441580 552 441586 604
rect 442166 592 442172 604
rect 442127 564 442172 592
rect 442166 552 442172 564
rect 442224 552 442230 604
rect 443822 592 443828 604
rect 443783 564 443828 592
rect 443822 552 443828 564
rect 443880 552 443886 604
rect 444466 552 444472 604
rect 444524 592 444530 604
rect 449866 592 449894 632
rect 454681 629 454693 632
rect 454727 629 454739 663
rect 454681 623 454739 629
rect 454773 663 454831 669
rect 454773 629 454785 663
rect 454819 660 454831 663
rect 456886 660 456892 672
rect 454819 632 456892 660
rect 454819 629 454831 632
rect 454773 623 454831 629
rect 456886 620 456892 632
rect 456944 620 456950 672
rect 457990 660 457996 672
rect 457951 632 457996 660
rect 457990 620 457996 632
rect 458048 620 458054 672
rect 458174 620 458180 672
rect 458232 660 458238 672
rect 460198 660 460204 672
rect 458232 632 458277 660
rect 460159 632 460204 660
rect 458232 620 458238 632
rect 460198 620 460204 632
rect 460256 620 460262 672
rect 444524 564 449894 592
rect 444524 552 444530 564
rect 449986 552 449992 604
rect 450044 592 450050 604
rect 451274 592 451280 604
rect 450044 564 450089 592
rect 451235 564 451280 592
rect 450044 552 450050 564
rect 451274 552 451280 564
rect 451332 552 451338 604
rect 452378 592 452384 604
rect 452339 564 452384 592
rect 452378 552 452384 564
rect 452436 552 452442 604
rect 454494 592 454500 604
rect 454455 564 454500 592
rect 454494 552 454500 564
rect 454552 552 454558 604
rect 455325 595 455383 601
rect 455325 561 455337 595
rect 455371 592 455383 595
rect 455690 592 455696 604
rect 455371 564 455696 592
rect 455371 561 455383 564
rect 455325 555 455383 561
rect 455690 552 455696 564
rect 455748 552 455754 604
rect 455877 595 455935 601
rect 455877 561 455889 595
rect 455923 592 455935 595
rect 459186 592 459192 604
rect 455923 564 459192 592
rect 455923 561 455935 564
rect 455877 555 455935 561
rect 459186 552 459192 564
rect 459244 552 459250 604
rect 460906 592 460934 768
rect 461949 731 462007 737
rect 461949 697 461961 731
rect 461995 728 462007 731
rect 461995 700 466132 728
rect 461995 697 462007 700
rect 461949 691 462007 697
rect 462225 663 462283 669
rect 462225 629 462237 663
rect 462271 660 462283 663
rect 462774 660 462780 672
rect 462271 632 462780 660
rect 462271 629 462283 632
rect 462225 623 462283 629
rect 462774 620 462780 632
rect 462832 620 462838 672
rect 465166 592 465172 604
rect 460906 564 465172 592
rect 465166 552 465172 564
rect 465224 552 465230 604
rect 466104 592 466132 700
rect 466196 660 466224 836
rect 466270 660 466276 672
rect 466196 632 466276 660
rect 466270 620 466276 632
rect 466328 620 466334 672
rect 466426 660 466454 904
rect 481453 901 481465 935
rect 481499 932 481511 935
rect 481499 904 493364 932
rect 481499 901 481511 904
rect 481453 895 481511 901
rect 486421 867 486479 873
rect 486421 864 486433 867
rect 473326 836 486433 864
rect 469585 731 469643 737
rect 469585 697 469597 731
rect 469631 728 469643 731
rect 473326 728 473354 836
rect 486421 833 486433 836
rect 486467 833 486479 867
rect 486421 827 486479 833
rect 475105 799 475163 805
rect 475105 765 475117 799
rect 475151 796 475163 799
rect 475151 768 489960 796
rect 475151 765 475163 768
rect 475105 759 475163 765
rect 489825 731 489883 737
rect 489825 728 489837 731
rect 469631 700 471284 728
rect 469631 697 469643 700
rect 469585 691 469643 697
rect 471054 660 471060 672
rect 466426 632 471060 660
rect 471054 620 471060 632
rect 471112 620 471118 672
rect 469858 592 469864 604
rect 466104 564 469864 592
rect 469858 552 469864 564
rect 469916 552 469922 604
rect 471256 592 471284 700
rect 471716 700 473354 728
rect 481606 700 489837 728
rect 471716 672 471744 700
rect 471698 620 471704 672
rect 471756 620 471762 672
rect 472250 660 472256 672
rect 472211 632 472256 660
rect 472250 620 472256 632
rect 472308 620 472314 672
rect 472802 660 472808 672
rect 472763 632 472808 660
rect 472802 620 472808 632
rect 472860 620 472866 672
rect 474550 660 474556 672
rect 474511 632 474556 660
rect 474550 620 474556 632
rect 474608 620 474614 672
rect 474921 663 474979 669
rect 474921 629 474933 663
rect 474967 660 474979 663
rect 480714 660 480720 672
rect 474967 632 480720 660
rect 474967 629 474979 632
rect 474921 623 474979 629
rect 480714 620 480720 632
rect 480772 620 480778 672
rect 481450 660 481456 672
rect 481411 632 481456 660
rect 481450 620 481456 632
rect 481508 620 481514 672
rect 475102 592 475108 604
rect 471256 564 474734 592
rect 475063 564 475108 592
rect 435775 496 439176 524
rect 435775 493 435787 496
rect 435729 487 435787 493
rect 443270 484 443276 536
rect 443328 524 443334 536
rect 453482 524 453488 536
rect 443328 496 449894 524
rect 453443 496 453488 524
rect 443328 484 443334 496
rect 430390 456 430396 468
rect 420604 428 429194 456
rect 430351 428 430396 456
rect 420604 416 420610 428
rect 430390 416 430396 428
rect 430448 416 430454 468
rect 434254 416 434260 468
rect 434312 456 434318 468
rect 447134 456 447140 468
rect 434312 428 447140 456
rect 434312 416 434318 428
rect 447134 416 447140 428
rect 447192 416 447198 468
rect 449866 456 449894 496
rect 453482 484 453488 496
rect 453540 484 453546 536
rect 453574 484 453580 536
rect 453632 524 453638 536
rect 466086 524 466092 536
rect 453632 496 466092 524
rect 453632 484 453638 496
rect 466086 484 466092 496
rect 466144 484 466150 536
rect 467190 484 467196 536
rect 467248 524 467254 536
rect 469769 527 469827 533
rect 469769 524 469781 527
rect 467248 496 469781 524
rect 467248 484 467254 496
rect 469769 493 469781 496
rect 469815 493 469827 527
rect 474706 524 474734 564
rect 475102 552 475108 564
rect 475160 552 475166 604
rect 476206 592 476212 604
rect 476167 564 476212 592
rect 476206 552 476212 564
rect 476264 552 476270 604
rect 476574 592 476580 604
rect 476535 564 476580 592
rect 476574 552 476580 564
rect 476632 552 476638 604
rect 477862 592 477868 604
rect 477236 564 477868 592
rect 477236 524 477264 564
rect 477862 552 477868 564
rect 477920 552 477926 604
rect 480622 552 480628 604
rect 480680 592 480686 604
rect 481606 592 481634 700
rect 489825 697 489837 700
rect 489871 697 489883 731
rect 489825 691 489883 697
rect 489932 672 489960 768
rect 490009 731 490067 737
rect 490009 697 490021 731
rect 490055 728 490067 731
rect 490055 700 491340 728
rect 490055 697 490067 700
rect 490009 691 490067 697
rect 491312 672 491340 700
rect 493336 672 493364 904
rect 483750 660 483756 672
rect 483711 632 483756 660
rect 483750 620 483756 632
rect 483808 620 483814 672
rect 485222 660 485228 672
rect 483952 632 485228 660
rect 481726 592 481732 604
rect 480680 564 481634 592
rect 481687 564 481732 592
rect 480680 552 480686 564
rect 481726 552 481732 564
rect 481784 552 481790 604
rect 474706 496 477264 524
rect 469769 487 469827 493
rect 477402 484 477408 536
rect 477460 524 477466 536
rect 483952 524 483980 632
rect 485222 620 485228 632
rect 485280 620 485286 672
rect 487706 660 487712 672
rect 487667 632 487712 660
rect 487706 620 487712 632
rect 487764 620 487770 672
rect 489914 620 489920 672
rect 489972 620 489978 672
rect 491110 660 491116 672
rect 491071 632 491116 660
rect 491110 620 491116 632
rect 491168 620 491174 672
rect 491294 620 491300 672
rect 491352 620 491358 672
rect 493229 663 493287 669
rect 493229 660 493241 663
rect 491404 632 493241 660
rect 484026 552 484032 604
rect 484084 552 484090 604
rect 486418 592 486424 604
rect 486379 564 486424 592
rect 486418 552 486424 564
rect 486476 552 486482 604
rect 487430 552 487436 604
rect 487488 592 487494 604
rect 491404 592 491432 632
rect 493229 629 493241 632
rect 493275 629 493287 663
rect 493229 623 493287 629
rect 493318 620 493324 672
rect 493376 620 493382 672
rect 487488 564 491432 592
rect 487488 552 487494 564
rect 492122 552 492128 604
rect 492180 592 492186 604
rect 493428 592 493456 972
rect 507305 969 507317 972
rect 507351 969 507363 1003
rect 507305 963 507363 969
rect 509237 1003 509295 1009
rect 509237 969 509249 1003
rect 509283 1000 509295 1003
rect 525153 1003 525211 1009
rect 525153 1000 525165 1003
rect 509283 972 525165 1000
rect 509283 969 509295 972
rect 509237 963 509295 969
rect 525153 969 525165 972
rect 525199 969 525211 1003
rect 525153 963 525211 969
rect 558733 1003 558791 1009
rect 558733 969 558745 1003
rect 558779 1000 558791 1003
rect 569862 1000 569868 1012
rect 558779 972 569868 1000
rect 558779 969 558791 972
rect 558733 963 558791 969
rect 569862 960 569868 972
rect 569920 960 569926 1012
rect 505741 935 505799 941
rect 505741 901 505753 935
rect 505787 932 505799 935
rect 521841 935 521899 941
rect 521841 932 521853 935
rect 505787 904 521853 932
rect 505787 901 505799 904
rect 505741 895 505799 901
rect 521841 901 521853 904
rect 521887 901 521899 935
rect 521841 895 521899 901
rect 531869 935 531927 941
rect 531869 901 531881 935
rect 531915 932 531927 935
rect 549073 935 549131 941
rect 549073 932 549085 935
rect 531915 904 549085 932
rect 531915 901 531927 904
rect 531869 895 531927 901
rect 549073 901 549085 904
rect 549119 901 549131 935
rect 549073 895 549131 901
rect 562597 935 562655 941
rect 562597 901 562609 935
rect 562643 932 562655 935
rect 575474 932 575480 944
rect 562643 904 575480 932
rect 562643 901 562655 904
rect 562597 895 562655 901
rect 575474 892 575480 904
rect 575532 892 575538 944
rect 513285 867 513343 873
rect 513285 833 513297 867
rect 513331 864 513343 867
rect 530121 867 530179 873
rect 530121 864 530133 867
rect 513331 836 530133 864
rect 513331 833 513343 836
rect 513285 827 513343 833
rect 530121 833 530133 836
rect 530167 833 530179 867
rect 530121 827 530179 833
rect 536469 867 536527 873
rect 536469 833 536481 867
rect 536515 864 536527 867
rect 548889 867 548947 873
rect 536515 836 546494 864
rect 536515 833 536527 836
rect 536469 827 536527 833
rect 515861 799 515919 805
rect 515861 765 515873 799
rect 515907 796 515919 799
rect 524141 799 524199 805
rect 524141 796 524153 799
rect 515907 768 524153 796
rect 515907 765 515919 768
rect 515861 759 515919 765
rect 524141 765 524153 768
rect 524187 765 524199 799
rect 540793 799 540851 805
rect 540793 796 540805 799
rect 524141 759 524199 765
rect 524386 768 540805 796
rect 524386 728 524414 768
rect 540793 765 540805 768
rect 540839 765 540851 799
rect 540793 759 540851 765
rect 492180 564 493456 592
rect 493520 700 506520 728
rect 492180 552 492186 564
rect 477460 496 483980 524
rect 477460 484 477466 496
rect 454773 459 454831 465
rect 454773 456 454785 459
rect 449866 428 454785 456
rect 454773 425 454785 428
rect 454819 425 454831 459
rect 454773 419 454831 425
rect 455322 416 455328 468
rect 455380 456 455386 468
rect 455417 459 455475 465
rect 455417 456 455429 459
rect 455380 428 455429 456
rect 455380 416 455386 428
rect 455417 425 455429 428
rect 455463 425 455475 459
rect 456518 456 456524 468
rect 456479 428 456524 456
rect 455417 419 455475 425
rect 456518 416 456524 428
rect 456576 416 456582 468
rect 468478 456 468484 468
rect 459526 428 468484 456
rect 396215 360 397868 388
rect 396215 357 396227 360
rect 396169 351 396227 357
rect 399938 348 399944 400
rect 399996 388 400002 400
rect 411714 388 411720 400
rect 399996 360 411720 388
rect 399996 348 400002 360
rect 411714 348 411720 360
rect 411772 348 411778 400
rect 416038 348 416044 400
rect 416096 388 416102 400
rect 428642 388 428648 400
rect 416096 360 428648 388
rect 416096 348 416102 360
rect 428642 348 428648 360
rect 428700 348 428706 400
rect 436462 388 436468 400
rect 432248 360 436468 388
rect 402238 320 402244 332
rect 396046 292 402244 320
rect 402238 280 402244 292
rect 402296 280 402302 332
rect 403434 280 403440 332
rect 403492 320 403498 332
rect 406473 323 406531 329
rect 406473 320 406485 323
rect 403492 292 406485 320
rect 403492 280 403498 292
rect 406473 289 406485 292
rect 406519 289 406531 323
rect 406473 283 406531 289
rect 409230 280 409236 332
rect 409288 320 409294 332
rect 421006 320 421012 332
rect 409288 292 421012 320
rect 409288 280 409294 292
rect 421006 280 421012 292
rect 421064 280 421070 332
rect 423490 280 423496 332
rect 423548 320 423554 332
rect 432248 320 432276 360
rect 436462 348 436468 360
rect 436520 348 436526 400
rect 437474 348 437480 400
rect 437532 388 437538 400
rect 450630 388 450636 400
rect 437532 360 450636 388
rect 437532 348 437538 360
rect 450630 348 450636 360
rect 450688 348 450694 400
rect 452286 388 452292 400
rect 450970 360 452292 388
rect 423548 292 432276 320
rect 423548 280 423554 292
rect 433058 280 433064 332
rect 433116 320 433122 332
rect 446030 320 446036 332
rect 433116 292 446036 320
rect 433116 280 433122 292
rect 446030 280 446036 292
rect 446088 280 446094 332
rect 450970 320 450998 360
rect 452286 348 452292 360
rect 452344 348 452350 400
rect 454218 348 454224 400
rect 454276 388 454282 400
rect 459526 388 459554 428
rect 468478 416 468484 428
rect 468536 416 468542 468
rect 469214 416 469220 468
rect 469272 456 469278 468
rect 484044 456 484072 552
rect 489730 484 489736 536
rect 489788 524 489794 536
rect 493413 527 493471 533
rect 493413 524 493425 527
rect 489788 496 493425 524
rect 489788 484 489794 496
rect 493413 493 493425 496
rect 493459 493 493471 527
rect 493413 487 493471 493
rect 469272 428 484072 456
rect 469272 416 469278 428
rect 490926 416 490932 468
rect 490984 456 490990 468
rect 493520 456 493548 700
rect 506492 672 506520 700
rect 507826 700 523080 728
rect 494422 660 494428 672
rect 494383 632 494428 660
rect 494422 620 494428 632
rect 494480 620 494486 672
rect 502978 660 502984 672
rect 494532 632 502984 660
rect 493597 595 493655 601
rect 493597 561 493609 595
rect 493643 592 493655 595
rect 494532 592 494560 632
rect 502978 620 502984 632
rect 503036 620 503042 672
rect 505738 660 505744 672
rect 505699 632 505744 660
rect 505738 620 505744 632
rect 505796 620 505802 672
rect 506474 620 506480 672
rect 506532 620 506538 672
rect 506934 620 506940 672
rect 506992 660 506998 672
rect 507826 660 507854 700
rect 523052 672 523080 700
rect 523972 700 524414 728
rect 525061 731 525119 737
rect 523972 672 524000 700
rect 525061 697 525073 731
rect 525107 728 525119 731
rect 525107 700 542216 728
rect 525107 697 525119 700
rect 525061 691 525119 697
rect 542188 672 542216 700
rect 509234 660 509240 672
rect 506992 632 507854 660
rect 509195 632 509240 660
rect 506992 620 506998 632
rect 509234 620 509240 632
rect 509292 620 509298 672
rect 509694 660 509700 672
rect 509655 632 509700 660
rect 509694 620 509700 632
rect 509752 620 509758 672
rect 511258 660 511264 672
rect 511219 632 511264 660
rect 511258 620 511264 632
rect 511316 620 511322 672
rect 512454 660 512460 672
rect 512415 632 512460 660
rect 512454 620 512460 632
rect 512512 620 512518 672
rect 513282 660 513288 672
rect 513243 632 513288 660
rect 513282 620 513288 632
rect 513340 620 513346 672
rect 515858 660 515864 672
rect 515819 632 515864 660
rect 515858 620 515864 632
rect 515916 620 515922 672
rect 517054 660 517060 672
rect 517015 632 517060 660
rect 517054 620 517060 632
rect 517112 620 517118 672
rect 519354 660 519360 672
rect 519315 632 519360 660
rect 519354 620 519360 632
rect 519412 620 519418 672
rect 521838 660 521844 672
rect 521799 632 521844 660
rect 521838 620 521844 632
rect 521896 620 521902 672
rect 523034 620 523040 672
rect 523092 620 523098 672
rect 523954 620 523960 672
rect 524012 620 524018 672
rect 528833 663 528891 669
rect 528833 660 528845 663
rect 524064 632 528845 660
rect 495342 592 495348 604
rect 493643 564 494560 592
rect 495303 564 495348 592
rect 493643 561 493655 564
rect 493597 555 493655 561
rect 495342 552 495348 564
rect 495400 552 495406 604
rect 496722 592 496728 604
rect 496683 564 496728 592
rect 496722 552 496728 564
rect 496780 552 496786 604
rect 498194 552 498200 604
rect 498252 592 498258 604
rect 499390 592 499396 604
rect 498252 564 498297 592
rect 499351 564 499396 592
rect 498252 552 498258 564
rect 499390 552 499396 564
rect 499448 552 499454 604
rect 500126 552 500132 604
rect 500184 592 500190 604
rect 516134 592 516140 604
rect 500184 564 516140 592
rect 500184 552 500190 564
rect 516134 552 516140 564
rect 516192 552 516198 604
rect 518158 552 518164 604
rect 518216 592 518222 604
rect 524064 592 524092 632
rect 528833 629 528845 632
rect 528879 629 528891 663
rect 532510 660 532516 672
rect 528833 623 528891 629
rect 528940 632 532516 660
rect 518216 564 524092 592
rect 524141 595 524199 601
rect 518216 552 518222 564
rect 524141 561 524153 595
rect 524187 592 524199 595
rect 528940 592 528968 632
rect 532510 620 532516 632
rect 532568 620 532574 672
rect 533062 620 533068 672
rect 533120 660 533126 672
rect 535822 660 535828 672
rect 533120 632 534856 660
rect 535783 632 535828 660
rect 533120 620 533126 632
rect 524187 564 528968 592
rect 524187 561 524199 564
rect 524141 555 524199 561
rect 529014 552 529020 604
rect 529072 552 529078 604
rect 530118 592 530124 604
rect 530079 564 530124 592
rect 530118 552 530124 564
rect 530176 552 530182 604
rect 531866 592 531872 604
rect 531827 564 531872 592
rect 531866 552 531872 564
rect 531924 552 531930 604
rect 533706 592 533712 604
rect 533667 564 533712 592
rect 533706 552 533712 564
rect 533764 552 533770 604
rect 534828 592 534856 632
rect 535822 620 535828 632
rect 535880 620 535886 672
rect 536466 660 536472 672
rect 536427 632 536472 660
rect 536466 620 536472 632
rect 536524 620 536530 672
rect 540790 660 540796 672
rect 540751 632 540796 660
rect 540790 620 540796 632
rect 540848 620 540854 672
rect 542170 620 542176 672
rect 542228 620 542234 672
rect 543182 660 543188 672
rect 543143 632 543188 660
rect 543182 620 543188 632
rect 543240 620 543246 672
rect 545482 660 545488 672
rect 545443 632 545488 660
rect 545482 620 545488 632
rect 545540 620 545546 672
rect 546466 660 546494 836
rect 548889 833 548901 867
rect 548935 864 548947 867
rect 562229 867 562287 873
rect 562229 864 562241 867
rect 548935 836 562241 864
rect 548935 833 548947 836
rect 548889 827 548947 833
rect 562229 833 562241 836
rect 562275 833 562287 867
rect 565906 864 565912 876
rect 562229 827 562287 833
rect 562336 836 565912 864
rect 551189 799 551247 805
rect 551189 765 551201 799
rect 551235 796 551247 799
rect 562336 796 562364 836
rect 565906 824 565912 836
rect 565964 824 565970 876
rect 551235 768 562364 796
rect 551235 765 551247 768
rect 551189 759 551247 765
rect 565814 756 565820 808
rect 565872 796 565878 808
rect 568022 796 568028 808
rect 565872 768 568028 796
rect 565872 756 565878 768
rect 568022 756 568028 768
rect 568080 756 568086 808
rect 548521 731 548579 737
rect 548521 697 548533 731
rect 548567 728 548579 731
rect 570322 728 570328 740
rect 548567 700 555188 728
rect 548567 697 548579 700
rect 548521 691 548579 697
rect 555160 672 555188 700
rect 556632 700 570328 728
rect 553762 660 553768 672
rect 546466 632 553768 660
rect 553762 620 553768 632
rect 553820 620 553826 672
rect 555142 620 555148 672
rect 555200 620 555206 672
rect 555786 660 555792 672
rect 555747 632 555792 660
rect 555786 620 555792 632
rect 555844 620 555850 672
rect 550266 592 550272 604
rect 534828 564 550272 592
rect 550266 552 550272 564
rect 550324 552 550330 604
rect 551186 592 551192 604
rect 551147 564 551192 592
rect 551186 552 551192 564
rect 551244 552 551250 604
rect 552382 552 552388 604
rect 552440 592 552446 604
rect 556632 592 556660 700
rect 570322 688 570328 700
rect 570380 688 570386 740
rect 556890 620 556896 672
rect 556948 660 556954 672
rect 575106 660 575112 672
rect 556948 632 575112 660
rect 556948 620 556954 632
rect 575106 620 575112 632
rect 575164 620 575170 672
rect 565814 592 565820 604
rect 552440 564 556660 592
rect 557506 564 565820 592
rect 552440 552 552446 564
rect 493689 527 493747 533
rect 493689 493 493701 527
rect 493735 524 493747 527
rect 505094 524 505100 536
rect 493735 496 505100 524
rect 493735 493 493747 496
rect 493689 487 493747 493
rect 505094 484 505100 496
rect 505152 484 505158 536
rect 507302 524 507308 536
rect 507263 496 507308 524
rect 507302 484 507308 496
rect 507360 484 507366 536
rect 512178 484 512184 536
rect 512236 524 512242 536
rect 529032 524 529060 552
rect 512236 496 529060 524
rect 512236 484 512242 496
rect 529658 484 529664 536
rect 529716 524 529722 536
rect 529716 496 536834 524
rect 529716 484 529722 496
rect 502334 456 502340 468
rect 490984 428 493548 456
rect 502295 428 502340 456
rect 490984 416 490990 428
rect 502334 416 502340 428
rect 502392 416 502398 468
rect 503530 416 503536 468
rect 503588 456 503594 468
rect 519722 456 519728 468
rect 503588 428 519728 456
rect 503588 416 503594 428
rect 519722 416 519728 428
rect 519780 416 519786 468
rect 525058 456 525064 468
rect 525019 428 525064 456
rect 525058 416 525064 428
rect 525116 416 525122 468
rect 525150 416 525156 468
rect 525208 456 525214 468
rect 528833 459 528891 465
rect 525208 428 525253 456
rect 525208 416 525214 428
rect 528833 425 528845 459
rect 528879 456 528891 459
rect 534534 456 534540 468
rect 528879 428 534540 456
rect 528879 425 528891 428
rect 528833 419 528891 425
rect 534534 416 534540 428
rect 534592 416 534598 468
rect 536806 456 536834 496
rect 538766 484 538772 536
rect 538824 524 538830 536
rect 548521 527 548579 533
rect 548521 524 548533 527
rect 538824 496 548533 524
rect 538824 484 538830 496
rect 548521 493 548533 496
rect 548567 493 548579 527
rect 548886 524 548892 536
rect 548847 496 548892 524
rect 548521 487 548579 493
rect 548886 484 548892 496
rect 548944 484 548950 536
rect 549073 527 549131 533
rect 549073 493 549085 527
rect 549119 524 549131 527
rect 549254 524 549260 536
rect 549119 496 549260 524
rect 549119 493 549131 496
rect 549073 487 549131 493
rect 549254 484 549260 496
rect 549312 484 549318 536
rect 550082 484 550088 536
rect 550140 524 550146 536
rect 557506 524 557534 564
rect 565814 552 565820 564
rect 565872 552 565878 604
rect 578602 552 578608 604
rect 578660 552 578666 604
rect 557994 524 558000 536
rect 550140 496 557534 524
rect 557955 496 558000 524
rect 550140 484 550146 496
rect 557994 484 558000 496
rect 558052 484 558058 536
rect 558730 524 558736 536
rect 558691 496 558736 524
rect 558730 484 558736 496
rect 558788 484 558794 536
rect 560202 484 560208 536
rect 560260 524 560266 536
rect 578620 524 578648 552
rect 560260 496 578648 524
rect 560260 484 560266 496
rect 546494 456 546500 468
rect 536806 428 546500 456
rect 546494 416 546500 428
rect 546552 416 546558 468
rect 547690 416 547696 468
rect 547748 456 547754 468
rect 562594 456 562600 468
rect 547748 428 561904 456
rect 562555 428 562600 456
rect 547748 416 547754 428
rect 454276 360 459554 388
rect 454276 348 454282 360
rect 465994 348 466000 400
rect 466052 388 466058 400
rect 474921 391 474979 397
rect 474921 388 474933 391
rect 466052 360 474933 388
rect 466052 348 466058 360
rect 474921 357 474933 360
rect 474967 357 474979 391
rect 474921 351 474979 357
rect 479610 348 479616 400
rect 479668 388 479674 400
rect 492769 391 492827 397
rect 492769 388 492781 391
rect 479668 360 492781 388
rect 479668 348 479674 360
rect 492769 357 492781 360
rect 492815 357 492827 391
rect 492769 351 492827 357
rect 493318 348 493324 400
rect 493376 388 493382 400
rect 508682 388 508688 400
rect 493376 360 508688 388
rect 493376 348 493382 360
rect 508682 348 508688 360
rect 508740 348 508746 400
rect 510246 388 510252 400
rect 510207 360 510252 388
rect 510246 348 510252 360
rect 510304 348 510310 400
rect 510982 348 510988 400
rect 511040 388 511046 400
rect 527634 388 527640 400
rect 511040 360 527640 388
rect 511040 348 511046 360
rect 527634 348 527640 360
rect 527692 348 527698 400
rect 528462 348 528468 400
rect 528520 388 528526 400
rect 545485 391 545543 397
rect 545485 388 545497 391
rect 528520 360 545497 388
rect 528520 348 528526 360
rect 545485 357 545497 360
rect 545531 357 545543 391
rect 561677 391 561735 397
rect 561677 388 561689 391
rect 545485 351 545543 357
rect 552584 360 561689 388
rect 447796 292 450998 320
rect 364794 252 364800 264
rect 356026 224 364800 252
rect 355229 215 355287 221
rect 364794 212 364800 224
rect 364852 212 364858 264
rect 372706 212 372712 264
rect 372764 252 372770 264
rect 383286 252 383292 264
rect 372764 224 383292 252
rect 372764 212 372770 224
rect 383286 212 383292 224
rect 383344 212 383350 264
rect 388070 252 388076 264
rect 383626 224 388076 252
rect 186958 184 186964 196
rect 184906 156 186964 184
rect 17402 76 17408 128
rect 17460 116 17466 128
rect 20070 116 20076 128
rect 17460 88 20076 116
rect 17460 76 17466 88
rect 20070 76 20076 88
rect 20128 76 20134 128
rect 45738 76 45744 128
rect 45796 116 45802 128
rect 47394 116 47400 128
rect 45796 88 47400 116
rect 45796 76 45802 88
rect 47394 76 47400 88
rect 47452 76 47458 128
rect 129826 76 129832 128
rect 129884 116 129890 128
rect 130286 116 130292 128
rect 129884 88 130292 116
rect 129884 76 129890 88
rect 130286 76 130292 88
rect 130344 76 130350 128
rect 155954 76 155960 128
rect 156012 116 156018 128
rect 157518 116 157524 128
rect 156012 88 157524 116
rect 156012 76 156018 88
rect 157518 76 157524 88
rect 157576 76 157582 128
rect 159358 76 159364 128
rect 159416 116 159422 128
rect 161474 116 161480 128
rect 159416 88 161480 116
rect 159416 76 159422 88
rect 161474 76 161480 88
rect 161532 76 161538 128
rect 184290 76 184296 128
rect 184348 116 184354 128
rect 184906 116 184934 156
rect 186958 144 186964 156
rect 187016 144 187022 196
rect 252002 144 252008 196
rect 252060 184 252066 196
rect 257246 184 257252 196
rect 252060 156 257252 184
rect 252060 144 252066 156
rect 257246 144 257252 156
rect 257304 144 257310 196
rect 257982 144 257988 196
rect 258040 184 258046 196
rect 263870 184 263876 196
rect 258040 156 263876 184
rect 258040 144 258046 156
rect 263870 144 263876 156
rect 263928 144 263934 196
rect 282914 144 282920 196
rect 282972 184 282978 196
rect 289998 184 290004 196
rect 282972 156 290004 184
rect 282972 144 282978 156
rect 289998 144 290004 156
rect 290056 144 290062 196
rect 302418 144 302424 196
rect 302476 184 302482 196
rect 310241 187 310299 193
rect 310241 184 310253 187
rect 302476 156 310253 184
rect 302476 144 302482 156
rect 310241 153 310253 156
rect 310287 153 310299 187
rect 310241 147 310299 153
rect 313642 144 313648 196
rect 313700 184 313706 196
rect 321830 184 321836 196
rect 313700 156 321836 184
rect 313700 144 313706 156
rect 321830 144 321836 156
rect 321888 144 321894 196
rect 333146 144 333152 196
rect 333204 184 333210 196
rect 342346 184 342352 196
rect 333204 156 342352 184
rect 333204 144 333210 156
rect 342346 144 342352 156
rect 342404 144 342410 196
rect 346762 144 346768 196
rect 346820 184 346826 196
rect 356054 184 356060 196
rect 346820 156 356060 184
rect 346820 144 346826 156
rect 356054 144 356060 156
rect 356112 144 356118 196
rect 356974 144 356980 196
rect 357032 184 357038 196
rect 365073 187 365131 193
rect 365073 184 365085 187
rect 357032 156 365085 184
rect 357032 144 357038 156
rect 365073 153 365085 156
rect 365119 153 365131 187
rect 365073 147 365131 153
rect 377398 144 377404 196
rect 377456 184 377462 196
rect 383626 184 383654 224
rect 388070 212 388076 224
rect 388128 212 388134 264
rect 389361 255 389419 261
rect 389361 221 389373 255
rect 389407 252 389419 255
rect 397914 252 397920 264
rect 389407 224 397920 252
rect 389407 221 389419 224
rect 389361 215 389419 221
rect 397914 212 397920 224
rect 397972 212 397978 264
rect 398009 255 398067 261
rect 398009 221 398021 255
rect 398055 252 398067 255
rect 404909 255 404967 261
rect 404909 252 404921 255
rect 398055 224 404921 252
rect 398055 221 398067 224
rect 398009 215 398067 221
rect 404909 221 404921 224
rect 404955 221 404967 255
rect 406565 255 406623 261
rect 406565 252 406577 255
rect 404909 215 404967 221
rect 405292 224 406577 252
rect 377456 156 383654 184
rect 377456 144 377462 156
rect 387610 144 387616 196
rect 387668 184 387674 196
rect 399202 184 399208 196
rect 387668 156 399208 184
rect 387668 144 387674 156
rect 399202 144 399208 156
rect 399260 144 399266 196
rect 402330 144 402336 196
rect 402388 184 402394 196
rect 405292 184 405320 224
rect 406565 221 406577 224
rect 406611 221 406623 255
rect 406565 215 406623 221
rect 410334 212 410340 264
rect 410392 252 410398 264
rect 410392 224 415532 252
rect 410392 212 410398 224
rect 402388 156 405320 184
rect 402388 144 402394 156
rect 405642 144 405648 196
rect 405700 184 405706 196
rect 415504 184 415532 224
rect 419442 212 419448 264
rect 419500 252 419506 264
rect 431770 252 431776 264
rect 419500 224 431776 252
rect 419500 212 419506 224
rect 431770 212 431776 224
rect 431828 212 431834 264
rect 431865 255 431923 261
rect 431865 221 431877 255
rect 431911 252 431923 255
rect 435729 255 435787 261
rect 435729 252 435741 255
rect 431911 224 435741 252
rect 431911 221 431923 224
rect 431865 215 431923 221
rect 435729 221 435741 224
rect 435775 221 435787 255
rect 435729 215 435787 221
rect 438762 212 438768 264
rect 438820 252 438826 264
rect 447796 252 447824 292
rect 451918 280 451924 332
rect 451976 320 451982 332
rect 456058 320 456064 332
rect 451976 292 456064 320
rect 451976 280 451982 292
rect 456058 280 456064 292
rect 456116 280 456122 332
rect 461026 280 461032 332
rect 461084 320 461090 332
rect 469769 323 469827 329
rect 461084 292 469720 320
rect 461084 280 461090 292
rect 438820 224 447824 252
rect 438820 212 438826 224
rect 447870 212 447876 264
rect 447928 252 447934 264
rect 461302 252 461308 264
rect 447928 224 461308 252
rect 447928 212 447934 224
rect 461302 212 461308 224
rect 461360 212 461366 264
rect 463602 212 463608 264
rect 463660 252 463666 264
rect 469585 255 469643 261
rect 469585 252 469597 255
rect 463660 224 469597 252
rect 463660 212 463666 224
rect 469585 221 469597 224
rect 469631 221 469643 255
rect 469692 252 469720 292
rect 469769 289 469781 323
rect 469815 320 469827 323
rect 481729 323 481787 329
rect 481729 320 481741 323
rect 469815 292 481741 320
rect 469815 289 469827 292
rect 469769 283 469827 289
rect 481729 289 481741 292
rect 481775 289 481787 323
rect 481729 283 481787 289
rect 482833 323 482891 329
rect 482833 289 482845 323
rect 482879 320 482891 323
rect 482968 320 482974 332
rect 482879 292 482974 320
rect 482879 289 482891 292
rect 482833 283 482891 289
rect 482968 280 482974 292
rect 483026 280 483032 332
rect 484854 280 484860 332
rect 484912 320 484918 332
rect 498010 320 498016 332
rect 484912 292 498016 320
rect 484912 280 484918 292
rect 498010 280 498016 292
rect 498068 280 498074 332
rect 501230 280 501236 332
rect 501288 320 501294 332
rect 508590 320 508596 332
rect 501288 292 508596 320
rect 501288 280 501294 292
rect 508590 280 508596 292
rect 508648 280 508654 332
rect 510338 280 510344 332
rect 510396 320 510402 332
rect 510396 292 519584 320
rect 510396 280 510402 292
rect 475470 252 475476 264
rect 469692 224 475476 252
rect 469585 215 469643 221
rect 475470 212 475476 224
rect 475528 212 475534 264
rect 478506 212 478512 264
rect 478564 252 478570 264
rect 492674 252 492680 264
rect 478564 224 492680 252
rect 478564 212 478570 224
rect 492674 212 492680 224
rect 492732 212 492738 264
rect 492769 255 492827 261
rect 492769 221 492781 255
rect 492815 252 492827 255
rect 494422 252 494428 264
rect 492815 224 494428 252
rect 492815 221 492827 224
rect 492769 215 492827 221
rect 494422 212 494428 224
rect 494480 212 494486 264
rect 497826 212 497832 264
rect 497884 252 497890 264
rect 513834 252 513840 264
rect 497884 224 513840 252
rect 497884 212 497890 224
rect 513834 212 513840 224
rect 513892 212 513898 264
rect 519556 252 519584 292
rect 520366 280 520372 332
rect 520424 320 520430 332
rect 536926 320 536932 332
rect 520424 292 536932 320
rect 520424 280 520430 292
rect 536926 280 536932 292
rect 536984 280 536990 332
rect 537570 280 537576 332
rect 537628 320 537634 332
rect 543458 320 543464 332
rect 537628 292 543464 320
rect 537628 280 537634 292
rect 543458 280 543464 292
rect 543516 280 543522 332
rect 545114 280 545120 332
rect 545172 320 545178 332
rect 552584 320 552612 360
rect 561677 357 561689 360
rect 561723 357 561735 391
rect 561677 351 561735 357
rect 561766 320 561772 332
rect 545172 292 552612 320
rect 552676 292 561772 320
rect 545172 280 545178 292
rect 526438 252 526444 264
rect 519556 224 526444 252
rect 526438 212 526444 224
rect 526496 212 526502 264
rect 543185 255 543243 261
rect 543185 252 543197 255
rect 527146 224 543197 252
rect 422754 184 422760 196
rect 405700 156 414612 184
rect 415504 156 422760 184
rect 405700 144 405706 156
rect 184348 88 184934 116
rect 184348 76 184354 88
rect 185486 76 185492 128
rect 185544 116 185550 128
rect 188246 116 188252 128
rect 185544 88 188252 116
rect 185544 76 185550 88
rect 188246 76 188252 88
rect 188304 76 188310 128
rect 215018 76 215024 128
rect 215076 116 215082 128
rect 219434 116 219440 128
rect 215076 88 219440 116
rect 215076 76 215082 88
rect 219434 76 219440 88
rect 219492 76 219498 128
rect 228542 76 228548 128
rect 228600 116 228606 128
rect 233234 116 233240 128
rect 228600 88 233240 116
rect 228600 76 228606 88
rect 233234 76 233240 88
rect 233292 76 233298 128
rect 266078 76 266084 128
rect 266136 116 266142 128
rect 272150 116 272156 128
rect 266136 88 272156 116
rect 266136 76 266142 88
rect 272150 76 272156 88
rect 272208 76 272214 128
rect 299382 116 299388 128
rect 292546 88 299388 116
rect 16298 8 16304 60
rect 16356 48 16362 60
rect 18966 48 18972 60
rect 16356 20 18972 48
rect 16356 8 16362 20
rect 18966 8 18972 20
rect 19024 8 19030 60
rect 44082 8 44088 60
rect 44140 48 44146 60
rect 46198 48 46204 60
rect 44140 20 46204 48
rect 44140 8 44146 20
rect 46198 8 46204 20
rect 46256 8 46262 60
rect 213822 8 213828 60
rect 213880 48 213886 60
rect 217686 48 217692 60
rect 213880 20 217692 48
rect 213880 8 213886 20
rect 217686 8 217692 20
rect 217744 8 217750 60
rect 227346 8 227352 60
rect 227404 48 227410 60
rect 232038 48 232044 60
rect 227404 20 232044 48
rect 227404 8 227410 20
rect 232038 8 232044 20
rect 232096 8 232102 60
rect 236546 8 236552 60
rect 236604 48 236610 60
rect 241422 48 241428 60
rect 236604 20 241428 48
rect 236604 8 236610 20
rect 241422 8 241428 20
rect 241480 8 241486 60
rect 292206 8 292212 60
rect 292264 48 292270 60
rect 292546 48 292574 88
rect 299382 76 299388 88
rect 299440 76 299446 128
rect 314746 76 314752 128
rect 314804 116 314810 128
rect 314804 88 316034 116
rect 314804 76 314810 88
rect 292264 20 292574 48
rect 316006 48 316034 88
rect 320634 76 320640 128
rect 320692 116 320698 128
rect 329006 116 329012 128
rect 320692 88 329012 116
rect 320692 76 320698 88
rect 329006 76 329012 88
rect 329064 76 329070 128
rect 330846 76 330852 128
rect 330904 116 330910 128
rect 336093 119 336151 125
rect 336093 116 336105 119
rect 330904 88 336105 116
rect 330904 76 330910 88
rect 336093 85 336105 88
rect 336139 85 336151 119
rect 336093 79 336151 85
rect 339494 76 339500 128
rect 339552 116 339558 128
rect 347774 116 347780 128
rect 339552 88 347780 116
rect 339552 76 339558 88
rect 347774 76 347780 88
rect 347832 76 347838 128
rect 358078 76 358084 128
rect 358136 116 358142 128
rect 368201 119 368259 125
rect 368201 116 368213 119
rect 358136 88 368213 116
rect 358136 76 358142 88
rect 368201 85 368213 88
rect 368247 85 368259 119
rect 368201 79 368259 85
rect 370406 76 370412 128
rect 370464 116 370470 128
rect 380894 116 380900 128
rect 370464 88 380900 116
rect 370464 76 370470 88
rect 380894 76 380900 88
rect 380952 76 380958 128
rect 384206 76 384212 128
rect 384264 116 384270 128
rect 384264 88 386414 116
rect 384264 76 384270 88
rect 322842 48 322848 60
rect 316006 20 322848 48
rect 292264 8 292270 20
rect 322842 8 322848 20
rect 322900 8 322906 60
rect 324038 8 324044 60
rect 324096 48 324102 60
rect 332502 48 332508 60
rect 324096 20 332508 48
rect 324096 8 324102 20
rect 332502 8 332508 20
rect 332560 8 332566 60
rect 337194 8 337200 60
rect 337252 48 337258 60
rect 345014 48 345020 60
rect 337252 20 345020 48
rect 337252 8 337258 20
rect 345014 8 345020 20
rect 345072 8 345078 60
rect 347682 8 347688 60
rect 347740 48 347746 60
rect 357342 48 357348 60
rect 347740 20 357348 48
rect 347740 8 347746 20
rect 357342 8 357348 20
rect 357400 8 357406 60
rect 360378 8 360384 60
rect 360436 48 360442 60
rect 370593 51 370651 57
rect 370593 48 370605 51
rect 360436 20 370605 48
rect 360436 8 360442 20
rect 370593 17 370605 20
rect 370639 17 370651 51
rect 370593 11 370651 17
rect 375098 8 375104 60
rect 375156 48 375162 60
rect 385678 48 385684 60
rect 375156 20 385684 48
rect 375156 8 375162 20
rect 385678 8 385684 20
rect 385736 8 385742 60
rect 386386 48 386414 88
rect 386506 76 386512 128
rect 386564 116 386570 128
rect 389361 119 389419 125
rect 389361 116 389373 119
rect 386564 88 389373 116
rect 386564 76 386570 88
rect 389361 85 389373 88
rect 389407 85 389419 119
rect 389361 79 389419 85
rect 390189 119 390247 125
rect 390189 85 390201 119
rect 390235 116 390247 119
rect 393777 119 393835 125
rect 393777 116 393789 119
rect 390235 88 393789 116
rect 390235 85 390247 88
rect 390189 79 390247 85
rect 393777 85 393789 88
rect 393823 85 393835 119
rect 393777 79 393835 85
rect 393958 76 393964 128
rect 394016 116 394022 128
rect 396169 119 396227 125
rect 396169 116 396181 119
rect 394016 88 396181 116
rect 394016 76 394022 88
rect 396169 85 396181 88
rect 396215 85 396227 119
rect 396169 79 396227 85
rect 397454 76 397460 128
rect 397512 116 397518 128
rect 405826 116 405832 128
rect 397512 88 405832 116
rect 397512 76 397518 88
rect 405826 76 405832 88
rect 405884 76 405890 128
rect 406930 76 406936 128
rect 406988 116 406994 128
rect 414584 116 414612 156
rect 422754 144 422760 156
rect 422812 144 422818 196
rect 426986 144 426992 196
rect 427044 184 427050 196
rect 440142 184 440148 196
rect 427044 156 440148 184
rect 427044 144 427050 156
rect 440142 144 440148 156
rect 440200 144 440206 196
rect 441062 144 441068 196
rect 441120 184 441126 196
rect 454497 187 454555 193
rect 454497 184 454509 187
rect 441120 156 454509 184
rect 441120 144 441126 156
rect 454497 153 454509 156
rect 454543 153 454555 187
rect 454497 147 454555 153
rect 462406 144 462412 196
rect 462464 184 462470 196
rect 476666 184 476672 196
rect 462464 156 476672 184
rect 462464 144 462470 156
rect 476666 144 476672 156
rect 476724 144 476730 196
rect 477402 144 477408 196
rect 477460 184 477466 196
rect 483658 184 483664 196
rect 477460 156 483664 184
rect 477460 144 477466 156
rect 483658 144 483664 156
rect 483716 144 483722 196
rect 486050 144 486056 196
rect 486108 184 486114 196
rect 501598 184 501604 196
rect 486108 156 501604 184
rect 486108 144 486114 156
rect 501598 144 501604 156
rect 501656 144 501662 196
rect 507854 144 507860 196
rect 507912 184 507918 196
rect 524046 184 524052 196
rect 507912 156 524052 184
rect 507912 144 507918 156
rect 524046 144 524052 156
rect 524104 144 524110 196
rect 526254 144 526260 196
rect 526312 184 526318 196
rect 527146 184 527174 224
rect 543185 221 543197 224
rect 543231 221 543243 255
rect 543185 215 543243 221
rect 544194 212 544200 264
rect 544252 252 544258 264
rect 552676 252 552704 292
rect 561766 280 561772 292
rect 561824 280 561830 332
rect 561876 320 561904 428
rect 562594 416 562600 428
rect 562652 416 562658 468
rect 561953 391 562011 397
rect 561953 357 561965 391
rect 561999 388 562011 391
rect 563054 388 563060 400
rect 561999 360 563060 388
rect 561999 357 562011 360
rect 561953 351 562011 357
rect 563054 348 563060 360
rect 563112 348 563118 400
rect 565446 320 565452 332
rect 561876 292 565452 320
rect 565446 280 565452 292
rect 565504 280 565510 332
rect 544252 224 552704 252
rect 544252 212 544258 224
rect 553302 212 553308 264
rect 553360 252 553366 264
rect 571150 252 571156 264
rect 553360 224 571156 252
rect 553360 212 553366 224
rect 571150 212 571156 224
rect 571208 212 571214 264
rect 526312 156 527174 184
rect 526312 144 526318 156
rect 535270 144 535276 196
rect 535328 184 535334 196
rect 552382 184 552388 196
rect 535328 156 552388 184
rect 535328 144 535334 156
rect 552382 144 552388 156
rect 552440 144 552446 196
rect 554590 144 554596 196
rect 554648 184 554654 196
rect 572898 184 572904 196
rect 554648 156 572904 184
rect 554648 144 554654 156
rect 572898 144 572904 156
rect 572956 144 572962 196
rect 417694 116 417700 128
rect 406988 88 411254 116
rect 414584 88 417700 116
rect 406988 76 406994 88
rect 395522 48 395528 60
rect 386386 20 395528 48
rect 395522 8 395528 20
rect 395580 8 395586 60
rect 396258 8 396264 60
rect 396316 48 396322 60
rect 405090 48 405096 60
rect 396316 20 405096 48
rect 396316 8 396322 20
rect 405090 8 405096 20
rect 405148 8 405154 60
rect 411226 48 411254 88
rect 417694 76 417700 88
rect 417752 76 417758 128
rect 428090 76 428096 128
rect 428148 116 428154 128
rect 431773 119 431831 125
rect 431773 116 431785 119
rect 428148 88 431785 116
rect 428148 76 428154 88
rect 431773 85 431785 88
rect 431819 85 431831 119
rect 431773 79 431831 85
rect 431862 76 431868 128
rect 431920 116 431926 128
rect 444742 116 444748 128
rect 431920 88 444748 116
rect 431920 76 431926 88
rect 444742 76 444748 88
rect 444800 76 444806 128
rect 445570 76 445576 128
rect 445628 116 445634 128
rect 455877 119 455935 125
rect 455877 116 455889 119
rect 445628 88 455889 116
rect 445628 76 445634 88
rect 455877 85 455889 88
rect 455923 85 455935 119
rect 455877 79 455935 85
rect 459002 76 459008 128
rect 459060 116 459066 128
rect 473262 116 473268 128
rect 459060 88 473268 116
rect 459060 76 459066 88
rect 473262 76 473268 88
rect 473320 76 473326 128
rect 473998 76 474004 128
rect 474056 116 474062 128
rect 483198 116 483204 128
rect 474056 88 483204 116
rect 474056 76 474062 88
rect 483198 76 483204 88
rect 483256 76 483262 128
rect 488534 76 488540 128
rect 488592 116 488598 128
rect 503990 116 503996 128
rect 488592 88 503996 116
rect 488592 76 488598 88
rect 503990 76 503996 88
rect 504048 76 504054 128
rect 504634 76 504640 128
rect 504692 116 504698 128
rect 520550 116 520556 128
rect 504692 88 520556 116
rect 504692 76 504698 88
rect 520550 76 520556 88
rect 520608 76 520614 128
rect 522850 76 522856 128
rect 522908 116 522914 128
rect 539778 116 539784 128
rect 522908 88 539784 116
rect 522908 76 522914 88
rect 539778 76 539784 88
rect 539836 76 539842 128
rect 546494 76 546500 128
rect 546552 116 546558 128
rect 564618 116 564624 128
rect 546552 88 564624 116
rect 546552 76 546558 88
rect 564618 76 564624 88
rect 564676 76 564682 128
rect 418798 48 418804 60
rect 411226 20 418804 48
rect 418798 8 418804 20
rect 418856 8 418862 60
rect 425790 8 425796 60
rect 425848 48 425854 60
rect 438854 48 438860 60
rect 425848 20 438860 48
rect 425848 8 425854 20
rect 438854 8 438860 20
rect 438912 8 438918 60
rect 439866 48 439872 60
rect 439827 20 439872 48
rect 439866 8 439872 20
rect 439924 8 439930 60
rect 449618 8 449624 60
rect 449676 48 449682 60
rect 462130 48 462136 60
rect 449676 20 462136 48
rect 449676 8 449682 20
rect 462130 8 462136 20
rect 462188 8 462194 60
rect 464890 8 464896 60
rect 464948 48 464954 60
rect 479518 48 479524 60
rect 464948 20 479524 48
rect 464948 8 464954 20
rect 479518 8 479524 20
rect 479576 8 479582 60
rect 482646 8 482652 60
rect 482704 48 482710 60
rect 498197 51 498255 57
rect 498197 48 498209 51
rect 482704 20 498209 48
rect 482704 8 482710 20
rect 498197 17 498209 20
rect 498243 17 498255 51
rect 498197 11 498255 17
rect 498930 8 498936 60
rect 498988 48 498994 60
rect 514938 48 514944 60
rect 498988 20 514944 48
rect 498988 8 498994 20
rect 514938 8 514944 20
rect 514996 8 515002 60
rect 521562 8 521568 60
rect 521620 48 521626 60
rect 538030 48 538036 60
rect 521620 20 538036 48
rect 521620 8 521626 20
rect 538030 8 538036 20
rect 538088 8 538094 60
rect 539870 8 539876 60
rect 539928 48 539934 60
rect 557166 48 557172 60
rect 539928 20 557172 48
rect 539928 8 539934 20
rect 557166 8 557172 20
rect 557224 8 557230 60
rect 561398 8 561404 60
rect 561456 48 561462 60
rect 580718 48 580724 60
rect 561456 20 580724 48
rect 561456 8 561462 20
rect 580718 8 580724 20
rect 580776 8 580782 60
<< via1 >>
rect 235448 703808 235500 703860
rect 300860 703808 300912 703860
rect 271788 703740 271840 703792
rect 364708 703740 364760 703792
rect 170496 703672 170548 703724
rect 315488 703672 315540 703724
rect 257252 703604 257304 703656
rect 429660 703604 429712 703656
rect 242440 703536 242492 703588
rect 494428 703536 494480 703588
rect 227628 703468 227680 703520
rect 503904 703468 503956 703520
rect 105452 703400 105504 703452
rect 330300 703400 330352 703452
rect 40500 703332 40552 703384
rect 345020 703332 345072 703384
rect 1584 703264 1636 703316
rect 359740 703264 359792 703316
rect 213000 703196 213052 703248
rect 576400 703196 576452 703248
rect 1676 703128 1728 703180
rect 374460 703128 374512 703180
rect 198280 703060 198332 703112
rect 575020 703060 575072 703112
rect 1768 702992 1820 703044
rect 389180 702992 389232 703044
rect 183376 702924 183428 702976
rect 573640 702924 573692 702976
rect 1860 702856 1912 702908
rect 403900 702856 403952 702908
rect 139308 702788 139360 702840
rect 572168 702788 572220 702840
rect 2504 702720 2556 702772
rect 448152 702720 448204 702772
rect 480 702652 532 702704
rect 477592 702652 477644 702704
rect 296 702584 348 702636
rect 507124 702584 507176 702636
rect 20 702516 72 702568
rect 536840 702516 536892 702568
rect 21456 702448 21508 702500
rect 576124 702448 576176 702500
rect 276020 702380 276072 702432
rect 305736 702380 305788 702432
rect 4344 702312 4396 702364
rect 472716 702312 472768 702364
rect 247408 702244 247460 702296
rect 313280 702244 313332 702296
rect 280988 702176 281040 702228
rect 384304 702176 384356 702228
rect 232688 702108 232740 702160
rect 349804 702108 349856 702160
rect 154028 702040 154080 702092
rect 291844 702040 291896 702092
rect 178592 701972 178644 702024
rect 325608 701972 325660 702024
rect 75460 701904 75512 701956
rect 232872 701904 232924 701956
rect 260840 701904 260892 701956
rect 399024 701904 399076 701956
rect 114284 701836 114336 701888
rect 277492 701836 277544 701888
rect 282920 701836 282972 701888
rect 320456 701836 320508 701888
rect 320916 701836 320968 701888
rect 482560 701836 482612 701888
rect 224960 701768 225012 701820
rect 414204 701768 414256 701820
rect 104808 701700 104860 701752
rect 340880 701700 340932 701752
rect 6644 701632 6696 701684
rect 252284 701632 252336 701684
rect 253204 701632 253256 701684
rect 453028 701632 453080 701684
rect 148968 701564 149020 701616
rect 567844 701564 567896 701616
rect 4252 701496 4304 701548
rect 428464 701496 428516 701548
rect 144276 701428 144328 701480
rect 574928 701428 574980 701480
rect 134432 701360 134484 701412
rect 576216 701360 576268 701412
rect 129464 701292 129516 701344
rect 573456 701292 573508 701344
rect 2412 701224 2464 701276
rect 458180 701224 458232 701276
rect 119712 701156 119764 701208
rect 574836 701156 574888 701208
rect 572 701088 624 701140
rect 467840 701088 467892 701140
rect 72976 700952 73028 701004
rect 335360 701020 335412 701072
rect 340972 701020 341024 701072
rect 512000 701020 512052 701072
rect 556896 701020 556948 701072
rect 564440 701020 564492 701072
rect 137836 700884 137888 700936
rect 282920 700884 282972 700936
rect 284116 700884 284168 700936
rect 295892 700884 295944 700936
rect 298008 700884 298060 700936
rect 300124 700884 300176 700936
rect 313280 700884 313332 700936
rect 462320 700884 462372 700936
rect 503904 700884 503956 700936
rect 559656 700884 559708 700936
rect 154120 700816 154172 700868
rect 325332 700816 325384 700868
rect 325608 700816 325660 700868
rect 580724 700816 580776 700868
rect 3792 700748 3844 700800
rect 207020 700748 207072 700800
rect 252284 700748 252336 700800
rect 478512 700748 478564 700800
rect 3332 700680 3384 700732
rect 253204 700680 253256 700732
rect 267004 700680 267056 700732
rect 413652 700680 413704 700732
rect 89168 700612 89220 700664
rect 340052 700612 340104 700664
rect 340880 700612 340932 700664
rect 580448 700612 580500 700664
rect 3148 700544 3200 700596
rect 260840 700544 260892 700596
rect 267648 700544 267700 700596
rect 2964 700476 3016 700528
rect 280988 700544 281040 700596
rect 332508 700544 332560 700596
rect 349804 700544 349856 700596
rect 527180 700544 527232 700596
rect 291384 700476 291436 700528
rect 291844 700476 291896 700528
rect 580632 700476 580684 700528
rect 4068 700408 4120 700460
rect 224960 700408 225012 700460
rect 237104 700408 237156 700460
rect 543464 700408 543516 700460
rect 24308 700340 24360 700392
rect 354956 700340 355008 700392
rect 8116 700272 8168 700324
rect 349896 700272 349948 700324
rect 262128 700204 262180 700256
rect 397460 700204 397512 700256
rect 218980 700136 219032 700188
rect 310934 700136 310986 700188
rect 202788 700068 202840 700120
rect 276020 700068 276072 700120
rect 276526 700068 276578 700120
rect 281494 700068 281546 700120
rect 348792 700068 348844 700120
rect 217876 700000 217928 700052
rect 563520 700000 563572 700052
rect 222844 699932 222896 699984
rect 579068 699932 579120 699984
rect 1032 699864 1084 699916
rect 364616 699864 364668 699916
rect 208124 699796 208176 699848
rect 570880 699796 570932 699848
rect 3056 699728 3108 699780
rect 369768 699728 369820 699780
rect 193220 699660 193272 699712
rect 578976 699660 579028 699712
rect 277492 699592 277544 699644
rect 580540 699592 580592 699644
rect 3976 699524 4028 699576
rect 320916 699524 320968 699576
rect 3700 699456 3752 699508
rect 340972 699456 341024 699508
rect 379520 699499 379572 699508
rect 379520 699465 379529 699499
rect 379529 699465 379563 699499
rect 379563 699465 379572 699499
rect 379520 699456 379572 699465
rect 386236 699499 386288 699508
rect 386236 699465 386245 699499
rect 386245 699465 386279 699499
rect 386279 699465 386288 699499
rect 386236 699456 386288 699465
rect 394148 699499 394200 699508
rect 394148 699465 394157 699499
rect 394157 699465 394191 699499
rect 394191 699465 394200 699499
rect 394148 699456 394200 699465
rect 408868 699499 408920 699508
rect 408868 699465 408877 699499
rect 408877 699465 408911 699499
rect 408911 699465 408920 699499
rect 408868 699456 408920 699465
rect 423680 699499 423732 699508
rect 423680 699465 423689 699499
rect 423689 699465 423723 699499
rect 423723 699465 423732 699499
rect 423680 699456 423732 699465
rect 438308 699499 438360 699508
rect 438308 699465 438317 699499
rect 438317 699465 438351 699499
rect 438351 699465 438360 699499
rect 438308 699456 438360 699465
rect 521844 699499 521896 699508
rect 521844 699465 521853 699499
rect 521853 699465 521887 699499
rect 521887 699465 521896 699499
rect 521844 699456 521896 699465
rect 232872 699388 232924 699440
rect 580356 699388 580408 699440
rect 35992 699363 36044 699372
rect 35992 699329 36001 699363
rect 36001 699329 36035 699363
rect 36035 699329 36044 699363
rect 35992 699320 36044 699329
rect 65616 699363 65668 699372
rect 65616 699329 65625 699363
rect 65625 699329 65659 699363
rect 65659 699329 65668 699363
rect 65616 699320 65668 699329
rect 70400 699363 70452 699372
rect 70400 699329 70409 699363
rect 70409 699329 70443 699363
rect 70443 699329 70452 699363
rect 70400 699320 70452 699329
rect 80152 699363 80204 699372
rect 80152 699329 80161 699363
rect 80161 699329 80195 699363
rect 80195 699329 80204 699363
rect 80152 699320 80204 699329
rect 85304 699363 85356 699372
rect 85304 699329 85313 699363
rect 85313 699329 85347 699363
rect 85347 699329 85356 699363
rect 85304 699320 85356 699329
rect 100024 699363 100076 699372
rect 100024 699329 100033 699363
rect 100033 699329 100067 699363
rect 100067 699329 100076 699363
rect 100024 699320 100076 699329
rect 109868 699363 109920 699372
rect 109868 699329 109877 699363
rect 109877 699329 109911 699363
rect 109911 699329 109920 699363
rect 109868 699320 109920 699329
rect 158812 699363 158864 699372
rect 158812 699329 158821 699363
rect 158821 699329 158855 699363
rect 158855 699329 158864 699363
rect 158812 699320 158864 699329
rect 168840 699363 168892 699372
rect 168840 699329 168849 699363
rect 168849 699329 168883 699363
rect 168883 699329 168892 699363
rect 168840 699320 168892 699329
rect 173716 699363 173768 699372
rect 173716 699329 173725 699363
rect 173725 699329 173759 699363
rect 173759 699329 173768 699363
rect 173716 699320 173768 699329
rect 188436 699363 188488 699372
rect 188436 699329 188445 699363
rect 188445 699329 188479 699363
rect 188479 699329 188488 699363
rect 188436 699320 188488 699329
rect 202972 699320 203024 699372
rect 573732 699320 573784 699372
rect 940 699252 992 699304
rect 569592 699184 569644 699236
rect 848 699116 900 699168
rect 565360 699048 565412 699100
rect 573548 698980 573600 699032
rect 756 698912 808 698964
rect 578884 698844 578936 698896
rect 664 698776 716 698828
rect 2596 698708 2648 698760
rect 569500 698640 569552 698692
rect 572076 698572 572128 698624
rect 571984 698504 572036 698556
rect 566740 698436 566792 698488
rect 569408 698368 569460 698420
rect 566556 698300 566608 698352
rect 563520 698232 563572 698284
rect 580172 698232 580224 698284
rect 204 697620 256 697672
rect 3424 697484 3476 697536
rect 574744 697552 574796 697604
rect 576400 671984 576452 672036
rect 579620 671984 579672 672036
rect 573732 644376 573784 644428
rect 580172 644376 580224 644428
rect 570880 632000 570932 632052
rect 580172 632000 580224 632052
rect 3056 619080 3108 619132
rect 4252 619080 4304 619132
rect 575020 618196 575072 618248
rect 580172 618196 580224 618248
rect 569592 591948 569644 592000
rect 580172 591948 580224 592000
rect 573640 564340 573692 564392
rect 580172 564340 580224 564392
rect 573548 538160 573600 538212
rect 580172 538160 580224 538212
rect 3148 514768 3200 514820
rect 4344 514768 4396 514820
rect 565360 511912 565412 511964
rect 580172 511912 580224 511964
rect 576308 471928 576360 471980
rect 579804 471928 579856 471980
rect 574928 431876 574980 431928
rect 579712 431876 579764 431928
rect 567844 419432 567896 419484
rect 580172 419432 580224 419484
rect 572168 405628 572220 405680
rect 580172 405628 580224 405680
rect 573456 379448 573508 379500
rect 579620 379448 579672 379500
rect 576216 365644 576268 365696
rect 580172 365644 580224 365696
rect 570788 353200 570840 353252
rect 580172 353200 580224 353252
rect 574836 313216 574888 313268
rect 579712 313216 579764 313268
rect 569500 299412 569552 299464
rect 579804 299412 579856 299464
rect 572076 273164 572128 273216
rect 580172 273164 580224 273216
rect 565268 245556 565320 245608
rect 580172 245556 580224 245608
rect 571984 233180 572036 233232
rect 580172 233180 580224 233232
rect 573364 219376 573416 219428
rect 580172 219376 580224 219428
rect 566740 206932 566792 206984
rect 579896 206932 579948 206984
rect 569408 193128 569460 193180
rect 580172 193128 580224 193180
rect 566556 166948 566608 167000
rect 580172 166948 580224 167000
rect 569316 153144 569368 153196
rect 579804 153144 579856 153196
rect 570696 139340 570748 139392
rect 580172 139340 580224 139392
rect 565176 126896 565228 126948
rect 580172 126896 580224 126948
rect 566648 113092 566700 113144
rect 580172 113092 580224 113144
rect 570604 100648 570656 100700
rect 580172 100648 580224 100700
rect 574744 86912 574796 86964
rect 580172 86912 580224 86964
rect 565084 73108 565136 73160
rect 579988 73108 580040 73160
rect 569224 60664 569276 60716
rect 580172 60664 580224 60716
rect 576124 46860 576176 46912
rect 580172 46860 580224 46912
rect 566464 33056 566516 33108
rect 580172 33056 580224 33108
rect 577504 20612 577556 20664
rect 579712 20612 579764 20664
rect 569868 3068 569920 3120
rect 577412 3068 577464 3120
rect 563704 3000 563756 3052
rect 583392 3000 583444 3052
rect 563520 2932 563572 2984
rect 573916 2932 573968 2984
rect 563612 2864 563664 2916
rect 575480 2864 575532 2916
rect 582196 2864 582248 2916
rect 576308 2796 576360 2848
rect 2964 2048 3016 2100
rect 564440 2048 564492 2100
rect 565912 1368 565964 1420
rect 569132 1368 569184 1420
rect 566832 1164 566884 1216
rect 563612 1096 563664 1148
rect 4068 688 4120 740
rect 1676 620 1728 672
rect 5356 620 5408 672
rect 7748 620 7800 672
rect 11060 620 11112 672
rect 14464 620 14516 672
rect 19432 620 19484 672
rect 22376 620 22428 672
rect 23020 620 23072 672
rect 25780 620 25832 672
rect 28816 620 28868 672
rect 31668 620 31720 672
rect 32404 620 32456 672
rect 34888 620 34940 672
rect 38384 620 38436 672
rect 572 552 624 604
rect 4252 552 4304 604
rect 5264 552 5316 604
rect 6460 552 6512 604
rect 7656 552 7708 604
rect 10324 484 10376 536
rect 12348 552 12400 604
rect 15568 552 15620 604
rect 18512 552 18564 604
rect 21272 552 21324 604
rect 21824 552 21876 604
rect 24860 552 24912 604
rect 25320 552 25372 604
rect 28080 552 28132 604
rect 28724 552 28776 604
rect 29184 552 29236 604
rect 30104 552 30156 604
rect 32588 552 32640 604
rect 33600 552 33652 604
rect 36084 552 36136 604
rect 37188 552 37240 604
rect 11520 484 11572 536
rect 13360 484 13412 536
rect 16672 484 16724 536
rect 31484 484 31536 536
rect 33784 484 33836 536
rect 3240 416 3292 468
rect 6644 416 6696 468
rect 24860 416 24912 468
rect 26884 416 26936 468
rect 8944 348 8996 400
rect 14556 348 14608 400
rect 17868 348 17920 400
rect 39580 552 39632 604
rect 40684 620 40736 672
rect 42800 620 42852 672
rect 46664 620 46716 672
rect 48504 620 48556 672
rect 48964 620 49016 672
rect 50804 620 50856 672
rect 63224 620 63276 672
rect 40776 552 40828 604
rect 41880 552 41932 604
rect 43996 552 44048 604
rect 47860 552 47912 604
rect 49608 552 49660 604
rect 50160 552 50212 604
rect 51356 552 51408 604
rect 53012 552 53064 604
rect 54944 552 54996 604
rect 56416 552 56468 604
rect 62028 552 62080 604
rect 63316 552 63368 604
rect 64328 620 64380 672
rect 65616 620 65668 672
rect 66720 620 66772 672
rect 68008 620 68060 672
rect 69112 620 69164 672
rect 70584 620 70636 672
rect 133236 620 133288 672
rect 134156 620 134208 672
rect 136180 620 136232 672
rect 137652 620 137704 672
rect 138756 620 138808 672
rect 140044 620 140096 672
rect 151360 620 151412 672
rect 153016 620 153068 672
rect 153660 620 153712 672
rect 155408 620 155460 672
rect 162768 620 162820 672
rect 164884 620 164936 672
rect 64420 552 64472 604
rect 65524 552 65576 604
rect 66812 552 66864 604
rect 70308 552 70360 604
rect 71228 552 71280 604
rect 76196 552 76248 604
rect 76932 552 76984 604
rect 77392 552 77444 604
rect 78036 552 78088 604
rect 78588 552 78640 604
rect 79140 552 79192 604
rect 79692 552 79744 604
rect 80336 552 80388 604
rect 80888 552 80940 604
rect 81440 552 81492 604
rect 82084 552 82136 604
rect 82728 552 82780 604
rect 121828 552 121880 604
rect 122288 552 122340 604
rect 124128 552 124180 604
rect 124680 552 124732 604
rect 125232 552 125284 604
rect 125876 552 125928 604
rect 126428 552 126480 604
rect 126980 552 127032 604
rect 127532 552 127584 604
rect 128176 552 128228 604
rect 128636 552 128688 604
rect 129372 552 129424 604
rect 133880 552 133932 604
rect 135260 552 135312 604
rect 136456 552 136508 604
rect 137560 552 137612 604
rect 138848 552 138900 604
rect 139952 552 140004 604
rect 141240 552 141292 604
rect 144552 552 144604 604
rect 145932 552 145984 604
rect 146852 552 146904 604
rect 148324 552 148376 604
rect 152556 552 152608 604
rect 154212 552 154264 604
rect 154764 552 154816 604
rect 156604 552 156656 604
rect 157064 552 157116 604
rect 158904 552 158956 604
rect 161572 552 161624 604
rect 163688 552 163740 604
rect 51908 484 51960 536
rect 67732 484 67784 536
rect 69388 484 69440 536
rect 134984 484 135036 536
rect 141056 484 141108 536
rect 142068 484 142120 536
rect 158168 484 158220 536
rect 159732 484 159784 536
rect 42156 416 42208 468
rect 163412 416 163464 468
rect 166080 620 166132 672
rect 167092 620 167144 672
rect 169576 620 169628 672
rect 180892 620 180944 672
rect 183744 620 183796 672
rect 165988 552 166040 604
rect 168380 552 168432 604
rect 170680 552 170732 604
rect 173164 552 173216 604
rect 179788 552 179840 604
rect 182548 552 182600 604
rect 183192 552 183244 604
rect 186136 620 186188 672
rect 191104 620 191156 672
rect 194416 620 194468 672
rect 211620 620 211672 672
rect 215668 620 215720 672
rect 220176 620 220228 672
rect 225328 620 225380 672
rect 226156 620 226208 672
rect 231032 620 231084 672
rect 190000 552 190052 604
rect 193220 552 193272 604
rect 196808 552 196860 604
rect 187700 484 187752 536
rect 191012 484 191064 536
rect 192944 484 192996 536
rect 39856 348 39908 400
rect 42892 348 42944 400
rect 45100 348 45152 400
rect 71320 348 71372 400
rect 72332 348 72384 400
rect 72424 348 72476 400
rect 73528 348 73580 400
rect 73620 348 73672 400
rect 74632 348 74684 400
rect 130936 348 130988 400
rect 131948 348 132000 400
rect 132040 348 132092 400
rect 133144 348 133196 400
rect 160468 348 160520 400
rect 162676 348 162728 400
rect 188804 348 188856 400
rect 192208 348 192260 400
rect 195244 348 195296 400
rect 199108 552 199160 604
rect 203616 552 203668 604
rect 204168 552 204220 604
rect 205732 552 205784 604
rect 209780 552 209832 604
rect 210424 552 210476 604
rect 212172 552 212224 604
rect 214472 552 214524 604
rect 219532 552 219584 604
rect 223948 552 224000 604
rect 225052 552 225104 604
rect 208400 484 208452 536
rect 218428 484 218480 536
rect 222936 484 222988 536
rect 227352 484 227404 536
rect 229836 552 229888 604
rect 229652 484 229704 536
rect 234620 620 234672 672
rect 235448 620 235500 672
rect 240508 620 240560 672
rect 241152 620 241204 672
rect 231860 552 231912 604
rect 237012 552 237064 604
rect 238116 552 238168 604
rect 238852 552 238904 604
rect 244096 552 244148 604
rect 233148 484 233200 536
rect 239956 484 240008 536
rect 245200 552 245252 604
rect 245752 620 245804 672
rect 247960 663 248012 672
rect 247960 629 247969 663
rect 247969 629 248003 663
rect 248003 629 248012 663
rect 247960 620 248012 629
rect 253480 620 253532 672
rect 254584 620 254636 672
rect 246028 552 246080 604
rect 244556 484 244608 536
rect 249984 552 250036 604
rect 251180 552 251232 604
rect 252376 595 252428 604
rect 252376 561 252385 595
rect 252385 561 252419 595
rect 252419 561 252428 595
rect 252376 552 252428 561
rect 254676 552 254728 604
rect 257068 552 257120 604
rect 257252 620 257304 672
rect 258264 620 258316 672
rect 260472 620 260524 672
rect 266544 620 266596 672
rect 260656 552 260708 604
rect 262680 552 262732 604
rect 268844 620 268896 672
rect 272892 620 272944 672
rect 267740 552 267792 604
rect 249064 484 249116 536
rect 261576 484 261628 536
rect 212540 416 212592 468
rect 216588 416 216640 468
rect 222476 416 222528 468
rect 234344 416 234396 468
rect 239036 416 239088 468
rect 253112 416 253164 468
rect 259092 416 259144 468
rect 263692 416 263744 468
rect 270040 552 270092 604
rect 270684 552 270736 604
rect 276756 552 276808 604
rect 277492 620 277544 672
rect 284300 620 284352 672
rect 279516 552 279568 604
rect 280712 595 280764 604
rect 280712 561 280721 595
rect 280721 561 280755 595
rect 280755 561 280764 595
rect 280712 552 280764 561
rect 281816 552 281868 604
rect 285404 552 285456 604
rect 268384 484 268436 536
rect 274548 484 274600 536
rect 278596 484 278648 536
rect 269488 416 269540 468
rect 276204 416 276256 468
rect 279240 416 279292 468
rect 286600 620 286652 672
rect 288992 620 289044 672
rect 291108 620 291160 672
rect 293408 620 293460 672
rect 287612 552 287664 604
rect 294880 552 294932 604
rect 294512 484 294564 536
rect 298468 620 298520 672
rect 300216 620 300268 672
rect 295616 552 295668 604
rect 303160 552 303212 604
rect 307668 620 307720 672
rect 307944 552 307996 604
rect 309048 552 309100 604
rect 309968 620 310020 672
rect 310244 595 310296 604
rect 310244 561 310253 595
rect 310253 561 310287 595
rect 310287 561 310296 595
rect 310244 552 310296 561
rect 311440 552 311492 604
rect 312636 595 312688 604
rect 312636 561 312645 595
rect 312645 561 312679 595
rect 312679 561 312688 595
rect 312636 552 312688 561
rect 288808 416 288860 468
rect 294604 416 294656 468
rect 300584 484 300636 536
rect 301320 484 301372 536
rect 301780 416 301832 468
rect 303620 416 303672 468
rect 315948 620 316000 672
rect 318524 620 318576 672
rect 324412 620 324464 672
rect 325148 620 325200 672
rect 333612 620 333664 672
rect 335360 620 335412 672
rect 316224 552 316276 604
rect 317144 552 317196 604
rect 325608 552 325660 604
rect 327448 552 327500 604
rect 319352 484 319404 536
rect 327816 484 327868 536
rect 329748 484 329800 536
rect 338672 620 338724 672
rect 340880 663 340932 672
rect 340880 629 340889 663
rect 340889 629 340923 663
rect 340923 629 340932 663
rect 340880 620 340932 629
rect 344560 620 344612 672
rect 339868 552 339920 604
rect 342076 552 342128 604
rect 347780 620 347832 672
rect 349252 620 349304 672
rect 349068 552 349120 604
rect 351276 552 351328 604
rect 360844 620 360896 672
rect 355232 595 355284 604
rect 355232 561 355241 595
rect 355241 561 355275 595
rect 355275 561 355284 595
rect 355232 552 355284 561
rect 355876 552 355928 604
rect 351184 484 351236 536
rect 352472 484 352524 536
rect 361948 484 362000 536
rect 312452 416 312504 468
rect 320732 416 320784 468
rect 322848 416 322900 468
rect 331220 416 331272 468
rect 331956 416 332008 468
rect 341156 416 341208 468
rect 343180 416 343232 468
rect 350632 416 350684 468
rect 353576 416 353628 468
rect 217232 348 217284 400
rect 221740 348 221792 400
rect 243360 348 243412 400
rect 248972 348 249024 400
rect 250904 348 250956 400
rect 259276 348 259328 400
rect 264980 348 265032 400
rect 271788 348 271840 400
rect 278504 348 278556 400
rect 280436 348 280488 400
rect 285680 348 285732 400
rect 299020 348 299072 400
rect 306932 348 306984 400
rect 311072 348 311124 400
rect 319536 348 319588 400
rect 321560 348 321612 400
rect 330116 348 330168 400
rect 336464 348 336516 400
rect 336556 348 336608 400
rect 345480 348 345532 400
rect 349068 348 349120 400
rect 358452 348 358504 400
rect 246764 280 246816 332
rect 256884 280 256936 332
rect 262772 280 262824 332
rect 275836 280 275888 332
rect 283288 280 283340 332
rect 284116 280 284168 332
rect 291200 280 291252 332
rect 296812 280 296864 332
rect 303988 280 304040 332
rect 304724 280 304776 332
rect 318340 280 318392 332
rect 326620 280 326672 332
rect 344376 280 344428 332
rect 353852 280 353904 332
rect 354680 280 354732 332
rect 359280 416 359332 468
rect 367008 552 367060 604
rect 368204 595 368256 604
rect 368204 561 368213 595
rect 368213 561 368247 595
rect 368247 561 368256 595
rect 368204 552 368256 561
rect 369308 620 369360 672
rect 371608 620 371660 672
rect 374276 620 374328 672
rect 375288 620 375340 672
rect 369400 552 369452 604
rect 370596 595 370648 604
rect 370596 561 370605 595
rect 370605 561 370639 595
rect 370639 561 370648 595
rect 370596 552 370648 561
rect 376484 552 376536 604
rect 377956 620 378008 672
rect 379520 620 379572 672
rect 390284 620 390336 672
rect 394240 620 394292 672
rect 395620 620 395672 672
rect 401140 620 401192 672
rect 380164 552 380216 604
rect 380808 552 380860 604
rect 383108 595 383160 604
rect 366088 527 366140 536
rect 366088 493 366097 527
rect 366097 493 366131 527
rect 366131 493 366140 527
rect 366088 484 366140 493
rect 366732 416 366784 468
rect 373816 484 373868 536
rect 380900 484 380952 536
rect 383108 561 383117 595
rect 383117 561 383151 595
rect 383151 561 383160 595
rect 383108 552 383160 561
rect 389456 595 389508 604
rect 389456 561 389465 595
rect 389465 561 389499 595
rect 389499 561 389508 595
rect 389456 552 389508 561
rect 389916 552 389968 604
rect 392400 552 392452 604
rect 393320 552 393372 604
rect 398840 552 398892 604
rect 391572 484 391624 536
rect 399944 484 399996 536
rect 400312 484 400364 536
rect 403440 484 403492 536
rect 404728 663 404780 672
rect 404728 629 404737 663
rect 404737 629 404771 663
rect 404771 629 404780 663
rect 404728 620 404780 629
rect 404912 663 404964 672
rect 404912 629 404921 663
rect 404921 629 404955 663
rect 404955 629 404964 663
rect 404912 620 404964 629
rect 407212 620 407264 672
rect 413744 663 413796 672
rect 410800 552 410852 604
rect 413100 552 413152 604
rect 413744 629 413753 663
rect 413753 629 413787 663
rect 413787 629 413796 663
rect 413744 620 413796 629
rect 414296 620 414348 672
rect 563520 1028 563572 1080
rect 415492 620 415544 672
rect 416688 620 416740 672
rect 417148 663 417200 672
rect 417148 629 417157 663
rect 417157 629 417191 663
rect 417191 629 417200 663
rect 417148 620 417200 629
rect 418344 620 418396 672
rect 430856 620 430908 672
rect 434444 620 434496 672
rect 419908 552 419960 604
rect 421656 595 421708 604
rect 421656 561 421665 595
rect 421665 561 421699 595
rect 421699 561 421708 595
rect 421656 552 421708 561
rect 422852 595 422904 604
rect 422852 561 422861 595
rect 422861 561 422895 595
rect 422895 561 422904 595
rect 422852 552 422904 561
rect 423772 595 423824 604
rect 423772 561 423781 595
rect 423781 561 423815 595
rect 423815 561 423824 595
rect 423772 552 423824 561
rect 424692 595 424744 604
rect 424692 561 424701 595
rect 424701 561 424735 595
rect 424735 561 424744 595
rect 424692 552 424744 561
rect 424968 552 425020 604
rect 414940 484 414992 536
rect 421748 484 421800 536
rect 424508 484 424560 536
rect 426348 527 426400 536
rect 426348 493 426357 527
rect 426357 493 426391 527
rect 426391 493 426400 527
rect 426348 484 426400 493
rect 429016 527 429068 536
rect 429016 493 429025 527
rect 429025 493 429059 527
rect 429059 493 429068 527
rect 429016 484 429068 493
rect 367836 416 367888 468
rect 375656 416 375708 468
rect 378416 416 378468 468
rect 365996 348 366048 400
rect 376300 348 376352 400
rect 386972 348 387024 400
rect 388812 348 388864 400
rect 391020 348 391072 400
rect 255688 212 255740 264
rect 261944 212 261996 264
rect 264888 212 264940 264
rect 271052 212 271104 264
rect 274088 212 274140 264
rect 289820 212 289872 264
rect 296996 212 297048 264
rect 297916 212 297968 264
rect 305736 212 305788 264
rect 308772 212 308824 264
rect 316592 212 316644 264
rect 326344 212 326396 264
rect 335360 212 335412 264
rect 345572 212 345624 264
rect 363696 280 363748 332
rect 364892 280 364944 332
rect 382004 280 382056 332
rect 393228 280 393280 332
rect 406200 416 406252 468
rect 408132 416 408184 468
rect 411536 416 411588 468
rect 420552 416 420604 468
rect 433248 552 433300 604
rect 435180 620 435232 672
rect 436468 620 436520 672
rect 437940 663 437992 672
rect 437940 629 437949 663
rect 437949 629 437983 663
rect 437983 629 437992 663
rect 437940 620 437992 629
rect 435548 552 435600 604
rect 442632 620 442684 672
rect 448244 620 448296 672
rect 448980 663 449032 672
rect 448980 629 448989 663
rect 448989 629 449023 663
rect 449023 629 449032 663
rect 448980 620 449032 629
rect 429476 484 429528 536
rect 441528 552 441580 604
rect 442172 595 442224 604
rect 442172 561 442181 595
rect 442181 561 442215 595
rect 442215 561 442224 595
rect 442172 552 442224 561
rect 443828 595 443880 604
rect 443828 561 443837 595
rect 443837 561 443871 595
rect 443871 561 443880 595
rect 443828 552 443880 561
rect 444472 552 444524 604
rect 456892 620 456944 672
rect 457996 663 458048 672
rect 457996 629 458005 663
rect 458005 629 458039 663
rect 458039 629 458048 663
rect 457996 620 458048 629
rect 458180 663 458232 672
rect 458180 629 458189 663
rect 458189 629 458223 663
rect 458223 629 458232 663
rect 460204 663 460256 672
rect 458180 620 458232 629
rect 460204 629 460213 663
rect 460213 629 460247 663
rect 460247 629 460256 663
rect 460204 620 460256 629
rect 449992 595 450044 604
rect 449992 561 450001 595
rect 450001 561 450035 595
rect 450035 561 450044 595
rect 451280 595 451332 604
rect 449992 552 450044 561
rect 451280 561 451289 595
rect 451289 561 451323 595
rect 451323 561 451332 595
rect 451280 552 451332 561
rect 452384 595 452436 604
rect 452384 561 452393 595
rect 452393 561 452427 595
rect 452427 561 452436 595
rect 452384 552 452436 561
rect 454500 595 454552 604
rect 454500 561 454509 595
rect 454509 561 454543 595
rect 454543 561 454552 595
rect 454500 552 454552 561
rect 455696 552 455748 604
rect 459192 552 459244 604
rect 462780 620 462832 672
rect 465172 552 465224 604
rect 466276 620 466328 672
rect 471060 620 471112 672
rect 469864 552 469916 604
rect 471704 620 471756 672
rect 472256 663 472308 672
rect 472256 629 472265 663
rect 472265 629 472299 663
rect 472299 629 472308 663
rect 472256 620 472308 629
rect 472808 663 472860 672
rect 472808 629 472817 663
rect 472817 629 472851 663
rect 472851 629 472860 663
rect 472808 620 472860 629
rect 474556 663 474608 672
rect 474556 629 474565 663
rect 474565 629 474599 663
rect 474599 629 474608 663
rect 474556 620 474608 629
rect 480720 620 480772 672
rect 481456 663 481508 672
rect 481456 629 481465 663
rect 481465 629 481499 663
rect 481499 629 481508 663
rect 481456 620 481508 629
rect 475108 595 475160 604
rect 443276 484 443328 536
rect 453488 527 453540 536
rect 430396 459 430448 468
rect 430396 425 430405 459
rect 430405 425 430439 459
rect 430439 425 430448 459
rect 430396 416 430448 425
rect 434260 416 434312 468
rect 447140 416 447192 468
rect 453488 493 453497 527
rect 453497 493 453531 527
rect 453531 493 453540 527
rect 453488 484 453540 493
rect 453580 484 453632 536
rect 466092 484 466144 536
rect 467196 484 467248 536
rect 475108 561 475117 595
rect 475117 561 475151 595
rect 475151 561 475160 595
rect 475108 552 475160 561
rect 476212 595 476264 604
rect 476212 561 476221 595
rect 476221 561 476255 595
rect 476255 561 476264 595
rect 476212 552 476264 561
rect 476580 595 476632 604
rect 476580 561 476589 595
rect 476589 561 476623 595
rect 476623 561 476632 595
rect 476580 552 476632 561
rect 477868 552 477920 604
rect 480628 552 480680 604
rect 483756 663 483808 672
rect 483756 629 483765 663
rect 483765 629 483799 663
rect 483799 629 483808 663
rect 483756 620 483808 629
rect 481732 595 481784 604
rect 481732 561 481741 595
rect 481741 561 481775 595
rect 481775 561 481784 595
rect 481732 552 481784 561
rect 477408 484 477460 536
rect 485228 620 485280 672
rect 487712 663 487764 672
rect 487712 629 487721 663
rect 487721 629 487755 663
rect 487755 629 487764 663
rect 487712 620 487764 629
rect 489920 620 489972 672
rect 491116 663 491168 672
rect 491116 629 491125 663
rect 491125 629 491159 663
rect 491159 629 491168 663
rect 491116 620 491168 629
rect 491300 620 491352 672
rect 484032 552 484084 604
rect 486424 595 486476 604
rect 486424 561 486433 595
rect 486433 561 486467 595
rect 486467 561 486476 595
rect 486424 552 486476 561
rect 487436 552 487488 604
rect 493324 620 493376 672
rect 492128 552 492180 604
rect 569868 960 569920 1012
rect 575480 892 575532 944
rect 455328 416 455380 468
rect 456524 459 456576 468
rect 456524 425 456533 459
rect 456533 425 456567 459
rect 456567 425 456576 459
rect 456524 416 456576 425
rect 399944 348 399996 400
rect 411720 348 411772 400
rect 416044 348 416096 400
rect 428648 348 428700 400
rect 402244 280 402296 332
rect 403440 280 403492 332
rect 409236 280 409288 332
rect 421012 280 421064 332
rect 423496 280 423548 332
rect 436468 348 436520 400
rect 437480 348 437532 400
rect 450636 348 450688 400
rect 433064 280 433116 332
rect 446036 280 446088 332
rect 452292 348 452344 400
rect 454224 348 454276 400
rect 468484 416 468536 468
rect 469220 416 469272 468
rect 489736 484 489788 536
rect 490932 416 490984 468
rect 494428 663 494480 672
rect 494428 629 494437 663
rect 494437 629 494471 663
rect 494471 629 494480 663
rect 494428 620 494480 629
rect 502984 620 503036 672
rect 505744 663 505796 672
rect 505744 629 505753 663
rect 505753 629 505787 663
rect 505787 629 505796 663
rect 505744 620 505796 629
rect 506480 620 506532 672
rect 506940 620 506992 672
rect 509240 663 509292 672
rect 509240 629 509249 663
rect 509249 629 509283 663
rect 509283 629 509292 663
rect 509240 620 509292 629
rect 509700 663 509752 672
rect 509700 629 509709 663
rect 509709 629 509743 663
rect 509743 629 509752 663
rect 509700 620 509752 629
rect 511264 663 511316 672
rect 511264 629 511273 663
rect 511273 629 511307 663
rect 511307 629 511316 663
rect 511264 620 511316 629
rect 512460 663 512512 672
rect 512460 629 512469 663
rect 512469 629 512503 663
rect 512503 629 512512 663
rect 512460 620 512512 629
rect 513288 663 513340 672
rect 513288 629 513297 663
rect 513297 629 513331 663
rect 513331 629 513340 663
rect 513288 620 513340 629
rect 515864 663 515916 672
rect 515864 629 515873 663
rect 515873 629 515907 663
rect 515907 629 515916 663
rect 515864 620 515916 629
rect 517060 663 517112 672
rect 517060 629 517069 663
rect 517069 629 517103 663
rect 517103 629 517112 663
rect 517060 620 517112 629
rect 519360 663 519412 672
rect 519360 629 519369 663
rect 519369 629 519403 663
rect 519403 629 519412 663
rect 519360 620 519412 629
rect 521844 663 521896 672
rect 521844 629 521853 663
rect 521853 629 521887 663
rect 521887 629 521896 663
rect 521844 620 521896 629
rect 523040 620 523092 672
rect 523960 620 524012 672
rect 495348 595 495400 604
rect 495348 561 495357 595
rect 495357 561 495391 595
rect 495391 561 495400 595
rect 495348 552 495400 561
rect 496728 595 496780 604
rect 496728 561 496737 595
rect 496737 561 496771 595
rect 496771 561 496780 595
rect 496728 552 496780 561
rect 498200 595 498252 604
rect 498200 561 498209 595
rect 498209 561 498243 595
rect 498243 561 498252 595
rect 499396 595 499448 604
rect 498200 552 498252 561
rect 499396 561 499405 595
rect 499405 561 499439 595
rect 499439 561 499448 595
rect 499396 552 499448 561
rect 500132 552 500184 604
rect 516140 552 516192 604
rect 518164 552 518216 604
rect 532516 620 532568 672
rect 533068 620 533120 672
rect 535828 663 535880 672
rect 529020 552 529072 604
rect 530124 595 530176 604
rect 530124 561 530133 595
rect 530133 561 530167 595
rect 530167 561 530176 595
rect 530124 552 530176 561
rect 531872 595 531924 604
rect 531872 561 531881 595
rect 531881 561 531915 595
rect 531915 561 531924 595
rect 531872 552 531924 561
rect 533712 595 533764 604
rect 533712 561 533721 595
rect 533721 561 533755 595
rect 533755 561 533764 595
rect 533712 552 533764 561
rect 535828 629 535837 663
rect 535837 629 535871 663
rect 535871 629 535880 663
rect 535828 620 535880 629
rect 536472 663 536524 672
rect 536472 629 536481 663
rect 536481 629 536515 663
rect 536515 629 536524 663
rect 536472 620 536524 629
rect 540796 663 540848 672
rect 540796 629 540805 663
rect 540805 629 540839 663
rect 540839 629 540848 663
rect 540796 620 540848 629
rect 542176 620 542228 672
rect 543188 663 543240 672
rect 543188 629 543197 663
rect 543197 629 543231 663
rect 543231 629 543240 663
rect 543188 620 543240 629
rect 545488 663 545540 672
rect 545488 629 545497 663
rect 545497 629 545531 663
rect 545531 629 545540 663
rect 545488 620 545540 629
rect 565912 824 565964 876
rect 565820 756 565872 808
rect 568028 756 568080 808
rect 553768 620 553820 672
rect 555148 620 555200 672
rect 555792 663 555844 672
rect 555792 629 555801 663
rect 555801 629 555835 663
rect 555835 629 555844 663
rect 555792 620 555844 629
rect 550272 552 550324 604
rect 551192 595 551244 604
rect 551192 561 551201 595
rect 551201 561 551235 595
rect 551235 561 551244 595
rect 551192 552 551244 561
rect 552388 552 552440 604
rect 570328 688 570380 740
rect 556896 620 556948 672
rect 575112 620 575164 672
rect 505100 484 505152 536
rect 507308 527 507360 536
rect 507308 493 507317 527
rect 507317 493 507351 527
rect 507351 493 507360 527
rect 507308 484 507360 493
rect 512184 484 512236 536
rect 529664 484 529716 536
rect 502340 459 502392 468
rect 502340 425 502349 459
rect 502349 425 502383 459
rect 502383 425 502392 459
rect 502340 416 502392 425
rect 503536 416 503588 468
rect 519728 416 519780 468
rect 525064 459 525116 468
rect 525064 425 525073 459
rect 525073 425 525107 459
rect 525107 425 525116 459
rect 525064 416 525116 425
rect 525156 459 525208 468
rect 525156 425 525165 459
rect 525165 425 525199 459
rect 525199 425 525208 459
rect 525156 416 525208 425
rect 534540 416 534592 468
rect 538772 484 538824 536
rect 548892 527 548944 536
rect 548892 493 548901 527
rect 548901 493 548935 527
rect 548935 493 548944 527
rect 548892 484 548944 493
rect 549260 484 549312 536
rect 550088 484 550140 536
rect 565820 552 565872 604
rect 578608 552 578660 604
rect 558000 527 558052 536
rect 558000 493 558009 527
rect 558009 493 558043 527
rect 558043 493 558052 527
rect 558000 484 558052 493
rect 558736 527 558788 536
rect 558736 493 558745 527
rect 558745 493 558779 527
rect 558779 493 558788 527
rect 558736 484 558788 493
rect 560208 484 560260 536
rect 546500 416 546552 468
rect 547696 416 547748 468
rect 562600 459 562652 468
rect 466000 348 466052 400
rect 479616 348 479668 400
rect 493324 348 493376 400
rect 508688 348 508740 400
rect 510252 391 510304 400
rect 510252 357 510261 391
rect 510261 357 510295 391
rect 510295 357 510304 391
rect 510252 348 510304 357
rect 510988 348 511040 400
rect 527640 348 527692 400
rect 528468 348 528520 400
rect 364800 212 364852 264
rect 372712 212 372764 264
rect 383292 212 383344 264
rect 17408 76 17460 128
rect 20076 76 20128 128
rect 45744 76 45796 128
rect 47400 76 47452 128
rect 129832 76 129884 128
rect 130292 76 130344 128
rect 155960 76 156012 128
rect 157524 76 157576 128
rect 159364 76 159416 128
rect 161480 76 161532 128
rect 184296 76 184348 128
rect 186964 144 187016 196
rect 252008 144 252060 196
rect 257252 144 257304 196
rect 257988 144 258040 196
rect 263876 144 263928 196
rect 282920 144 282972 196
rect 290004 144 290056 196
rect 302424 144 302476 196
rect 313648 144 313700 196
rect 321836 144 321888 196
rect 333152 144 333204 196
rect 342352 144 342404 196
rect 346768 144 346820 196
rect 356060 144 356112 196
rect 356980 144 357032 196
rect 377404 144 377456 196
rect 388076 212 388128 264
rect 397920 212 397972 264
rect 387616 144 387668 196
rect 399208 144 399260 196
rect 402336 144 402388 196
rect 410340 212 410392 264
rect 405648 144 405700 196
rect 419448 212 419500 264
rect 431776 212 431828 264
rect 438768 212 438820 264
rect 451924 280 451976 332
rect 456064 280 456116 332
rect 461032 280 461084 332
rect 447876 212 447928 264
rect 461308 212 461360 264
rect 463608 212 463660 264
rect 482974 280 483026 332
rect 484860 280 484912 332
rect 498016 280 498068 332
rect 501236 280 501288 332
rect 508596 280 508648 332
rect 510344 280 510396 332
rect 475476 212 475528 264
rect 478512 212 478564 264
rect 492680 212 492732 264
rect 494428 212 494480 264
rect 497832 212 497884 264
rect 513840 212 513892 264
rect 520372 280 520424 332
rect 536932 280 536984 332
rect 537576 280 537628 332
rect 543464 280 543516 332
rect 545120 280 545172 332
rect 526444 212 526496 264
rect 185492 76 185544 128
rect 188252 76 188304 128
rect 215024 76 215076 128
rect 219440 76 219492 128
rect 228548 76 228600 128
rect 233240 76 233292 128
rect 266084 76 266136 128
rect 272156 76 272208 128
rect 16304 8 16356 60
rect 18972 8 19024 60
rect 44088 8 44140 60
rect 46204 8 46256 60
rect 213828 8 213880 60
rect 217692 8 217744 60
rect 227352 8 227404 60
rect 232044 8 232096 60
rect 236552 8 236604 60
rect 241428 8 241480 60
rect 292212 8 292264 60
rect 299388 76 299440 128
rect 314752 76 314804 128
rect 320640 76 320692 128
rect 329012 76 329064 128
rect 330852 76 330904 128
rect 339500 76 339552 128
rect 347780 76 347832 128
rect 358084 76 358136 128
rect 370412 76 370464 128
rect 380900 76 380952 128
rect 384212 76 384264 128
rect 322848 8 322900 60
rect 324044 8 324096 60
rect 332508 8 332560 60
rect 337200 8 337252 60
rect 345020 8 345072 60
rect 347688 8 347740 60
rect 357348 8 357400 60
rect 360384 8 360436 60
rect 375104 8 375156 60
rect 385684 8 385736 60
rect 386512 76 386564 128
rect 393964 76 394016 128
rect 397460 76 397512 128
rect 405832 76 405884 128
rect 406936 76 406988 128
rect 422760 144 422812 196
rect 426992 144 427044 196
rect 440148 144 440200 196
rect 441068 144 441120 196
rect 462412 144 462464 196
rect 476672 144 476724 196
rect 477408 144 477460 196
rect 483664 144 483716 196
rect 486056 144 486108 196
rect 501604 144 501656 196
rect 507860 144 507912 196
rect 524052 144 524104 196
rect 526260 144 526312 196
rect 544200 212 544252 264
rect 561772 280 561824 332
rect 562600 425 562609 459
rect 562609 425 562643 459
rect 562643 425 562652 459
rect 562600 416 562652 425
rect 563060 348 563112 400
rect 565452 280 565504 332
rect 553308 212 553360 264
rect 571156 212 571208 264
rect 535276 144 535328 196
rect 552388 144 552440 196
rect 554596 144 554648 196
rect 572904 144 572956 196
rect 395528 8 395580 60
rect 396264 8 396316 60
rect 405096 8 405148 60
rect 417700 76 417752 128
rect 428096 76 428148 128
rect 431868 76 431920 128
rect 444748 76 444800 128
rect 445576 76 445628 128
rect 459008 76 459060 128
rect 473268 76 473320 128
rect 474004 76 474056 128
rect 483204 76 483256 128
rect 488540 76 488592 128
rect 503996 76 504048 128
rect 504640 76 504692 128
rect 520556 76 520608 128
rect 522856 76 522908 128
rect 539784 76 539836 128
rect 546500 76 546552 128
rect 564624 76 564676 128
rect 418804 8 418856 60
rect 425796 8 425848 60
rect 438860 8 438912 60
rect 439872 51 439924 60
rect 439872 17 439881 51
rect 439881 17 439915 51
rect 439915 17 439924 51
rect 439872 8 439924 17
rect 449624 8 449676 60
rect 462136 8 462188 60
rect 464896 8 464948 60
rect 479524 8 479576 60
rect 482652 8 482704 60
rect 498936 8 498988 60
rect 514944 8 514996 60
rect 521568 8 521620 60
rect 538036 8 538088 60
rect 539876 8 539928 60
rect 557172 8 557224 60
rect 561404 8 561456 60
rect 580724 8 580776 60
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 170496 703724 170548 703730
rect 170496 703666 170548 703672
rect 1584 703316 1636 703322
rect 1584 703258 1636 703264
rect 480 702704 532 702710
rect 480 702646 532 702652
rect 296 702636 348 702642
rect 296 702578 348 702584
rect 20 702568 72 702574
rect 20 702510 72 702516
rect 32 71913 60 702510
rect 110 701720 166 701729
rect 110 701655 166 701664
rect 124 85241 152 701655
rect 204 697672 256 697678
rect 204 697614 256 697620
rect 216 111217 244 697614
rect 308 171134 336 702578
rect 386 701992 442 702001
rect 386 701927 442 701936
rect 400 258074 428 701927
rect 492 267186 520 702646
rect 572 701140 624 701146
rect 572 701082 624 701088
rect 584 293185 612 701082
rect 1032 699916 1084 699922
rect 1032 699858 1084 699864
rect 940 699304 992 699310
rect 940 699246 992 699252
rect 848 699168 900 699174
rect 848 699110 900 699116
rect 756 698964 808 698970
rect 756 698906 808 698912
rect 664 698828 716 698834
rect 664 698770 716 698776
rect 676 449585 704 698770
rect 768 501809 796 698906
rect 860 553897 888 699110
rect 952 606121 980 699246
rect 1044 658209 1072 699858
rect 1596 684321 1624 703258
rect 1676 703180 1728 703186
rect 1676 703122 1728 703128
rect 1582 684312 1638 684321
rect 1582 684247 1638 684256
rect 1030 658200 1086 658209
rect 1030 658135 1086 658144
rect 1688 632097 1716 703122
rect 1768 703044 1820 703050
rect 1768 702986 1820 702992
rect 1674 632088 1730 632097
rect 1674 632023 1730 632032
rect 938 606112 994 606121
rect 938 606047 994 606056
rect 1780 580009 1808 702986
rect 1860 702908 1912 702914
rect 1860 702850 1912 702856
rect 1766 580000 1822 580009
rect 1766 579935 1822 579944
rect 846 553888 902 553897
rect 846 553823 902 553832
rect 1872 527921 1900 702850
rect 2504 702772 2556 702778
rect 2504 702714 2556 702720
rect 2226 701856 2282 701865
rect 2226 701791 2282 701800
rect 2042 701448 2098 701457
rect 2042 701383 2098 701392
rect 1950 698048 2006 698057
rect 1950 697983 2006 697992
rect 1858 527912 1914 527921
rect 1858 527847 1914 527856
rect 754 501800 810 501809
rect 754 501735 810 501744
rect 1964 475697 1992 697983
rect 1950 475688 2006 475697
rect 1950 475623 2006 475632
rect 662 449576 718 449585
rect 662 449511 718 449520
rect 570 293176 626 293185
rect 570 293111 626 293120
rect 570 267200 626 267209
rect 492 267158 570 267186
rect 570 267135 626 267144
rect 400 258046 612 258074
rect 584 254153 612 258046
rect 570 254144 626 254153
rect 570 254079 626 254088
rect 308 171106 612 171134
rect 584 162897 612 171106
rect 570 162888 626 162897
rect 570 162823 626 162832
rect 202 111208 258 111217
rect 202 111143 258 111152
rect 110 85232 166 85241
rect 110 85167 166 85176
rect 18 71904 74 71913
rect 18 71839 74 71848
rect 2056 58585 2084 701383
rect 2134 697640 2190 697649
rect 2134 697575 2190 697584
rect 2148 214985 2176 697575
rect 2134 214976 2190 214985
rect 2134 214911 2190 214920
rect 2240 188873 2268 701791
rect 2412 701276 2464 701282
rect 2412 701218 2464 701224
rect 2318 697912 2374 697921
rect 2318 697847 2374 697856
rect 2332 319297 2360 697847
rect 2424 358465 2452 701218
rect 2516 371385 2544 702714
rect 4344 702364 4396 702370
rect 4344 702306 4396 702312
rect 4252 701548 4304 701554
rect 4252 701490 4304 701496
rect 3792 700800 3844 700806
rect 3792 700742 3844 700748
rect 3332 700732 3384 700738
rect 3332 700674 3384 700680
rect 3148 700596 3200 700602
rect 3148 700538 3200 700544
rect 2964 700528 3016 700534
rect 2964 700470 3016 700476
rect 2596 698760 2648 698766
rect 2596 698702 2648 698708
rect 2608 397497 2636 698702
rect 2686 698184 2742 698193
rect 2686 698119 2742 698128
rect 2700 423609 2728 698119
rect 2976 619177 3004 700470
rect 3056 699780 3108 699786
rect 3056 699722 3108 699728
rect 3068 671265 3096 699722
rect 3054 671256 3110 671265
rect 3054 671191 3110 671200
rect 2962 619168 3018 619177
rect 2962 619103 3018 619112
rect 3056 619132 3108 619138
rect 3056 619074 3108 619080
rect 3068 462641 3096 619074
rect 3160 566953 3188 700538
rect 3238 700496 3294 700505
rect 3238 700431 3294 700440
rect 3146 566944 3202 566953
rect 3146 566879 3202 566888
rect 3148 514820 3200 514826
rect 3148 514762 3200 514768
rect 3054 462632 3110 462641
rect 3054 462567 3110 462576
rect 2686 423600 2742 423609
rect 2686 423535 2742 423544
rect 2594 397488 2650 397497
rect 2594 397423 2650 397432
rect 2502 371376 2558 371385
rect 2502 371311 2558 371320
rect 2410 358456 2466 358465
rect 2410 358391 2466 358400
rect 2318 319288 2374 319297
rect 2318 319223 2374 319232
rect 3160 306241 3188 514762
rect 3252 410553 3280 700431
rect 3238 410544 3294 410553
rect 3238 410479 3294 410488
rect 3344 345409 3372 700674
rect 3606 699952 3662 699961
rect 3606 699887 3662 699896
rect 3514 698456 3570 698465
rect 3514 698391 3570 698400
rect 3424 697536 3476 697542
rect 3424 697478 3476 697484
rect 3330 345400 3386 345409
rect 3330 345335 3386 345344
rect 3146 306232 3202 306241
rect 3146 306167 3202 306176
rect 2226 188864 2282 188873
rect 2226 188799 2282 188808
rect 2042 58576 2098 58585
rect 2042 58511 2098 58520
rect 3436 19417 3464 697478
rect 3528 45529 3556 698391
rect 3620 97617 3648 699887
rect 3700 699508 3752 699514
rect 3700 699450 3752 699456
rect 3712 136785 3740 699450
rect 3804 149841 3832 700742
rect 4068 700460 4120 700466
rect 4068 700402 4120 700408
rect 3882 700224 3938 700233
rect 3882 700159 3938 700168
rect 3896 201929 3924 700159
rect 3976 699576 4028 699582
rect 3976 699518 4028 699524
rect 3988 241097 4016 699518
rect 4080 514865 4108 700402
rect 4264 619138 4292 701490
rect 4252 619132 4304 619138
rect 4252 619074 4304 619080
rect 4066 514856 4122 514865
rect 4356 514826 4384 702306
rect 6644 701684 6696 701690
rect 6644 701626 6696 701632
rect 4434 701312 4490 701321
rect 4434 701247 4490 701256
rect 4066 514791 4122 514800
rect 4344 514820 4396 514826
rect 4344 514762 4396 514768
rect 4448 412634 4476 701247
rect 6656 699938 6684 701626
rect 8128 700330 8156 703520
rect 21456 702500 21508 702506
rect 21456 702442 21508 702448
rect 16302 702400 16358 702409
rect 16302 702335 16358 702344
rect 8116 700324 8168 700330
rect 8116 700266 8168 700272
rect 16316 699938 16344 702335
rect 21468 699938 21496 702442
rect 24320 700398 24348 703520
rect 40512 703390 40540 703520
rect 40500 703384 40552 703390
rect 40500 703326 40552 703332
rect 31206 701584 31262 701593
rect 31206 701519 31262 701528
rect 24308 700392 24360 700398
rect 24308 700334 24360 700340
rect 31220 699938 31248 701519
rect 72988 701010 73016 703520
rect 75460 701956 75512 701962
rect 75460 701898 75512 701904
rect 72976 701004 73028 701010
rect 72976 700946 73028 700952
rect 60646 700088 60702 700097
rect 60646 700023 60702 700032
rect 60660 699938 60688 700023
rect 75472 699938 75500 701898
rect 89180 700670 89208 703520
rect 105464 703458 105492 703520
rect 105452 703452 105504 703458
rect 105452 703394 105504 703400
rect 114284 701888 114336 701894
rect 114284 701830 114336 701836
rect 104808 701752 104860 701758
rect 104808 701694 104860 701700
rect 89168 700664 89220 700670
rect 89168 700606 89220 700612
rect 90178 700360 90234 700369
rect 90178 700295 90234 700304
rect 90192 699938 90220 700295
rect 104820 699938 104848 701694
rect 6440 699910 6684 699938
rect 16192 699910 16344 699938
rect 21160 699910 21496 699938
rect 30912 699910 31248 699938
rect 60444 699910 60688 699938
rect 75164 699910 75500 699938
rect 89884 699910 90220 699938
rect 104604 699910 104848 699938
rect 26146 699816 26202 699825
rect 26036 699774 26146 699802
rect 26146 699751 26202 699760
rect 114296 699666 114324 701830
rect 134432 701412 134484 701418
rect 134432 701354 134484 701360
rect 129464 701344 129516 701350
rect 129464 701286 129516 701292
rect 119712 701208 119764 701214
rect 119712 701150 119764 701156
rect 119724 699938 119752 701150
rect 129476 699938 129504 701286
rect 134444 699938 134472 701354
rect 137848 700942 137876 703520
rect 139308 702840 139360 702846
rect 139308 702782 139360 702788
rect 137836 700936 137888 700942
rect 137836 700878 137888 700884
rect 139320 699938 139348 702782
rect 154028 702092 154080 702098
rect 154028 702034 154080 702040
rect 148968 701616 149020 701622
rect 148968 701558 149020 701564
rect 144276 701480 144328 701486
rect 144276 701422 144328 701428
rect 144288 699938 144316 701422
rect 148980 699938 149008 701558
rect 154040 699938 154068 702034
rect 154132 700874 154160 703520
rect 170324 703474 170352 703520
rect 170508 703474 170536 703666
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 227628 703520 227680 703526
rect 235142 703520 235254 704960
rect 235448 703860 235500 703866
rect 235448 703802 235500 703808
rect 235460 703610 235488 703802
rect 235368 703582 235488 703610
rect 242440 703588 242492 703594
rect 170324 703446 170536 703474
rect 198280 703112 198332 703118
rect 198280 703054 198332 703060
rect 183376 702976 183428 702982
rect 183376 702918 183428 702924
rect 178592 702024 178644 702030
rect 178592 701966 178644 701972
rect 154120 700868 154172 700874
rect 154120 700810 154172 700816
rect 163870 700632 163926 700641
rect 163870 700567 163926 700576
rect 163884 699938 163912 700567
rect 178604 699938 178632 701966
rect 183388 699938 183416 702918
rect 198292 699938 198320 703054
rect 202800 700126 202828 703520
rect 213000 703248 213052 703254
rect 213000 703190 213052 703196
rect 207018 702128 207074 702137
rect 207018 702063 207074 702072
rect 207032 700806 207060 702063
rect 207020 700800 207072 700806
rect 207020 700742 207072 700748
rect 202788 700120 202840 700126
rect 202788 700062 202840 700068
rect 213012 699938 213040 703190
rect 218992 700194 219020 703520
rect 227628 703462 227680 703468
rect 235184 703474 235212 703520
rect 235368 703474 235396 703582
rect 242440 703530 242492 703536
rect 224960 701820 225012 701826
rect 224960 701762 225012 701768
rect 224972 700466 225000 701762
rect 224960 700460 225012 700466
rect 224960 700402 225012 700408
rect 218980 700188 219032 700194
rect 218980 700130 219032 700136
rect 217876 700052 217928 700058
rect 217876 699994 217928 700000
rect 217888 699938 217916 699994
rect 222844 699984 222896 699990
rect 119416 699910 119752 699938
rect 129168 699910 129504 699938
rect 134136 699910 134472 699938
rect 139012 699910 139348 699938
rect 143980 699910 144316 699938
rect 148856 699910 149008 699938
rect 153732 699910 154068 699938
rect 163576 699910 163912 699938
rect 178296 699910 178632 699938
rect 183264 699910 183416 699938
rect 197984 699910 198320 699938
rect 212704 699910 213040 699938
rect 217580 699910 217916 699938
rect 222548 699932 222844 699938
rect 227640 699938 227668 703462
rect 235184 703446 235396 703474
rect 232688 702160 232740 702166
rect 232688 702102 232740 702108
rect 232700 699938 232728 702102
rect 232872 701956 232924 701962
rect 232872 701898 232924 701904
rect 222548 699926 222896 699932
rect 222548 699910 222884 699926
rect 227424 699910 227668 699938
rect 232392 699910 232728 699938
rect 208124 699848 208176 699854
rect 207828 699796 208124 699802
rect 207828 699790 208176 699796
rect 207828 699774 208164 699790
rect 193220 699712 193272 699718
rect 114296 699638 114448 699666
rect 193108 699660 193220 699666
rect 193108 699654 193272 699660
rect 193108 699638 193260 699654
rect 232884 699446 232912 701898
rect 237104 700460 237156 700466
rect 237104 700402 237156 700408
rect 237116 699666 237144 700402
rect 242452 699938 242480 703530
rect 251426 703520 251538 704960
rect 257252 703656 257304 703662
rect 257252 703598 257304 703604
rect 247408 702296 247460 702302
rect 247408 702238 247460 702244
rect 247420 699938 247448 702238
rect 252284 701684 252336 701690
rect 252284 701626 252336 701632
rect 253204 701684 253256 701690
rect 253204 701626 253256 701632
rect 252296 701185 252324 701626
rect 252282 701176 252338 701185
rect 252282 701111 252338 701120
rect 252284 700800 252336 700806
rect 252284 700742 252336 700748
rect 252296 699938 252324 700742
rect 253216 700738 253244 701626
rect 253204 700732 253256 700738
rect 253204 700674 253256 700680
rect 257264 699938 257292 703598
rect 267618 703520 267730 704960
rect 271788 703792 271840 703798
rect 271788 703734 271840 703740
rect 260840 701956 260892 701962
rect 260840 701898 260892 701904
rect 260852 700602 260880 701898
rect 267004 700732 267056 700738
rect 267004 700674 267056 700680
rect 260840 700596 260892 700602
rect 260840 700538 260892 700544
rect 262128 700256 262180 700262
rect 262128 700198 262180 700204
rect 262140 699938 262168 700198
rect 267016 699938 267044 700674
rect 267660 700602 267688 703520
rect 267648 700596 267700 700602
rect 267648 700538 267700 700544
rect 271800 699938 271828 703734
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 300860 703860 300912 703866
rect 300860 703802 300912 703808
rect 276020 702432 276072 702438
rect 283852 702434 283880 703520
rect 283852 702406 284156 702434
rect 276020 702374 276072 702380
rect 276032 700126 276060 702374
rect 280988 702228 281040 702234
rect 280988 702170 281040 702176
rect 277492 701888 277544 701894
rect 277492 701830 277544 701836
rect 276020 700120 276072 700126
rect 276020 700062 276072 700068
rect 276526 700120 276578 700126
rect 276526 700062 276578 700068
rect 242144 699910 242480 699938
rect 247112 699910 247448 699938
rect 251988 699910 252324 699938
rect 256956 699910 257292 699938
rect 261832 699910 262168 699938
rect 266708 699910 267044 699938
rect 271676 699910 271828 699938
rect 276538 699924 276566 700062
rect 237116 699638 237268 699666
rect 277504 699650 277532 701830
rect 281000 700602 281028 702170
rect 282920 701888 282972 701894
rect 282920 701830 282972 701836
rect 282932 700942 282960 701830
rect 284128 700942 284156 702406
rect 291844 702092 291896 702098
rect 291844 702034 291896 702040
rect 286690 701176 286746 701185
rect 286690 701111 286746 701120
rect 282920 700936 282972 700942
rect 282920 700878 282972 700884
rect 284116 700936 284168 700942
rect 284116 700878 284168 700884
rect 280988 700596 281040 700602
rect 280988 700538 281040 700544
rect 281494 700120 281546 700126
rect 281494 700062 281546 700068
rect 281506 699924 281534 700062
rect 286704 699938 286732 701111
rect 291856 700534 291884 702034
rect 298006 701176 298062 701185
rect 298006 701111 298062 701120
rect 298020 700942 298048 701111
rect 300136 700942 300164 703520
rect 295892 700936 295944 700942
rect 295892 700878 295944 700884
rect 298008 700936 298060 700942
rect 298008 700878 298060 700884
rect 300124 700936 300176 700942
rect 300124 700878 300176 700884
rect 291384 700528 291436 700534
rect 291384 700470 291436 700476
rect 291844 700528 291896 700534
rect 291844 700470 291896 700476
rect 286396 699910 286732 699938
rect 291396 699666 291424 700470
rect 295904 699938 295932 700878
rect 300872 699938 300900 703802
rect 315488 703724 315540 703730
rect 315488 703666 315540 703672
rect 305736 702432 305788 702438
rect 305736 702374 305788 702380
rect 305748 699938 305776 702374
rect 313280 702296 313332 702302
rect 313280 702238 313332 702244
rect 313292 700942 313320 702238
rect 313280 700936 313332 700942
rect 313280 700878 313332 700884
rect 310934 700188 310986 700194
rect 310934 700130 310986 700136
rect 295904 699910 296240 699938
rect 300872 699910 301116 699938
rect 305748 699910 306084 699938
rect 310946 699924 310974 700130
rect 315500 699938 315528 703666
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364708 703792 364760 703798
rect 364708 703734 364760 703740
rect 364720 703610 364748 703734
rect 364720 703582 364840 703610
rect 330300 703452 330352 703458
rect 330300 703394 330352 703400
rect 325608 702024 325660 702030
rect 325608 701966 325660 701972
rect 320456 701888 320508 701894
rect 320456 701830 320508 701836
rect 320916 701888 320968 701894
rect 320916 701830 320968 701836
rect 320468 699938 320496 701830
rect 315500 699910 315836 699938
rect 320468 699910 320804 699938
rect 277492 699644 277544 699650
rect 291272 699638 291424 699666
rect 277492 699586 277544 699592
rect 320928 699582 320956 701830
rect 325620 700874 325648 701966
rect 325332 700868 325384 700874
rect 325332 700810 325384 700816
rect 325608 700868 325660 700874
rect 325608 700810 325660 700816
rect 325344 699938 325372 700810
rect 330312 699938 330340 703394
rect 332520 700602 332548 703520
rect 345020 703384 345072 703390
rect 345020 703326 345072 703332
rect 340880 701752 340932 701758
rect 340880 701694 340932 701700
rect 335360 701072 335412 701078
rect 335360 701014 335412 701020
rect 332508 700596 332560 700602
rect 332508 700538 332560 700544
rect 325344 699910 325680 699938
rect 330312 699910 330648 699938
rect 335372 699802 335400 701014
rect 340892 700670 340920 701694
rect 340972 701072 341024 701078
rect 340972 701014 341024 701020
rect 340052 700664 340104 700670
rect 340052 700606 340104 700612
rect 340880 700664 340932 700670
rect 340880 700606 340932 700612
rect 340064 699938 340092 700606
rect 340064 699910 340400 699938
rect 335372 699774 335524 699802
rect 320916 699576 320968 699582
rect 320916 699518 320968 699524
rect 340984 699514 341012 701014
rect 345032 699938 345060 703326
rect 348804 700126 348832 703520
rect 364812 703474 364840 703582
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429660 703656 429712 703662
rect 429660 703598 429712 703604
rect 364996 703474 365024 703520
rect 364812 703446 365024 703474
rect 359740 703316 359792 703322
rect 359740 703258 359792 703264
rect 349804 702160 349856 702166
rect 349804 702102 349856 702108
rect 349816 700602 349844 702102
rect 349804 700596 349856 700602
rect 349804 700538 349856 700544
rect 354956 700392 355008 700398
rect 354956 700334 355008 700340
rect 349896 700324 349948 700330
rect 349896 700266 349948 700272
rect 348792 700120 348844 700126
rect 348792 700062 348844 700068
rect 349908 699938 349936 700266
rect 354968 699938 354996 700334
rect 359752 699938 359780 703258
rect 374460 703180 374512 703186
rect 374460 703122 374512 703128
rect 374472 699938 374500 703122
rect 389180 703044 389232 703050
rect 389180 702986 389232 702992
rect 384304 702228 384356 702234
rect 384304 702170 384356 702176
rect 384316 699938 384344 702170
rect 389192 699938 389220 702986
rect 397472 700262 397500 703520
rect 403900 702908 403952 702914
rect 403900 702850 403952 702856
rect 399024 701956 399076 701962
rect 399024 701898 399076 701904
rect 397460 700256 397512 700262
rect 397460 700198 397512 700204
rect 399036 699938 399064 701898
rect 403912 699938 403940 702850
rect 413664 700738 413692 703520
rect 429672 703474 429700 703598
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494440 703594 494652 703610
rect 494428 703588 494652 703594
rect 494480 703582 494652 703588
rect 494428 703530 494480 703536
rect 429856 703474 429884 703520
rect 429672 703446 429884 703474
rect 448152 702772 448204 702778
rect 448152 702714 448204 702720
rect 414204 701820 414256 701826
rect 414204 701762 414256 701768
rect 413652 700732 413704 700738
rect 413652 700674 413704 700680
rect 345032 699910 345368 699938
rect 349908 699910 350244 699938
rect 354968 699910 355212 699938
rect 359752 699910 360088 699938
rect 364628 699922 364964 699938
rect 364616 699916 364964 699922
rect 364668 699910 364964 699916
rect 374472 699910 374808 699938
rect 384316 699910 384652 699938
rect 389192 699910 389528 699938
rect 399036 699910 399372 699938
rect 403912 699910 404248 699938
rect 364616 699858 364668 699864
rect 369780 699786 369932 699802
rect 369768 699780 369932 699786
rect 369820 699774 369932 699780
rect 369768 699722 369820 699728
rect 414216 699666 414244 701762
rect 428464 701548 428516 701554
rect 428464 701490 428516 701496
rect 428476 699938 428504 701490
rect 443274 700496 443330 700505
rect 443274 700431 443330 700440
rect 443288 699938 443316 700431
rect 448164 699938 448192 702714
rect 453028 701684 453080 701690
rect 453028 701626 453080 701632
rect 453040 699938 453068 701626
rect 458180 701276 458232 701282
rect 458180 701218 458232 701224
rect 458192 699938 458220 701218
rect 462332 700942 462360 703520
rect 477592 702704 477644 702710
rect 477592 702646 477644 702652
rect 472716 702364 472768 702370
rect 472716 702306 472768 702312
rect 467840 701140 467892 701146
rect 467840 701082 467892 701088
rect 462320 700936 462372 700942
rect 462320 700878 462372 700884
rect 467852 699938 467880 701082
rect 472728 699938 472756 702306
rect 477604 699938 477632 702646
rect 478524 700806 478552 703520
rect 494624 703474 494652 703582
rect 494766 703520 494878 704960
rect 503904 703520 503956 703526
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 494808 703474 494836 703520
rect 494624 703446 494836 703474
rect 503904 703462 503956 703468
rect 487434 701992 487490 702001
rect 487434 701927 487490 701936
rect 482560 701888 482612 701894
rect 482560 701830 482612 701836
rect 478512 700800 478564 700806
rect 478512 700742 478564 700748
rect 482572 699938 482600 701830
rect 487448 699938 487476 701927
rect 497278 701856 497334 701865
rect 497278 701791 497334 701800
rect 497292 699938 497320 701791
rect 503916 700942 503944 703462
rect 507124 702636 507176 702642
rect 507124 702578 507176 702584
rect 503904 700936 503956 700942
rect 503904 700878 503956 700884
rect 502476 700224 502532 700233
rect 502476 700159 502532 700168
rect 428476 699910 428812 699938
rect 443288 699910 443624 699938
rect 448164 699910 448500 699938
rect 453040 699910 453376 699938
rect 458192 699910 458344 699938
rect 467852 699910 468188 699938
rect 472728 699910 473064 699938
rect 477604 699910 477940 699938
rect 482572 699910 482908 699938
rect 487448 699910 487784 699938
rect 497292 699910 497628 699938
rect 502490 699924 502518 700159
rect 507136 699938 507164 702578
rect 516966 702128 517022 702137
rect 516966 702063 517022 702072
rect 512000 701072 512052 701078
rect 512000 701014 512052 701020
rect 512012 699938 512040 701014
rect 516980 699938 517008 702063
rect 526718 701720 526774 701729
rect 526718 701655 526774 701664
rect 526732 699938 526760 701655
rect 527192 700602 527220 703520
rect 536840 702568 536892 702574
rect 536840 702510 536892 702516
rect 527180 700596 527232 700602
rect 527180 700538 527232 700544
rect 536852 700210 536880 702510
rect 543476 700466 543504 703520
rect 546498 701448 546554 701457
rect 546498 701383 546554 701392
rect 543464 700460 543516 700466
rect 543464 700402 543516 700408
rect 536852 700182 536926 700210
rect 531686 699952 531742 699961
rect 507136 699910 507472 699938
rect 512012 699910 512348 699938
rect 516980 699910 517316 699938
rect 526732 699910 527068 699938
rect 531742 699910 532036 699938
rect 536898 699924 536926 700182
rect 546512 699938 546540 701383
rect 551282 701312 551338 701321
rect 551282 701247 551338 701256
rect 551296 699938 551324 701247
rect 556896 701072 556948 701078
rect 556896 701014 556948 701020
rect 556908 699938 556936 701014
rect 559668 700942 559696 703520
rect 576400 703248 576452 703254
rect 576400 703190 576452 703196
rect 575020 703112 575072 703118
rect 575020 703054 575072 703060
rect 573640 702976 573692 702982
rect 573640 702918 573692 702924
rect 572168 702840 572220 702846
rect 572168 702782 572220 702788
rect 561126 702264 561182 702273
rect 561126 702199 561182 702208
rect 559656 700936 559708 700942
rect 559656 700878 559708 700884
rect 546512 699910 546756 699938
rect 551296 699910 551632 699938
rect 556600 699910 556936 699938
rect 561140 699938 561168 702199
rect 567844 701616 567896 701622
rect 567844 701558 567896 701564
rect 569222 701584 569278 701593
rect 564440 701072 564492 701078
rect 564440 701014 564492 701020
rect 563520 700052 563572 700058
rect 563520 699994 563572 700000
rect 561140 699910 561476 699938
rect 531686 699887 531742 699896
rect 414092 699638 414244 699666
rect 386234 699544 386290 699553
rect 379532 699514 379776 699530
rect 340972 699508 341024 699514
rect 340972 699450 341024 699456
rect 379520 699508 379776 699514
rect 379572 699502 379776 699508
rect 394160 699514 394496 699530
rect 408880 699514 409216 699530
rect 423692 699514 423936 699530
rect 438320 699514 438656 699530
rect 521856 699514 522192 699530
rect 386234 699479 386236 699488
rect 379520 699450 379572 699456
rect 386288 699479 386290 699488
rect 394148 699508 394496 699514
rect 386236 699450 386288 699456
rect 394200 699502 394496 699508
rect 408868 699508 409216 699514
rect 394148 699450 394200 699456
rect 408920 699502 409216 699508
rect 423680 699508 423936 699514
rect 408868 699450 408920 699456
rect 423732 699502 423936 699508
rect 438308 699508 438656 699514
rect 423680 699450 423732 699456
rect 438360 699502 438656 699508
rect 521844 699508 522192 699514
rect 438308 699450 438360 699456
rect 521896 699502 522192 699508
rect 521844 699450 521896 699456
rect 232872 699440 232924 699446
rect 11610 699408 11666 699417
rect 11316 699366 11610 699394
rect 41050 699408 41106 699417
rect 35880 699378 36032 699394
rect 35880 699372 36044 699378
rect 35880 699366 35992 699372
rect 11610 699343 11666 699352
rect 40756 699366 41050 699394
rect 46018 699408 46074 699417
rect 45724 699366 46018 699394
rect 41050 699343 41106 699352
rect 50894 699408 50950 699417
rect 50600 699366 50894 699394
rect 46018 699343 46074 699352
rect 55770 699408 55826 699417
rect 55476 699366 55770 699394
rect 50894 699343 50950 699352
rect 95146 699408 95202 699417
rect 65320 699378 65656 699394
rect 70288 699378 70440 699394
rect 80040 699378 80192 699394
rect 85008 699378 85344 699394
rect 65320 699372 65668 699378
rect 65320 699366 65616 699372
rect 55770 699343 55826 699352
rect 35992 699314 36044 699320
rect 70288 699372 70452 699378
rect 70288 699366 70400 699372
rect 65616 699314 65668 699320
rect 80040 699372 80204 699378
rect 80040 699366 80152 699372
rect 70400 699314 70452 699320
rect 85008 699372 85356 699378
rect 85008 699366 85304 699372
rect 80152 699314 80204 699320
rect 94852 699366 95146 699394
rect 124586 699408 124642 699417
rect 99728 699378 100064 699394
rect 109572 699378 109908 699394
rect 99728 699372 100076 699378
rect 99728 699366 100024 699372
rect 95146 699343 95202 699352
rect 85304 699314 85356 699320
rect 109572 699372 109920 699378
rect 109572 699366 109868 699372
rect 100024 699314 100076 699320
rect 124292 699366 124586 699394
rect 158700 699378 158852 699394
rect 168544 699378 168880 699394
rect 173420 699378 173756 699394
rect 188140 699378 188476 699394
rect 202860 699378 203012 699394
rect 232872 699382 232924 699388
rect 418710 699408 418766 699417
rect 158700 699372 158864 699378
rect 158700 699366 158812 699372
rect 124586 699343 124642 699352
rect 109868 699314 109920 699320
rect 168544 699372 168892 699378
rect 168544 699366 168840 699372
rect 158812 699314 158864 699320
rect 173420 699372 173768 699378
rect 173420 699366 173716 699372
rect 168840 699314 168892 699320
rect 188140 699372 188488 699378
rect 188140 699366 188436 699372
rect 173716 699314 173768 699320
rect 202860 699372 203024 699378
rect 202860 699366 202972 699372
rect 188436 699314 188488 699320
rect 433430 699408 433486 699417
rect 418766 699366 419060 699394
rect 418710 699343 418766 699352
rect 462870 699408 462926 699417
rect 433486 699366 433780 699394
rect 433430 699343 433486 699352
rect 492586 699408 492642 699417
rect 462926 699366 463220 699394
rect 462870 699343 462926 699352
rect 541530 699408 541586 699417
rect 492642 699366 492752 699394
rect 492586 699343 492642 699352
rect 541586 699366 541880 699394
rect 541530 699343 541586 699352
rect 202972 699314 203024 699320
rect 563532 698290 563560 699994
rect 563520 698284 563572 698290
rect 563520 698226 563572 698232
rect 4172 412606 4476 412634
rect 4172 409986 4200 412606
rect 4080 409958 4200 409986
rect 3974 241088 4030 241097
rect 3974 241023 4030 241032
rect 3882 201920 3938 201929
rect 3882 201855 3938 201864
rect 3790 149832 3846 149841
rect 3790 149767 3846 149776
rect 3698 136776 3754 136785
rect 3698 136711 3754 136720
rect 3606 97608 3662 97617
rect 3606 97543 3662 97552
rect 3514 45520 3570 45529
rect 3514 45455 3570 45464
rect 4080 32473 4108 409958
rect 4066 32464 4122 32473
rect 4066 32399 4122 32408
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 2962 6488 3018 6497
rect 2962 6423 3018 6432
rect 2976 2106 3004 6423
rect 563704 3052 563756 3058
rect 563704 2994 563756 3000
rect 563520 2984 563572 2990
rect 563520 2926 563572 2932
rect 2964 2100 3016 2106
rect 2964 2042 3016 2048
rect 563532 1086 563560 2926
rect 563612 2916 563664 2922
rect 563612 2858 563664 2864
rect 563624 1154 563652 2858
rect 563612 1148 563664 1154
rect 563612 1090 563664 1096
rect 563520 1080 563572 1086
rect 563520 1022 563572 1028
rect 563716 762 563744 2994
rect 564452 2106 564480 701014
rect 565082 699816 565138 699825
rect 565082 699751 565138 699760
rect 565096 73166 565124 699751
rect 565360 699100 565412 699106
rect 565360 699042 565412 699048
rect 565174 698864 565230 698873
rect 565174 698799 565230 698808
rect 565188 126954 565216 698799
rect 565266 697776 565322 697785
rect 565266 697711 565322 697720
rect 565280 245614 565308 697711
rect 565372 511970 565400 699042
rect 566646 698592 566702 698601
rect 566646 698527 566702 698536
rect 566556 698352 566608 698358
rect 566462 698320 566518 698329
rect 566556 698294 566608 698300
rect 566462 698255 566518 698264
rect 565360 511964 565412 511970
rect 565360 511906 565412 511912
rect 565268 245608 565320 245614
rect 565268 245550 565320 245556
rect 565176 126948 565228 126954
rect 565176 126890 565228 126896
rect 565084 73160 565136 73166
rect 565084 73102 565136 73108
rect 566476 33114 566504 698255
rect 566568 167006 566596 698294
rect 566556 167000 566608 167006
rect 566556 166942 566608 166948
rect 566660 113150 566688 698527
rect 566740 698488 566792 698494
rect 566740 698430 566792 698436
rect 566752 206990 566780 698430
rect 567856 419490 567884 701558
rect 569222 701519 569278 701528
rect 567844 419484 567896 419490
rect 567844 419426 567896 419432
rect 566740 206984 566792 206990
rect 566740 206926 566792 206932
rect 566648 113144 566700 113150
rect 566648 113086 566700 113092
rect 569236 60722 569264 701519
rect 570694 700088 570750 700097
rect 570694 700023 570750 700032
rect 569592 699236 569644 699242
rect 569592 699178 569644 699184
rect 569314 699000 569370 699009
rect 569314 698935 569370 698944
rect 569328 153202 569356 698935
rect 569500 698692 569552 698698
rect 569500 698634 569552 698640
rect 569408 698420 569460 698426
rect 569408 698362 569460 698368
rect 569420 193186 569448 698362
rect 569512 299470 569540 698634
rect 569604 592006 569632 699178
rect 570602 698728 570658 698737
rect 570602 698663 570658 698672
rect 569592 592000 569644 592006
rect 569592 591942 569644 591948
rect 569500 299464 569552 299470
rect 569500 299406 569552 299412
rect 569408 193180 569460 193186
rect 569408 193122 569460 193128
rect 569316 153196 569368 153202
rect 569316 153138 569368 153144
rect 570616 100706 570644 698663
rect 570708 139398 570736 700023
rect 570880 699848 570932 699854
rect 570880 699790 570932 699796
rect 570786 698048 570842 698057
rect 570786 697983 570842 697992
rect 570800 353258 570828 697983
rect 570892 632058 570920 699790
rect 572076 698624 572128 698630
rect 572076 698566 572128 698572
rect 571984 698556 572036 698562
rect 571984 698498 572036 698504
rect 570880 632052 570932 632058
rect 570880 631994 570932 632000
rect 570788 353252 570840 353258
rect 570788 353194 570840 353200
rect 571996 233238 572024 698498
rect 572088 273222 572116 698566
rect 572180 405686 572208 702782
rect 573456 701344 573508 701350
rect 573456 701286 573508 701292
rect 573362 700360 573418 700369
rect 573362 700295 573418 700304
rect 572168 405680 572220 405686
rect 572168 405622 572220 405628
rect 572076 273216 572128 273222
rect 572076 273158 572128 273164
rect 571984 233232 572036 233238
rect 571984 233174 572036 233180
rect 573376 219434 573404 700295
rect 573468 379506 573496 701286
rect 573548 699032 573600 699038
rect 573548 698974 573600 698980
rect 573560 538218 573588 698974
rect 573652 564398 573680 702918
rect 574928 701480 574980 701486
rect 574928 701422 574980 701428
rect 574836 701208 574888 701214
rect 574836 701150 574888 701156
rect 573732 699372 573784 699378
rect 573732 699314 573784 699320
rect 573744 644434 573772 699314
rect 574744 697604 574796 697610
rect 574744 697546 574796 697552
rect 573732 644428 573784 644434
rect 573732 644370 573784 644376
rect 573640 564392 573692 564398
rect 573640 564334 573692 564340
rect 573548 538212 573600 538218
rect 573548 538154 573600 538160
rect 573456 379500 573508 379506
rect 573456 379442 573508 379448
rect 573364 219428 573416 219434
rect 573364 219370 573416 219376
rect 570696 139392 570748 139398
rect 570696 139334 570748 139340
rect 570604 100700 570656 100706
rect 570604 100642 570656 100648
rect 574756 86970 574784 697546
rect 574848 313274 574876 701150
rect 574940 431934 574968 701422
rect 575032 618254 575060 703054
rect 576124 702500 576176 702506
rect 576124 702442 576176 702448
rect 575020 618248 575072 618254
rect 575020 618190 575072 618196
rect 574928 431928 574980 431934
rect 574928 431870 574980 431876
rect 574836 313268 574888 313274
rect 574836 313210 574888 313216
rect 574744 86964 574796 86970
rect 574744 86906 574796 86912
rect 569224 60716 569276 60722
rect 569224 60658 569276 60664
rect 576136 46918 576164 702442
rect 576216 701412 576268 701418
rect 576216 701354 576268 701360
rect 576228 365702 576256 701354
rect 576306 700632 576362 700641
rect 576306 700567 576362 700576
rect 576320 471986 576348 700567
rect 576412 672042 576440 703190
rect 577502 702400 577558 702409
rect 577502 702335 577558 702344
rect 576400 672036 576452 672042
rect 576400 671978 576452 671984
rect 576308 471980 576360 471986
rect 576308 471922 576360 471928
rect 576216 365696 576268 365702
rect 576216 365638 576268 365644
rect 576124 46912 576176 46918
rect 576124 46854 576176 46860
rect 566464 33108 566516 33114
rect 566464 33050 566516 33056
rect 577516 20670 577544 702335
rect 580724 700868 580776 700874
rect 580724 700810 580776 700816
rect 580448 700664 580500 700670
rect 580448 700606 580500 700612
rect 579068 699984 579120 699990
rect 579068 699926 579120 699932
rect 578976 699712 579028 699718
rect 578976 699654 579028 699660
rect 578884 698896 578936 698902
rect 578884 698838 578936 698844
rect 578896 484673 578924 698838
rect 578988 577697 579016 699654
rect 579080 683913 579108 699926
rect 580356 699440 580408 699446
rect 580356 699382 580408 699388
rect 580262 699136 580318 699145
rect 580262 699071 580318 699080
rect 580172 698284 580224 698290
rect 580172 698226 580224 698232
rect 580184 697241 580212 698226
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 579066 683904 579122 683913
rect 579066 683839 579122 683848
rect 579620 672036 579672 672042
rect 579620 671978 579672 671984
rect 579632 670721 579660 671978
rect 579618 670712 579674 670721
rect 579618 670647 579674 670656
rect 580172 644428 580224 644434
rect 580172 644370 580224 644376
rect 580184 644065 580212 644370
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580172 632052 580224 632058
rect 580172 631994 580224 632000
rect 580184 630873 580212 631994
rect 580170 630864 580226 630873
rect 580170 630799 580226 630808
rect 580172 618248 580224 618254
rect 580172 618190 580224 618196
rect 580184 617545 580212 618190
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580172 592000 580224 592006
rect 580172 591942 580224 591948
rect 580184 591025 580212 591942
rect 580170 591016 580226 591025
rect 580170 590951 580226 590960
rect 578974 577688 579030 577697
rect 578974 577623 579030 577632
rect 580172 564392 580224 564398
rect 580170 564360 580172 564369
rect 580224 564360 580226 564369
rect 580170 564295 580226 564304
rect 580172 538212 580224 538218
rect 580172 538154 580224 538160
rect 580184 537849 580212 538154
rect 580170 537840 580226 537849
rect 580170 537775 580226 537784
rect 580172 511964 580224 511970
rect 580172 511906 580224 511912
rect 580184 511329 580212 511906
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 578882 484664 578938 484673
rect 578882 484599 578938 484608
rect 579804 471980 579856 471986
rect 579804 471922 579856 471928
rect 579816 471481 579844 471922
rect 579802 471472 579858 471481
rect 579802 471407 579858 471416
rect 579712 431928 579764 431934
rect 579712 431870 579764 431876
rect 579724 431633 579752 431870
rect 579710 431624 579766 431633
rect 579710 431559 579766 431568
rect 580172 419484 580224 419490
rect 580172 419426 580224 419432
rect 580184 418305 580212 419426
rect 580170 418296 580226 418305
rect 580170 418231 580226 418240
rect 580172 405680 580224 405686
rect 580172 405622 580224 405628
rect 580184 404977 580212 405622
rect 580170 404968 580226 404977
rect 580170 404903 580226 404912
rect 579620 379500 579672 379506
rect 579620 379442 579672 379448
rect 579632 378457 579660 379442
rect 579618 378448 579674 378457
rect 579618 378383 579674 378392
rect 580172 365696 580224 365702
rect 580172 365638 580224 365644
rect 580184 365129 580212 365638
rect 580170 365120 580226 365129
rect 580170 365055 580226 365064
rect 580172 353252 580224 353258
rect 580172 353194 580224 353200
rect 580184 351937 580212 353194
rect 580170 351928 580226 351937
rect 580170 351863 580226 351872
rect 579712 313268 579764 313274
rect 579712 313210 579764 313216
rect 579724 312089 579752 313210
rect 579710 312080 579766 312089
rect 579710 312015 579766 312024
rect 579804 299464 579856 299470
rect 579804 299406 579856 299412
rect 579816 298761 579844 299406
rect 579802 298752 579858 298761
rect 579802 298687 579858 298696
rect 580172 273216 580224 273222
rect 580172 273158 580224 273164
rect 580184 272241 580212 273158
rect 580170 272232 580226 272241
rect 580170 272167 580226 272176
rect 580172 245608 580224 245614
rect 580170 245576 580172 245585
rect 580224 245576 580226 245585
rect 580170 245511 580226 245520
rect 580172 233232 580224 233238
rect 580172 233174 580224 233180
rect 580184 232393 580212 233174
rect 580170 232384 580226 232393
rect 580170 232319 580226 232328
rect 580172 219428 580224 219434
rect 580172 219370 580224 219376
rect 580184 219065 580212 219370
rect 580170 219056 580226 219065
rect 580170 218991 580226 219000
rect 579896 206984 579948 206990
rect 579896 206926 579948 206932
rect 579908 205737 579936 206926
rect 579894 205728 579950 205737
rect 579894 205663 579950 205672
rect 580172 193180 580224 193186
rect 580172 193122 580224 193128
rect 580184 192545 580212 193122
rect 580170 192536 580226 192545
rect 580170 192471 580226 192480
rect 580172 167000 580224 167006
rect 580172 166942 580224 166948
rect 580184 165889 580212 166942
rect 580170 165880 580226 165889
rect 580170 165815 580226 165824
rect 579804 153196 579856 153202
rect 579804 153138 579856 153144
rect 579816 152697 579844 153138
rect 579802 152688 579858 152697
rect 579802 152623 579858 152632
rect 580172 139392 580224 139398
rect 580170 139360 580172 139369
rect 580224 139360 580226 139369
rect 580170 139295 580226 139304
rect 580172 126948 580224 126954
rect 580172 126890 580224 126896
rect 580184 126041 580212 126890
rect 580170 126032 580226 126041
rect 580170 125967 580226 125976
rect 580172 113144 580224 113150
rect 580172 113086 580224 113092
rect 580184 112849 580212 113086
rect 580170 112840 580226 112849
rect 580170 112775 580226 112784
rect 580172 100700 580224 100706
rect 580172 100642 580224 100648
rect 580184 99521 580212 100642
rect 580170 99512 580226 99521
rect 580170 99447 580226 99456
rect 580172 86964 580224 86970
rect 580172 86906 580224 86912
rect 580184 86193 580212 86906
rect 580170 86184 580226 86193
rect 580170 86119 580226 86128
rect 579988 73160 580040 73166
rect 579988 73102 580040 73108
rect 580000 73001 580028 73102
rect 579986 72992 580042 73001
rect 579986 72927 580042 72936
rect 580172 60716 580224 60722
rect 580172 60658 580224 60664
rect 580184 59673 580212 60658
rect 580170 59664 580226 59673
rect 580170 59599 580226 59608
rect 580172 46912 580224 46918
rect 580172 46854 580224 46860
rect 580184 46345 580212 46854
rect 580170 46336 580226 46345
rect 580170 46271 580226 46280
rect 580170 33144 580226 33153
rect 580170 33079 580172 33088
rect 580224 33079 580226 33088
rect 580172 33050 580224 33056
rect 577504 20664 577556 20670
rect 577504 20606 577556 20612
rect 579712 20664 579764 20670
rect 579712 20606 579764 20612
rect 579724 19825 579752 20606
rect 579710 19816 579766 19825
rect 579710 19751 579766 19760
rect 580276 6633 580304 699071
rect 580368 179217 580396 699382
rect 580460 258913 580488 700606
rect 580632 700528 580684 700534
rect 580632 700470 580684 700476
rect 580540 699644 580592 699650
rect 580540 699586 580592 699592
rect 580552 325281 580580 699586
rect 580644 458153 580672 700470
rect 580736 524521 580764 700810
rect 580722 524512 580778 524521
rect 580722 524447 580778 524456
rect 580630 458144 580686 458153
rect 580630 458079 580686 458088
rect 580538 325272 580594 325281
rect 580538 325207 580594 325216
rect 580446 258904 580502 258913
rect 580446 258839 580502 258848
rect 580354 179208 580410 179217
rect 580354 179143 580410 179152
rect 580262 6624 580318 6633
rect 580262 6559 580318 6568
rect 569868 3120 569920 3126
rect 569868 3062 569920 3068
rect 577412 3120 577464 3126
rect 577412 3062 577464 3068
rect 564440 2100 564492 2106
rect 564440 2042 564492 2048
rect 565912 1420 565964 1426
rect 565912 1362 565964 1368
rect 569132 1420 569184 1426
rect 569132 1362 569184 1368
rect 565924 882 565952 1362
rect 566832 1216 566884 1222
rect 566832 1158 566884 1164
rect 565912 876 565964 882
rect 565912 818 565964 824
rect 4068 740 4120 746
rect 563408 734 563744 762
rect 565820 808 565872 814
rect 565820 750 565872 756
rect 4068 682 4120 688
rect 1676 672 1728 678
rect 1676 614 1728 620
rect 572 604 624 610
rect 572 546 624 552
rect 584 480 612 546
rect 1688 480 1716 614
rect 2884 598 3096 626
rect 2884 480 2912 598
rect 3068 490 3096 598
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 3068 474 3280 490
rect 4080 480 4108 682
rect 5356 672 5408 678
rect 4264 610 4600 626
rect 7748 672 7800 678
rect 5408 620 5704 626
rect 5356 614 5704 620
rect 11060 672 11112 678
rect 8758 640 8814 649
rect 7800 620 8004 626
rect 7748 614 8004 620
rect 4252 604 4600 610
rect 4304 598 4600 604
rect 5264 604 5316 610
rect 4252 546 4304 552
rect 5368 598 5704 614
rect 6460 604 6512 610
rect 5264 546 5316 552
rect 6460 546 6512 552
rect 7656 604 7708 610
rect 7760 598 8004 614
rect 8758 575 8814 584
rect 9954 640 10010 649
rect 14464 672 14516 678
rect 13266 640 13322 649
rect 11112 620 11192 626
rect 11060 614 11192 620
rect 11072 598 11192 614
rect 9954 575 10010 584
rect 7656 546 7708 552
rect 5276 480 5304 546
rect 6472 480 6500 546
rect 3068 468 3292 474
rect 3068 462 3240 468
rect 3240 410 3292 416
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 6656 474 6808 490
rect 7668 480 7696 546
rect 8772 480 8800 575
rect 9968 480 9996 575
rect 10324 536 10376 542
rect 10212 484 10324 490
rect 6644 468 6808 474
rect 6696 462 6808 468
rect 6644 410 6696 416
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 8944 400 8996 406
rect 8996 348 9108 354
rect 8944 342 9108 348
rect 8956 326 9108 342
rect 9926 -960 10038 480
rect 10212 478 10376 484
rect 11164 480 11192 598
rect 12348 604 12400 610
rect 13322 598 13616 626
rect 19432 672 19484 678
rect 14516 620 14812 626
rect 14464 614 14812 620
rect 14476 598 14812 614
rect 15580 610 15916 626
rect 15568 604 15916 610
rect 13266 575 13322 584
rect 12348 546 12400 552
rect 15620 598 15916 604
rect 16684 598 17020 626
rect 17880 598 18216 626
rect 22376 672 22428 678
rect 19432 614 19484 620
rect 20626 640 20682 649
rect 18512 604 18564 610
rect 15568 546 15620 552
rect 11520 536 11572 542
rect 11408 484 11520 490
rect 10212 462 10364 478
rect 11122 -960 11234 480
rect 11408 478 11572 484
rect 12360 480 12388 546
rect 16684 542 16712 598
rect 13360 536 13412 542
rect 12622 504 12678 513
rect 11408 462 11560 478
rect 12318 -960 12430 480
rect 12512 462 12622 490
rect 13360 478 13412 484
rect 16672 536 16724 542
rect 12622 439 12678 448
rect 13372 354 13400 478
rect 13514 354 13626 480
rect 13372 326 13626 354
rect 14556 400 14608 406
rect 14710 354 14822 480
rect 14608 348 14822 354
rect 14556 342 14822 348
rect 14568 326 14822 342
rect 13514 -960 13626 326
rect 14710 -960 14822 326
rect 15906 82 16018 480
rect 16672 478 16724 484
rect 17010 82 17122 480
rect 17880 406 17908 598
rect 18512 546 18564 552
rect 17868 400 17920 406
rect 17868 342 17920 348
rect 18206 218 18318 480
rect 18524 218 18552 546
rect 19444 480 19472 614
rect 21284 610 21620 626
rect 23020 672 23072 678
rect 22428 620 22724 626
rect 22376 614 22724 620
rect 25780 672 25832 678
rect 23020 614 23072 620
rect 23478 640 23534 649
rect 20626 575 20682 584
rect 21272 604 21620 610
rect 20640 480 20668 575
rect 21324 598 21620 604
rect 21824 604 21876 610
rect 21272 546 21324 552
rect 22388 598 22724 614
rect 21824 546 21876 552
rect 21836 480 21864 546
rect 23032 480 23060 614
rect 23534 598 23828 626
rect 24872 610 25024 626
rect 28816 672 28868 678
rect 26514 640 26570 649
rect 25832 620 26128 626
rect 25780 614 26128 620
rect 24860 604 25024 610
rect 23478 575 23534 584
rect 24228 564 24440 592
rect 24228 480 24256 564
rect 24412 490 24440 564
rect 24912 598 25024 604
rect 25320 604 25372 610
rect 24860 546 24912 552
rect 25792 598 26128 614
rect 28722 640 28778 649
rect 28092 610 28428 626
rect 28080 604 28428 610
rect 26514 575 26570 584
rect 25320 546 25372 552
rect 18206 190 18552 218
rect 17408 128 17460 134
rect 15906 66 16344 82
rect 17010 76 17408 82
rect 17010 70 17460 76
rect 15906 60 16356 66
rect 15906 54 16304 60
rect 15906 -960 16018 54
rect 16304 2 16356 8
rect 17010 54 17448 70
rect 17010 -960 17122 54
rect 18206 -960 18318 190
rect 18984 66 19320 82
rect 18972 60 19320 66
rect 19024 54 19320 60
rect 18972 2 19024 8
rect 19402 -960 19514 480
rect 20076 128 20128 134
rect 20128 76 20424 82
rect 20076 70 20424 76
rect 20088 54 20424 70
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 24412 474 24900 490
rect 25332 480 25360 546
rect 26528 480 26556 575
rect 27724 564 27936 592
rect 24412 468 24912 474
rect 24412 462 24860 468
rect 24860 410 24912 416
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 26896 474 27232 490
rect 27724 480 27752 564
rect 27908 513 27936 564
rect 28132 598 28428 604
rect 31668 672 31720 678
rect 30286 640 30342 649
rect 28868 620 28948 626
rect 28816 614 28948 620
rect 28828 598 28948 614
rect 29196 610 29532 626
rect 28722 575 28724 584
rect 28080 546 28132 552
rect 28776 575 28778 584
rect 28724 546 28776 552
rect 27894 504 27950 513
rect 26884 468 27232 474
rect 26936 462 27232 468
rect 26884 410 26936 416
rect 27682 -960 27794 480
rect 28920 480 28948 598
rect 29184 604 29532 610
rect 29236 598 29532 604
rect 30104 604 30156 610
rect 29184 546 29236 552
rect 30342 598 30636 626
rect 31312 598 31524 626
rect 32404 672 32456 678
rect 31720 620 31832 626
rect 31668 614 31832 620
rect 34888 672 34940 678
rect 34794 640 34850 649
rect 32404 614 32456 620
rect 31680 598 31832 614
rect 30286 575 30342 584
rect 30104 546 30156 552
rect 30116 480 30144 546
rect 31312 480 31340 598
rect 31496 542 31524 598
rect 31484 536 31536 542
rect 27894 439 27950 448
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 31484 478 31536 484
rect 32416 480 32444 614
rect 32600 610 32936 626
rect 32588 604 32936 610
rect 32640 598 32936 604
rect 33600 604 33652 610
rect 32588 546 32640 552
rect 38384 672 38436 678
rect 35990 640 36046 649
rect 34940 620 35236 626
rect 34888 614 35236 620
rect 34900 598 35236 614
rect 34794 575 34850 584
rect 36096 610 36340 626
rect 40684 672 40736 678
rect 38384 614 38436 620
rect 38474 640 38530 649
rect 35990 575 36046 584
rect 36084 604 36340 610
rect 33600 546 33652 552
rect 33612 480 33640 546
rect 33784 536 33836 542
rect 33836 484 34132 490
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 33784 478 34132 484
rect 34808 480 34836 575
rect 36004 480 36032 575
rect 36136 598 36340 604
rect 37188 604 37240 610
rect 36084 546 36136 552
rect 37188 546 37240 552
rect 37200 480 37228 546
rect 37370 504 37426 513
rect 33796 462 34132 478
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 37426 462 37536 490
rect 38396 480 38424 614
rect 38530 598 38640 626
rect 42800 672 42852 678
rect 40684 614 40736 620
rect 39580 604 39632 610
rect 38474 575 38530 584
rect 39580 546 39632 552
rect 39592 480 39620 546
rect 40696 480 40724 614
rect 40788 610 40940 626
rect 46664 672 46716 678
rect 42852 620 43148 626
rect 42800 614 43148 620
rect 40776 604 40940 610
rect 40828 598 40940 604
rect 41880 604 41932 610
rect 40776 546 40828 552
rect 42812 598 43148 614
rect 44008 610 44344 626
rect 43996 604 44344 610
rect 41880 546 41932 552
rect 44048 598 44344 604
rect 45112 598 45448 626
rect 46664 614 46716 620
rect 48504 672 48556 678
rect 48964 672 49016 678
rect 48556 620 48852 626
rect 48504 614 48852 620
rect 50804 672 50856 678
rect 48964 614 49016 620
rect 43996 546 44048 552
rect 41892 480 41920 546
rect 37370 439 37426 448
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 39856 400 39908 406
rect 39744 348 39856 354
rect 39744 342 39908 348
rect 39744 326 39896 342
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 42044 474 42196 490
rect 42044 468 42208 474
rect 42044 462 42156 468
rect 42156 410 42208 416
rect 42892 400 42944 406
rect 43046 354 43158 480
rect 42944 348 43158 354
rect 42892 342 43158 348
rect 42904 326 43158 342
rect 43046 -960 43158 326
rect 44242 82 44354 480
rect 45112 406 45140 598
rect 46676 480 46704 614
rect 47860 604 47912 610
rect 48516 598 48852 614
rect 47860 546 47912 552
rect 47872 480 47900 546
rect 48976 480 49004 614
rect 49620 610 49956 626
rect 63224 672 63276 678
rect 52550 640 52606 649
rect 50856 620 51152 626
rect 50804 614 51152 620
rect 49608 604 49956 610
rect 49660 598 49956 604
rect 50160 604 50212 610
rect 49608 546 49660 552
rect 50816 598 51152 614
rect 51356 604 51408 610
rect 50160 546 50212 552
rect 54206 640 54262 649
rect 53024 610 53360 626
rect 52550 575 52606 584
rect 53012 604 53360 610
rect 51356 546 51408 552
rect 50172 480 50200 546
rect 51368 480 51396 546
rect 51908 536 51960 542
rect 51960 484 52256 490
rect 45100 400 45152 406
rect 45100 342 45152 348
rect 44100 66 44354 82
rect 44088 60 44354 66
rect 44140 54 44354 60
rect 44088 2 44140 8
rect 44242 -960 44354 54
rect 45438 82 45550 480
rect 45744 128 45796 134
rect 45438 76 45744 82
rect 45438 70 45796 76
rect 45438 54 45784 70
rect 46216 66 46552 82
rect 46204 60 46552 66
rect 45438 -960 45550 54
rect 46256 54 46552 60
rect 46204 2 46256 8
rect 46634 -960 46746 480
rect 47400 128 47452 134
rect 47452 76 47748 82
rect 47400 70 47748 76
rect 47412 54 47748 70
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 51908 478 52256 484
rect 52564 480 52592 575
rect 53064 598 53360 604
rect 53576 598 53788 626
rect 53012 546 53064 552
rect 53576 513 53604 598
rect 53562 504 53618 513
rect 51920 462 52256 478
rect 52522 -960 52634 480
rect 53760 480 53788 598
rect 56046 640 56102 649
rect 54262 598 54556 626
rect 54944 604 54996 610
rect 54206 575 54262 584
rect 57610 640 57666 649
rect 56428 610 56764 626
rect 56046 575 56102 584
rect 56416 604 56764 610
rect 54944 546 54996 552
rect 54956 480 54984 546
rect 55310 504 55366 513
rect 53562 439 53618 448
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 55366 462 55660 490
rect 56060 480 56088 575
rect 56468 598 56764 604
rect 56416 546 56468 552
rect 57256 564 57468 592
rect 58438 640 58494 649
rect 57666 598 57960 626
rect 57610 575 57666 584
rect 59818 640 59874 649
rect 58438 575 58494 584
rect 57256 480 57284 564
rect 57440 513 57468 564
rect 57426 504 57482 513
rect 55310 439 55366 448
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58452 480 58480 575
rect 59464 564 59676 592
rect 60830 640 60886 649
rect 59874 598 60168 626
rect 59818 575 59874 584
rect 62118 640 62174 649
rect 60830 575 60886 584
rect 62028 604 62080 610
rect 59464 513 59492 564
rect 58806 504 58862 513
rect 57426 439 57482 448
rect 58410 -960 58522 480
rect 59450 504 59506 513
rect 58862 462 59064 490
rect 58806 439 58862 448
rect 59648 480 59676 564
rect 60844 480 60872 575
rect 62174 598 62468 626
rect 64328 672 64380 678
rect 63224 614 63276 620
rect 62118 575 62174 584
rect 62028 546 62080 552
rect 61106 504 61162 513
rect 59450 439 59506 448
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61162 462 61364 490
rect 62040 480 62068 546
rect 63236 480 63264 614
rect 63328 610 63664 626
rect 65616 672 65668 678
rect 64328 614 64380 620
rect 63316 604 63664 610
rect 63368 598 63664 604
rect 63316 546 63368 552
rect 64340 480 64368 614
rect 64432 610 64768 626
rect 66720 672 66772 678
rect 65668 620 65872 626
rect 65616 614 65872 620
rect 68008 672 68060 678
rect 66720 614 66772 620
rect 64420 604 64768 610
rect 64472 598 64768 604
rect 65524 604 65576 610
rect 64420 546 64472 552
rect 65628 598 65872 614
rect 65524 546 65576 552
rect 65536 480 65564 546
rect 66732 480 66760 614
rect 66824 610 67068 626
rect 66812 604 67068 610
rect 66864 598 67068 604
rect 67744 598 67956 626
rect 69112 672 69164 678
rect 68060 620 68172 626
rect 68008 614 68172 620
rect 70584 672 70636 678
rect 69112 614 69164 620
rect 70472 620 70584 626
rect 133236 672 133288 678
rect 70472 614 70636 620
rect 68020 598 68172 614
rect 66812 546 66864 552
rect 67744 542 67772 598
rect 67732 536 67784 542
rect 61106 439 61162 448
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67732 478 67784 484
rect 67928 480 67956 598
rect 69124 480 69152 614
rect 70308 604 70360 610
rect 70472 598 70624 614
rect 71240 610 71576 626
rect 71228 604 71576 610
rect 70308 546 70360 552
rect 71280 598 71576 604
rect 72344 598 72680 626
rect 73540 598 73876 626
rect 74644 598 74980 626
rect 76944 610 77280 626
rect 78048 610 78384 626
rect 79152 610 79488 626
rect 80348 610 80684 626
rect 81452 610 81788 626
rect 82740 610 82892 626
rect 76196 604 76248 610
rect 71228 546 71280 552
rect 69388 536 69440 542
rect 69276 484 69388 490
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 69276 478 69440 484
rect 70320 480 70348 546
rect 69276 462 69428 478
rect 70278 -960 70390 480
rect 71320 400 71372 406
rect 71474 354 71586 480
rect 72344 406 72372 598
rect 71372 348 71586 354
rect 71320 342 71586 348
rect 72332 400 72384 406
rect 72332 342 72384 348
rect 72424 400 72476 406
rect 72578 354 72690 480
rect 73540 406 73568 598
rect 72476 348 72690 354
rect 72424 342 72690 348
rect 73528 400 73580 406
rect 73528 342 73580 348
rect 73620 400 73672 406
rect 73774 354 73886 480
rect 74644 406 74672 598
rect 76196 546 76248 552
rect 76932 604 77280 610
rect 76984 598 77280 604
rect 77392 604 77444 610
rect 76932 546 76984 552
rect 77392 546 77444 552
rect 78036 604 78384 610
rect 78088 598 78384 604
rect 78588 604 78640 610
rect 78036 546 78088 552
rect 78588 546 78640 552
rect 79140 604 79488 610
rect 79192 598 79488 604
rect 79692 604 79744 610
rect 79140 546 79192 552
rect 79692 546 79744 552
rect 80336 604 80684 610
rect 80388 598 80684 604
rect 80888 604 80940 610
rect 80336 546 80388 552
rect 80888 546 80940 552
rect 81440 604 81788 610
rect 81492 598 81788 604
rect 82084 604 82136 610
rect 81440 546 81492 552
rect 82084 546 82136 552
rect 82728 604 82892 610
rect 82780 598 82892 604
rect 83292 598 83504 626
rect 82728 546 82780 552
rect 76208 480 76236 546
rect 77404 480 77432 546
rect 78600 480 78628 546
rect 79704 480 79732 546
rect 80900 480 80928 546
rect 82096 480 82124 546
rect 83292 480 83320 598
rect 83476 490 83504 598
rect 84488 598 85192 626
rect 85684 598 85896 626
rect 73672 348 73886 354
rect 73620 342 73886 348
rect 74632 400 74684 406
rect 74632 342 74684 348
rect 71332 326 71586 342
rect 72436 326 72690 342
rect 73632 326 73886 342
rect 71474 -960 71586 326
rect 72578 -960 72690 326
rect 73774 -960 73886 326
rect 74970 82 75082 480
rect 74970 54 76084 82
rect 74970 -960 75082 54
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 83476 462 84088 490
rect 84488 480 84516 598
rect 85684 480 85712 598
rect 85868 490 85896 598
rect 86880 598 87492 626
rect 87984 598 88596 626
rect 89180 598 89392 626
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 85868 462 86296 490
rect 86880 480 86908 598
rect 87984 480 88012 598
rect 89180 480 89208 598
rect 89364 490 89392 598
rect 90376 598 90896 626
rect 91572 598 92000 626
rect 92768 598 93196 626
rect 93964 598 94300 626
rect 95160 598 95404 626
rect 96264 598 96600 626
rect 97460 598 97704 626
rect 98656 598 98808 626
rect 99852 598 100004 626
rect 105616 598 105768 626
rect 106812 598 106964 626
rect 107916 598 108160 626
rect 109020 598 109356 626
rect 110216 598 110552 626
rect 111320 598 111656 626
rect 112424 598 112852 626
rect 113620 598 114048 626
rect 114724 598 115244 626
rect 115828 598 116440 626
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 89364 462 89792 490
rect 90376 480 90404 598
rect 91572 480 91600 598
rect 92768 480 92796 598
rect 93964 480 93992 598
rect 95160 480 95188 598
rect 96264 480 96292 598
rect 97460 480 97488 598
rect 98656 480 98684 598
rect 99852 480 99880 598
rect 105740 480 105768 598
rect 106936 480 106964 598
rect 108132 480 108160 598
rect 109328 480 109356 598
rect 110524 480 110552 598
rect 111628 480 111656 598
rect 112824 480 112852 598
rect 114020 480 114048 598
rect 115216 480 115244 598
rect 116412 480 116440 598
rect 117424 598 117636 626
rect 118128 598 118832 626
rect 119324 598 119936 626
rect 117424 490 117452 598
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117024 462 117452 490
rect 117608 480 117636 598
rect 118804 480 118832 598
rect 119908 480 119936 598
rect 120920 598 121132 626
rect 121532 610 121868 626
rect 121532 604 121880 610
rect 121532 598 121828 604
rect 120920 490 120948 598
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 120428 462 120948 490
rect 121104 480 121132 598
rect 121828 546 121880 552
rect 122288 604 122340 610
rect 122288 546 122340 552
rect 123312 598 123524 626
rect 123832 610 124168 626
rect 124936 610 125272 626
rect 126132 610 126468 626
rect 127236 610 127572 626
rect 128340 610 128676 626
rect 123832 604 124180 610
rect 123832 598 124128 604
rect 122300 480 122328 546
rect 123312 490 123340 598
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 122728 462 123340 490
rect 123496 480 123524 598
rect 124128 546 124180 552
rect 124680 604 124732 610
rect 124936 604 125284 610
rect 124936 598 125232 604
rect 124680 546 124732 552
rect 125232 546 125284 552
rect 125876 604 125928 610
rect 126132 604 126480 610
rect 126132 598 126428 604
rect 125876 546 125928 552
rect 126428 546 126480 552
rect 126980 604 127032 610
rect 127236 604 127584 610
rect 127236 598 127532 604
rect 126980 546 127032 552
rect 127532 546 127584 552
rect 128176 604 128228 610
rect 128340 604 128688 610
rect 128340 598 128636 604
rect 128176 546 128228 552
rect 128636 546 128688 552
rect 129372 604 129424 610
rect 130640 598 130976 626
rect 131744 598 132080 626
rect 132940 620 133236 626
rect 134156 672 134208 678
rect 132940 614 133288 620
rect 132940 598 133276 614
rect 133892 610 134044 626
rect 134156 614 134208 620
rect 136180 672 136232 678
rect 137652 672 137704 678
rect 136232 620 136344 626
rect 136180 614 136344 620
rect 133880 604 134044 610
rect 129372 546 129424 552
rect 124692 480 124720 546
rect 125888 480 125916 546
rect 126992 480 127020 546
rect 128188 480 128216 546
rect 129384 480 129412 546
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 129832 128 129884 134
rect 129536 76 129832 82
rect 129536 70 129884 76
rect 130292 128 130344 134
rect 130538 82 130650 480
rect 130948 406 130976 598
rect 130936 400 130988 406
rect 130936 342 130988 348
rect 131734 354 131846 480
rect 132052 406 132080 598
rect 133932 598 134044 604
rect 133880 546 133932 552
rect 134168 480 134196 614
rect 135260 604 135312 610
rect 136192 598 136344 614
rect 137448 610 137600 626
rect 138756 672 138808 678
rect 137652 614 137704 620
rect 138552 620 138756 626
rect 140044 672 140096 678
rect 138552 614 138808 620
rect 136456 604 136508 610
rect 135260 546 135312 552
rect 137448 604 137612 610
rect 137448 598 137560 604
rect 136456 546 136508 552
rect 137560 546 137612 552
rect 134984 536 135036 542
rect 135036 484 135148 490
rect 131948 400 132000 406
rect 131734 348 131948 354
rect 131734 342 132000 348
rect 132040 400 132092 406
rect 132040 342 132092 348
rect 132930 354 133042 480
rect 133144 400 133196 406
rect 132930 348 133144 354
rect 132930 342 133196 348
rect 130344 76 130650 82
rect 130292 70 130650 76
rect 129536 54 129872 70
rect 130304 54 130650 70
rect 130538 -960 130650 54
rect 131734 326 131988 342
rect 132930 326 133184 342
rect 131734 -960 131846 326
rect 132930 -960 133042 326
rect 134126 -960 134238 480
rect 134984 478 135148 484
rect 135272 480 135300 546
rect 136468 480 136496 546
rect 137664 480 137692 614
rect 138552 598 138796 614
rect 139748 610 139992 626
rect 151360 672 151412 678
rect 142066 640 142122 649
rect 140044 614 140096 620
rect 138848 604 138900 610
rect 139748 604 140004 610
rect 139748 598 139952 604
rect 138848 546 138900 552
rect 139952 546 140004 552
rect 138860 480 138888 546
rect 140056 480 140084 614
rect 141240 604 141292 610
rect 141956 598 142066 626
rect 143446 640 143502 649
rect 142066 575 142122 584
rect 142264 598 142476 626
rect 143152 598 143446 626
rect 141240 546 141292 552
rect 141056 536 141108 542
rect 140852 484 141056 490
rect 134996 462 135148 478
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 140852 478 141108 484
rect 141252 480 141280 546
rect 142068 536 142120 542
rect 142264 490 142292 598
rect 142120 484 142292 490
rect 140852 462 141096 478
rect 141210 -960 141322 480
rect 142068 478 142292 484
rect 142448 480 142476 598
rect 144734 640 144790 649
rect 143446 575 143502 584
rect 143552 598 143764 626
rect 144256 610 144592 626
rect 144256 604 144604 610
rect 144256 598 144552 604
rect 143552 480 143580 598
rect 143736 513 143764 598
rect 145746 640 145802 649
rect 145452 598 145746 626
rect 144734 575 144790 584
rect 147126 640 147182 649
rect 146556 610 146892 626
rect 145746 575 145802 584
rect 145932 604 145984 610
rect 144552 546 144604 552
rect 143722 504 143778 513
rect 142080 462 142292 478
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144748 480 144776 575
rect 146556 604 146904 610
rect 146556 598 146852 604
rect 145932 546 145984 552
rect 148966 640 149022 649
rect 147126 575 147182 584
rect 148324 604 148376 610
rect 146852 546 146904 552
rect 145944 480 145972 546
rect 147140 480 147168 575
rect 148856 598 148966 626
rect 150622 640 150678 649
rect 148966 575 149022 584
rect 149348 598 149560 626
rect 148324 546 148376 552
rect 147770 504 147826 513
rect 143722 439 143778 448
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 147660 462 147770 490
rect 148336 480 148364 546
rect 149348 513 149376 598
rect 149334 504 149390 513
rect 147770 439 147826 448
rect 148294 -960 148406 480
rect 149532 480 149560 598
rect 151064 620 151360 626
rect 153016 672 153068 678
rect 151064 614 151412 620
rect 151818 640 151874 649
rect 151064 598 151400 614
rect 150622 575 150678 584
rect 152260 610 152596 626
rect 153660 672 153712 678
rect 153016 614 153068 620
rect 153364 620 153660 626
rect 155408 672 155460 678
rect 153364 614 153712 620
rect 152260 604 152608 610
rect 152260 598 152556 604
rect 151818 575 151874 584
rect 150254 504 150310 513
rect 149334 439 149390 448
rect 149490 -960 149602 480
rect 149960 462 150254 490
rect 150636 480 150664 575
rect 151832 480 151860 575
rect 152556 546 152608 552
rect 153028 480 153056 614
rect 153364 598 153700 614
rect 154468 610 154804 626
rect 162768 672 162820 678
rect 155408 614 155460 620
rect 154212 604 154264 610
rect 154468 604 154816 610
rect 154468 598 154764 604
rect 154212 546 154264 552
rect 154764 546 154816 552
rect 154224 480 154252 546
rect 155420 480 155448 614
rect 156768 610 157104 626
rect 156604 604 156656 610
rect 156768 604 157116 610
rect 156768 598 157064 604
rect 156604 546 156656 552
rect 157872 598 158208 626
rect 157064 546 157116 552
rect 156616 480 156644 546
rect 158180 542 158208 598
rect 158904 604 158956 610
rect 160172 598 160508 626
rect 161276 610 161612 626
rect 162472 620 162768 626
rect 164884 672 164936 678
rect 164790 640 164846 649
rect 162472 614 162820 620
rect 161276 604 161624 610
rect 161276 598 161572 604
rect 158904 546 158956 552
rect 158168 536 158220 542
rect 150254 439 150310 448
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 155960 128 156012 134
rect 155664 76 155960 82
rect 155664 70 156012 76
rect 155664 54 156000 70
rect 156574 -960 156686 480
rect 157524 128 157576 134
rect 157770 82 157882 480
rect 158168 478 158220 484
rect 158916 480 158944 546
rect 159732 536 159784 542
rect 157576 76 157882 82
rect 157524 70 157882 76
rect 157536 54 157882 70
rect 157770 -960 157882 54
rect 158874 -960 158986 480
rect 159732 478 159784 484
rect 159744 354 159772 478
rect 160070 354 160182 480
rect 160480 406 160508 598
rect 162472 598 162808 614
rect 163688 604 163740 610
rect 161572 546 161624 552
rect 164680 598 164790 626
rect 166080 672 166132 678
rect 164884 614 164936 620
rect 164790 575 164846 584
rect 163688 546 163740 552
rect 159744 326 160182 354
rect 160468 400 160520 406
rect 160468 342 160520 348
rect 159364 128 159416 134
rect 159068 76 159364 82
rect 159068 70 159416 76
rect 159068 54 159404 70
rect 160070 -960 160182 326
rect 161266 82 161378 480
rect 162462 354 162574 480
rect 163424 474 163576 490
rect 163700 480 163728 546
rect 164896 480 164924 614
rect 165876 610 166028 626
rect 167092 672 167144 678
rect 166080 614 166132 620
rect 166980 620 167092 626
rect 169576 672 169628 678
rect 167366 640 167422 649
rect 166980 614 167144 620
rect 165876 604 166040 610
rect 165876 598 165988 604
rect 165988 546 166040 552
rect 166092 480 166120 614
rect 166980 598 167132 614
rect 167196 598 167366 626
rect 167196 480 167224 598
rect 169482 640 169538 649
rect 167366 575 167422 584
rect 168380 604 168432 610
rect 169280 598 169482 626
rect 180892 672 180944 678
rect 171966 640 172022 649
rect 169576 614 169628 620
rect 169482 575 169538 584
rect 168380 546 168432 552
rect 168392 480 168420 546
rect 169588 480 169616 614
rect 170384 610 170720 626
rect 170384 604 170732 610
rect 170384 598 170680 604
rect 170680 546 170732 552
rect 170784 598 170996 626
rect 170784 480 170812 598
rect 163412 468 163576 474
rect 163464 462 163576 468
rect 163412 410 163464 416
rect 162676 400 162728 406
rect 162462 348 162676 354
rect 162462 342 162728 348
rect 162462 326 162716 342
rect 161480 128 161532 134
rect 161266 76 161480 82
rect 161266 70 161532 76
rect 161266 54 161520 70
rect 161266 -960 161378 54
rect 162462 -960 162574 326
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168194 368 168250 377
rect 168084 326 168194 354
rect 168194 303 168250 312
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 170968 377 170996 598
rect 172978 640 173034 649
rect 172684 598 172978 626
rect 171966 575 172022 584
rect 175462 640 175518 649
rect 172978 575 173034 584
rect 173164 604 173216 610
rect 171980 480 172008 575
rect 173164 546 173216 552
rect 174096 598 174308 626
rect 173176 480 173204 546
rect 173898 504 173954 513
rect 170954 368 171010 377
rect 171690 368 171746 377
rect 171488 326 171690 354
rect 170954 303 171010 312
rect 171690 303 171746 312
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 173788 462 173898 490
rect 174096 490 174124 598
rect 173898 439 173954 448
rect 174004 462 174124 490
rect 174280 480 174308 598
rect 176382 640 176438 649
rect 176088 598 176382 626
rect 175462 575 175518 584
rect 179050 640 179106 649
rect 176382 575 176438 584
rect 176672 598 176884 626
rect 175476 480 175504 575
rect 176672 480 176700 598
rect 176856 513 176884 598
rect 177684 598 177896 626
rect 176842 504 176898 513
rect 174004 377 174032 462
rect 173990 368 174046 377
rect 173990 303 174046 312
rect 174238 -960 174350 480
rect 175186 368 175242 377
rect 174984 326 175186 354
rect 175186 303 175242 312
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177486 504 177542 513
rect 177192 462 177486 490
rect 176842 439 176898 448
rect 177486 439 177542 448
rect 177684 377 177712 598
rect 177868 480 177896 598
rect 180246 640 180302 649
rect 179492 610 179828 626
rect 179492 604 179840 610
rect 179492 598 179788 604
rect 179050 575 179106 584
rect 179064 480 179092 575
rect 180596 620 180892 626
rect 183744 672 183796 678
rect 182086 640 182142 649
rect 180596 614 180944 620
rect 180596 598 180932 614
rect 181272 598 181484 626
rect 181792 598 182086 626
rect 180246 575 180302 584
rect 179788 546 179840 552
rect 180260 480 180288 575
rect 177670 368 177726 377
rect 177670 303 177726 312
rect 177826 -960 177938 480
rect 178682 368 178738 377
rect 178388 326 178682 354
rect 178682 303 178738 312
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181272 377 181300 598
rect 181456 480 181484 598
rect 182896 610 183232 626
rect 186136 672 186188 678
rect 183744 614 183796 620
rect 184938 640 184994 649
rect 182086 575 182142 584
rect 182548 604 182600 610
rect 182896 604 183244 610
rect 182896 598 183192 604
rect 182548 546 182600 552
rect 183192 546 183244 552
rect 182560 480 182588 546
rect 183756 480 183784 614
rect 191104 672 191156 678
rect 186136 614 186188 620
rect 184938 575 184994 584
rect 184952 480 184980 575
rect 186148 480 186176 614
rect 187404 598 187740 626
rect 188600 598 188844 626
rect 189704 610 190040 626
rect 190808 620 191104 626
rect 194416 672 194468 678
rect 192298 640 192354 649
rect 190808 614 191156 620
rect 189704 604 190052 610
rect 189704 598 190000 604
rect 187712 542 187740 598
rect 187700 536 187752 542
rect 186594 504 186650 513
rect 181258 368 181314 377
rect 181258 303 181314 312
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184296 128 184348 134
rect 184000 76 184296 82
rect 184000 70 184348 76
rect 184000 54 184336 70
rect 184910 -960 185022 480
rect 185492 128 185544 134
rect 185196 76 185492 82
rect 185196 70 185544 76
rect 185196 54 185532 70
rect 186106 -960 186218 480
rect 186300 462 186594 490
rect 186594 439 186650 448
rect 187302 218 187414 480
rect 187700 478 187752 484
rect 186976 202 187414 218
rect 186964 196 187414 202
rect 187016 190 187414 196
rect 186964 138 187016 144
rect 187302 -960 187414 190
rect 188252 128 188304 134
rect 188498 82 188610 480
rect 188816 406 188844 598
rect 190808 598 191144 614
rect 192004 598 192298 626
rect 211620 672 211672 678
rect 194416 614 194468 620
rect 195610 640 195666 649
rect 192298 575 192354 584
rect 193220 604 193272 610
rect 190000 546 190052 552
rect 193220 546 193272 552
rect 191012 536 191064 542
rect 189906 504 189962 513
rect 188804 400 188856 406
rect 188804 342 188856 348
rect 188304 76 188610 82
rect 188252 70 188610 76
rect 188264 54 188610 70
rect 188498 -960 188610 54
rect 189694 218 189806 480
rect 189906 439 189962 448
rect 189920 218 189948 439
rect 189694 190 189948 218
rect 190798 354 190910 480
rect 191012 478 191064 484
rect 192944 536 192996 542
rect 192996 484 193108 490
rect 191024 354 191052 478
rect 190798 326 191052 354
rect 191994 354 192106 480
rect 192944 478 193108 484
rect 193232 480 193260 546
rect 194046 504 194102 513
rect 192956 462 193108 478
rect 192208 400 192260 406
rect 191994 348 192208 354
rect 191994 342 192260 348
rect 191994 326 192248 342
rect 189694 -960 189806 190
rect 190798 -960 190910 326
rect 191994 -960 192106 326
rect 193190 -960 193302 480
rect 194102 462 194212 490
rect 194428 480 194456 614
rect 197910 640 197966 649
rect 195610 575 195666 584
rect 196808 604 196860 610
rect 195624 480 195652 575
rect 200026 640 200082 649
rect 197910 575 197966 584
rect 199108 604 199160 610
rect 196808 546 196860 552
rect 196820 480 196848 546
rect 197924 480 197952 575
rect 199916 598 200026 626
rect 203890 640 203946 649
rect 203320 610 203656 626
rect 203320 604 203668 610
rect 203320 598 203616 604
rect 200026 575 200082 584
rect 199108 546 199160 552
rect 200132 564 200344 592
rect 198922 504 198978 513
rect 194046 439 194102 448
rect 194386 -960 194498 480
rect 195244 400 195296 406
rect 195296 348 195408 354
rect 195244 342 195408 348
rect 195256 326 195408 342
rect 195582 -960 195694 480
rect 196622 368 196678 377
rect 196512 326 196622 354
rect 196622 303 196678 312
rect 196778 -960 196890 480
rect 197726 96 197782 105
rect 197616 54 197726 82
rect 197726 31 197782 40
rect 197882 -960 197994 480
rect 198812 462 198922 490
rect 199120 480 199148 546
rect 198922 439 198978 448
rect 199078 -960 199190 480
rect 200132 377 200160 564
rect 200316 480 200344 564
rect 201512 564 201724 592
rect 201314 504 201370 513
rect 200118 368 200174 377
rect 200118 303 200174 312
rect 200274 -960 200386 480
rect 201112 462 201314 490
rect 201512 480 201540 564
rect 201314 439 201370 448
rect 201470 -960 201582 480
rect 201696 105 201724 564
rect 202524 564 202736 592
rect 202524 377 202552 564
rect 202708 480 202736 564
rect 203890 575 203946 584
rect 204166 640 204222 649
rect 207386 640 207442 649
rect 205620 610 205772 626
rect 205620 604 205784 610
rect 205620 598 205732 604
rect 204166 575 204168 584
rect 203616 546 203668 552
rect 203904 480 203932 575
rect 204220 575 204222 584
rect 204168 546 204220 552
rect 204916 564 205128 592
rect 204916 513 204944 564
rect 204902 504 204958 513
rect 202510 368 202566 377
rect 202510 303 202566 312
rect 202418 232 202474 241
rect 202216 190 202418 218
rect 202418 167 202474 176
rect 201682 96 201738 105
rect 201682 31 201738 40
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205100 480 205128 564
rect 205732 546 205784 552
rect 206020 564 206232 592
rect 208214 640 208270 649
rect 207920 598 208214 626
rect 207386 575 207442 584
rect 208214 575 208270 584
rect 208398 640 208454 649
rect 209318 640 209374 649
rect 208398 575 208454 584
rect 208596 598 208808 626
rect 209024 598 209318 626
rect 204902 439 204958 448
rect 204810 368 204866 377
rect 204516 326 204810 354
rect 204810 303 204866 312
rect 205058 -960 205170 480
rect 206020 241 206048 564
rect 206204 480 206232 564
rect 206926 504 206982 513
rect 206006 232 206062 241
rect 206006 167 206062 176
rect 206162 -960 206274 480
rect 206724 462 206926 490
rect 207400 480 207428 575
rect 208412 542 208440 575
rect 208400 536 208452 542
rect 206926 439 206982 448
rect 207358 -960 207470 480
rect 208400 478 208452 484
rect 208596 480 208624 598
rect 208554 -960 208666 480
rect 208780 377 208808 598
rect 210128 610 210464 626
rect 209318 575 209374 584
rect 209780 604 209832 610
rect 210128 604 210476 610
rect 210128 598 210424 604
rect 209780 546 209832 552
rect 210424 546 210476 552
rect 210804 598 211016 626
rect 211324 620 211620 626
rect 215668 672 215720 678
rect 211324 614 211672 620
rect 213366 640 213422 649
rect 211324 598 211660 614
rect 212172 604 212224 610
rect 209792 480 209820 546
rect 210804 513 210832 598
rect 210790 504 210846 513
rect 208766 368 208822 377
rect 208766 303 208822 312
rect 209750 -960 209862 480
rect 210988 480 211016 598
rect 220176 672 220228 678
rect 216126 640 216182 649
rect 215668 614 215720 620
rect 213366 575 213422 584
rect 214472 604 214524 610
rect 212172 546 212224 552
rect 212184 480 212212 546
rect 210790 439 210846 448
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 212428 474 212580 490
rect 213380 480 213408 575
rect 214472 546 214524 552
rect 214484 480 214512 546
rect 215680 480 215708 614
rect 215832 598 216126 626
rect 216936 598 217272 626
rect 218132 598 218468 626
rect 219236 610 219572 626
rect 225328 672 225380 678
rect 220726 640 220782 649
rect 220228 620 220340 626
rect 220176 614 220340 620
rect 219236 604 219584 610
rect 219236 598 219532 604
rect 216126 575 216182 584
rect 212428 468 212592 474
rect 212428 462 212540 468
rect 212540 410 212592 416
rect 213338 -960 213450 480
rect 213532 66 213868 82
rect 213532 60 213880 66
rect 213532 54 213828 60
rect 213828 2 213880 8
rect 214442 -960 214554 480
rect 215024 128 215076 134
rect 214728 76 215024 82
rect 214728 70 215076 76
rect 214728 54 215064 70
rect 215638 -960 215750 480
rect 216588 468 216640 474
rect 216588 410 216640 416
rect 216600 354 216628 410
rect 216834 354 216946 480
rect 217244 406 217272 598
rect 218440 542 218468 598
rect 220188 598 220340 614
rect 220464 598 220726 626
rect 219532 546 219584 552
rect 218428 536 218480 542
rect 216600 326 216946 354
rect 217232 400 217284 406
rect 217232 342 217284 348
rect 216834 -960 216946 326
rect 218030 82 218142 480
rect 218428 478 218480 484
rect 220464 480 220492 598
rect 221830 640 221886 649
rect 221536 598 221830 626
rect 220726 575 220782 584
rect 221830 575 221886 584
rect 222764 598 222976 626
rect 224940 610 225092 626
rect 225156 620 225328 626
rect 226156 672 226208 678
rect 225156 614 225380 620
rect 226044 620 226156 626
rect 231032 672 231084 678
rect 226044 614 226208 620
rect 226338 640 226394 649
rect 217704 66 218142 82
rect 217692 60 218142 66
rect 217744 54 218142 60
rect 217692 2 217744 8
rect 218030 -960 218142 54
rect 219226 82 219338 480
rect 219440 128 219492 134
rect 219226 76 219440 82
rect 219226 70 219492 76
rect 219226 54 219480 70
rect 219226 -960 219338 54
rect 220422 -960 220534 480
rect 221526 354 221638 480
rect 222488 474 222640 490
rect 222764 480 222792 598
rect 222948 542 222976 598
rect 223948 604 224000 610
rect 224940 604 225104 610
rect 224940 598 225052 604
rect 223948 546 224000 552
rect 225052 546 225104 552
rect 225156 598 225368 614
rect 226044 598 226196 614
rect 222936 536 222988 542
rect 222476 468 222640 474
rect 222528 462 222640 468
rect 222476 410 222528 416
rect 221740 400 221792 406
rect 221526 348 221740 354
rect 221526 342 221792 348
rect 221526 326 221780 342
rect 221526 -960 221638 326
rect 222722 -960 222834 480
rect 222936 478 222988 484
rect 223578 504 223634 513
rect 223634 462 223744 490
rect 223960 480 223988 546
rect 225156 480 225184 598
rect 228730 640 228786 649
rect 226338 575 226394 584
rect 227364 598 227576 626
rect 226352 480 226380 575
rect 227364 542 227392 598
rect 227352 536 227404 542
rect 223578 439 223634 448
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227352 478 227404 484
rect 227548 480 227576 598
rect 230938 640 230994 649
rect 228730 575 228786 584
rect 229836 604 229888 610
rect 228744 480 228772 575
rect 230644 598 230938 626
rect 234620 672 234672 678
rect 231032 614 231084 620
rect 230938 575 230994 584
rect 229836 546 229888 552
rect 229652 536 229704 542
rect 229448 484 229652 490
rect 227148 66 227392 82
rect 227148 60 227404 66
rect 227148 54 227352 60
rect 227352 2 227404 8
rect 227506 -960 227618 480
rect 228548 128 228600 134
rect 228344 76 228548 82
rect 228344 70 228600 76
rect 228344 54 228588 70
rect 228702 -960 228814 480
rect 229448 478 229704 484
rect 229848 480 229876 546
rect 231044 480 231072 614
rect 231748 610 231900 626
rect 231748 604 231912 610
rect 231748 598 231860 604
rect 231860 546 231912 552
rect 232056 598 232268 626
rect 229448 462 229692 478
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232056 66 232084 598
rect 232240 480 232268 598
rect 233252 598 233464 626
rect 235448 672 235500 678
rect 234620 614 234672 620
rect 235152 620 235448 626
rect 240508 672 240560 678
rect 235152 614 235500 620
rect 235814 640 235870 649
rect 233148 536 233200 542
rect 232852 484 233148 490
rect 232044 60 232096 66
rect 232044 2 232096 8
rect 232198 -960 232310 480
rect 232852 478 233200 484
rect 232852 462 233188 478
rect 233252 134 233280 598
rect 233436 480 233464 598
rect 233240 128 233292 134
rect 233240 70 233292 76
rect 233394 -960 233506 480
rect 234048 474 234384 490
rect 234632 480 234660 614
rect 235152 598 235488 614
rect 237746 640 237802 649
rect 235814 575 235870 584
rect 237012 604 237064 610
rect 235828 480 235856 575
rect 237452 598 237746 626
rect 238556 610 238892 626
rect 241152 672 241204 678
rect 240508 614 240560 620
rect 240856 620 241152 626
rect 245752 672 245804 678
rect 240856 614 241204 620
rect 242898 640 242954 649
rect 237746 575 237802 584
rect 238116 604 238168 610
rect 237012 546 237064 552
rect 238556 604 238904 610
rect 238556 598 238852 604
rect 238116 546 238168 552
rect 238852 546 238904 552
rect 239048 564 239352 592
rect 237024 480 237052 546
rect 238128 480 238156 546
rect 234048 468 234396 474
rect 234048 462 234344 468
rect 234344 410 234396 416
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236256 66 236592 82
rect 236256 60 236604 66
rect 236256 54 236552 60
rect 236552 2 236604 8
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239048 474 239076 564
rect 239324 480 239352 564
rect 239956 536 240008 542
rect 239660 484 239956 490
rect 239036 468 239088 474
rect 239036 410 239088 416
rect 239282 -960 239394 480
rect 239660 478 240008 484
rect 240520 480 240548 614
rect 240856 598 241192 614
rect 241532 564 241744 592
rect 245364 620 245752 626
rect 247960 672 248012 678
rect 245364 614 245804 620
rect 242898 575 242954 584
rect 244096 604 244148 610
rect 239660 462 239996 478
rect 240478 -960 240590 480
rect 241532 218 241560 564
rect 241716 480 241744 564
rect 242254 504 242310 513
rect 241440 190 241560 218
rect 241440 66 241468 190
rect 241428 60 241480 66
rect 241428 2 241480 8
rect 241674 -960 241786 480
rect 241960 462 242254 490
rect 242912 480 242940 575
rect 244096 546 244148 552
rect 245200 604 245252 610
rect 245364 598 245792 614
rect 246028 604 246080 610
rect 245200 546 245252 552
rect 246468 598 246804 626
rect 247664 620 247960 626
rect 253480 672 253532 678
rect 249706 640 249762 649
rect 247664 614 248012 620
rect 247664 598 248000 614
rect 248768 598 249104 626
rect 246028 546 246080 552
rect 244108 480 244136 546
rect 244556 536 244608 542
rect 244260 484 244556 490
rect 242254 439 242310 448
rect 242870 -960 242982 480
rect 243360 400 243412 406
rect 243064 348 243360 354
rect 243064 342 243412 348
rect 243064 326 243400 342
rect 244066 -960 244178 480
rect 244260 478 244608 484
rect 245212 480 245240 546
rect 244260 462 244596 478
rect 245170 -960 245282 480
rect 246040 354 246068 546
rect 246366 354 246478 480
rect 246040 326 246478 354
rect 246776 338 246804 598
rect 249076 542 249104 598
rect 249762 598 249872 626
rect 254584 672 254636 678
rect 253480 614 253532 620
rect 254472 620 254584 626
rect 257252 672 257304 678
rect 254472 614 254636 620
rect 255870 640 255926 649
rect 249984 604 250036 610
rect 249706 575 249762 584
rect 249984 546 250036 552
rect 251180 604 251232 610
rect 251180 546 251232 552
rect 252376 604 252428 610
rect 252376 546 252428 552
rect 249064 536 249116 542
rect 247314 504 247370 513
rect 247314 439 247370 448
rect 246366 -960 246478 326
rect 246764 332 246816 338
rect 246764 274 246816 280
rect 247328 218 247356 439
rect 247562 218 247674 480
rect 247328 190 247674 218
rect 247562 -960 247674 190
rect 248758 354 248870 480
rect 249064 478 249116 484
rect 249996 480 250024 546
rect 251192 480 251220 546
rect 252388 480 252416 546
rect 248972 400 249024 406
rect 248758 348 248972 354
rect 248758 342 249024 348
rect 248758 326 249012 342
rect 248758 -960 248870 326
rect 249954 -960 250066 480
rect 250904 400 250956 406
rect 250956 348 251068 354
rect 250904 342 251068 348
rect 250916 326 251068 342
rect 251150 -960 251262 480
rect 252020 202 252172 218
rect 252008 196 252172 202
rect 252060 190 252172 196
rect 252008 138 252060 144
rect 252346 -960 252458 480
rect 253124 474 253276 490
rect 253492 480 253520 614
rect 254472 598 254624 614
rect 254676 604 254728 610
rect 257252 614 257304 620
rect 258264 672 258316 678
rect 260472 672 260524 678
rect 258264 614 258316 620
rect 260176 620 260472 626
rect 266544 672 266596 678
rect 260176 614 260524 620
rect 255870 575 255926 584
rect 257068 604 257120 610
rect 254676 546 254728 552
rect 254688 480 254716 546
rect 255884 480 255912 575
rect 257068 546 257120 552
rect 257080 480 257108 546
rect 253112 468 253276 474
rect 253164 462 253276 468
rect 253112 410 253164 416
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255688 264 255740 270
rect 255576 212 255688 218
rect 255576 206 255740 212
rect 255576 190 255728 206
rect 255842 -960 255954 480
rect 256772 338 256924 354
rect 256772 332 256936 338
rect 256772 326 256884 332
rect 256884 274 256936 280
rect 257038 -960 257150 480
rect 257264 202 257292 614
rect 258276 480 258304 614
rect 260176 598 260512 614
rect 262384 610 262720 626
rect 268844 672 268896 678
rect 267278 640 267334 649
rect 266544 614 266596 620
rect 260656 604 260708 610
rect 259288 564 259500 592
rect 259288 490 259316 564
rect 257876 202 258028 218
rect 257252 196 257304 202
rect 257876 196 258040 202
rect 257876 190 257988 196
rect 257252 138 257304 144
rect 257988 138 258040 144
rect 258234 -960 258346 480
rect 259104 474 259316 490
rect 259472 480 259500 564
rect 262384 604 262732 610
rect 262384 598 262680 604
rect 260656 546 260708 552
rect 261772 564 261984 592
rect 260668 480 260696 546
rect 261576 536 261628 542
rect 261280 484 261576 490
rect 259092 468 259316 474
rect 259144 462 259316 468
rect 259092 410 259144 416
rect 259276 400 259328 406
rect 258980 348 259276 354
rect 258980 342 259328 348
rect 258980 326 259316 342
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261280 478 261628 484
rect 261772 480 261800 564
rect 261280 462 261616 478
rect 261730 -960 261842 480
rect 261956 270 261984 564
rect 262680 546 262732 552
rect 262784 564 262996 592
rect 262784 338 262812 564
rect 262968 480 262996 564
rect 263980 564 264192 592
rect 262772 332 262824 338
rect 262772 274 262824 280
rect 261944 264 261996 270
rect 261944 206 261996 212
rect 262926 -960 263038 480
rect 263580 474 263732 490
rect 263580 468 263744 474
rect 263580 462 263692 468
rect 263692 410 263744 416
rect 263980 354 264008 564
rect 264164 480 264192 564
rect 265176 564 265388 592
rect 265176 490 265204 564
rect 263888 326 264008 354
rect 263888 202 263916 326
rect 263876 196 263928 202
rect 263876 138 263928 144
rect 264122 -960 264234 480
rect 264992 462 265204 490
rect 265360 480 265388 564
rect 266556 480 266584 614
rect 266984 598 267278 626
rect 272892 672 272944 678
rect 268844 614 268896 620
rect 267278 575 267334 584
rect 267740 604 267792 610
rect 267740 546 267792 552
rect 267752 480 267780 546
rect 268384 536 268436 542
rect 268088 484 268384 490
rect 264992 406 265020 462
rect 264980 400 265032 406
rect 264980 342 265032 348
rect 264888 264 264940 270
rect 264684 212 264888 218
rect 264684 206 264940 212
rect 264684 190 264928 206
rect 265318 -960 265430 480
rect 266084 128 266136 134
rect 265788 76 266084 82
rect 265788 70 266136 76
rect 265788 54 266124 70
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268088 478 268436 484
rect 268856 480 268884 614
rect 270388 610 270724 626
rect 270040 604 270092 610
rect 270388 604 270736 610
rect 270388 598 270684 604
rect 270040 546 270092 552
rect 270684 546 270736 552
rect 271064 598 271276 626
rect 268088 462 268424 478
rect 268814 -960 268926 480
rect 269192 474 269528 490
rect 270052 480 270080 546
rect 269192 468 269540 474
rect 269192 462 269488 468
rect 269488 410 269540 416
rect 270010 -960 270122 480
rect 271064 270 271092 598
rect 271248 480 271276 598
rect 272260 598 272472 626
rect 272596 620 272892 626
rect 277492 672 277544 678
rect 272596 614 272944 620
rect 273626 640 273682 649
rect 272596 598 272932 614
rect 271052 264 271104 270
rect 271052 206 271104 212
rect 271206 -960 271318 480
rect 271788 400 271840 406
rect 271492 348 271788 354
rect 272260 354 272288 598
rect 272444 480 272472 598
rect 275190 640 275246 649
rect 274896 598 275190 626
rect 273626 575 273682 584
rect 275190 575 275246 584
rect 275848 598 276000 626
rect 277196 620 277492 626
rect 284300 672 284352 678
rect 282090 640 282146 649
rect 277196 614 277544 620
rect 276756 604 276808 610
rect 273640 480 273668 575
rect 274548 536 274600 542
rect 271492 342 271840 348
rect 271492 326 271828 342
rect 272168 326 272288 354
rect 272168 134 272196 326
rect 272156 128 272208 134
rect 272156 70 272208 76
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274548 478 274600 484
rect 274560 354 274588 478
rect 274794 354 274906 480
rect 274560 326 274906 354
rect 275848 338 275876 598
rect 277196 598 277532 614
rect 278300 598 278636 626
rect 281704 610 281856 626
rect 276756 546 276808 552
rect 275990 354 276102 480
rect 276204 468 276256 474
rect 276204 410 276256 416
rect 276216 354 276244 410
rect 274088 264 274140 270
rect 273792 212 274088 218
rect 273792 206 274140 212
rect 273792 190 274128 206
rect 274794 -960 274906 326
rect 275836 332 275888 338
rect 275836 274 275888 280
rect 275990 326 276244 354
rect 276768 354 276796 546
rect 278608 542 278636 598
rect 279516 604 279568 610
rect 279516 546 279568 552
rect 280712 604 280764 610
rect 281704 604 281868 610
rect 281704 598 281816 604
rect 280712 546 280764 552
rect 281816 546 281868 552
rect 281920 598 282090 626
rect 278596 536 278648 542
rect 277094 354 277206 480
rect 276768 326 277206 354
rect 275990 -960 276102 326
rect 277094 -960 277206 326
rect 278290 354 278402 480
rect 278596 478 278648 484
rect 279252 474 279404 490
rect 279528 480 279556 546
rect 280724 480 280752 546
rect 281920 480 281948 598
rect 286600 672 286652 678
rect 284300 614 284352 620
rect 285678 640 285734 649
rect 282090 575 282146 584
rect 283116 564 283328 592
rect 283116 480 283144 564
rect 279240 468 279404 474
rect 279292 462 279404 468
rect 279240 410 279292 416
rect 278504 400 278556 406
rect 278290 348 278504 354
rect 278290 342 278556 348
rect 278290 326 278544 342
rect 278290 -960 278402 326
rect 279486 -960 279598 480
rect 280436 400 280488 406
rect 280488 348 280600 354
rect 280436 342 280600 348
rect 280448 326 280600 342
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 282808 202 282960 218
rect 282808 196 282972 202
rect 282808 190 282920 196
rect 282920 138 282972 144
rect 283074 -960 283186 480
rect 283300 338 283328 564
rect 284312 480 284340 614
rect 285404 604 285456 610
rect 288992 672 289044 678
rect 287794 640 287850 649
rect 286600 614 286652 620
rect 285678 575 285734 584
rect 285404 546 285456 552
rect 285218 504 285274 513
rect 284004 338 284156 354
rect 283288 332 283340 338
rect 284004 332 284168 338
rect 284004 326 284116 332
rect 283288 274 283340 280
rect 284116 274 284168 280
rect 284270 -960 284382 480
rect 285108 462 285218 490
rect 285416 480 285444 546
rect 285218 439 285274 448
rect 285374 -960 285486 480
rect 285692 406 285720 575
rect 286612 480 286640 614
rect 287408 610 287652 626
rect 287408 604 287664 610
rect 287408 598 287612 604
rect 291108 672 291160 678
rect 288992 614 289044 620
rect 287794 575 287850 584
rect 287612 546 287664 552
rect 287808 480 287836 575
rect 285680 400 285732 406
rect 286414 368 286470 377
rect 285680 342 285732 348
rect 286304 326 286414 354
rect 286414 303 286470 312
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288512 474 288848 490
rect 289004 480 289032 614
rect 290016 598 290228 626
rect 290812 620 291108 626
rect 293408 672 293460 678
rect 292578 640 292634 649
rect 290812 614 291160 620
rect 290812 598 291148 614
rect 291212 598 291424 626
rect 288512 468 288860 474
rect 288512 462 288808 468
rect 288808 410 288860 416
rect 288962 -960 289074 480
rect 289820 264 289872 270
rect 289708 212 289820 218
rect 289708 206 289872 212
rect 289708 190 289860 206
rect 290016 202 290044 598
rect 290200 480 290228 598
rect 290004 196 290056 202
rect 290004 138 290056 144
rect 290158 -960 290270 480
rect 291212 338 291240 598
rect 291396 480 291424 598
rect 293112 620 293408 626
rect 298468 672 298520 678
rect 294602 640 294658 649
rect 293112 614 293460 620
rect 293112 598 293448 614
rect 293512 598 293724 626
rect 292578 575 292634 584
rect 292592 480 292620 575
rect 291200 332 291252 338
rect 291200 274 291252 280
rect 291354 -960 291466 480
rect 291916 66 292252 82
rect 291916 60 292264 66
rect 291916 54 292212 60
rect 292212 2 292264 8
rect 292550 -960 292662 480
rect 293406 368 293462 377
rect 293512 354 293540 598
rect 293696 480 293724 598
rect 296074 640 296130 649
rect 295320 610 295656 626
rect 294602 575 294658 584
rect 294880 604 294932 610
rect 294512 536 294564 542
rect 294216 484 294512 490
rect 293462 326 293540 354
rect 293406 303 293462 312
rect 293654 -960 293766 480
rect 294216 478 294564 484
rect 294216 462 294552 478
rect 294616 474 294644 575
rect 295320 604 295668 610
rect 295320 598 295616 604
rect 294880 546 294932 552
rect 300216 672 300268 678
rect 298468 614 298520 620
rect 299920 620 300216 626
rect 307668 672 307720 678
rect 305826 640 305882 649
rect 299920 614 300268 620
rect 296074 575 296130 584
rect 295616 546 295668 552
rect 294892 480 294920 546
rect 296088 480 296116 575
rect 297008 564 297312 592
rect 294604 468 294656 474
rect 294604 410 294656 416
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 296516 338 296852 354
rect 296516 332 296864 338
rect 296516 326 296812 332
rect 296812 274 296864 280
rect 297008 270 297036 564
rect 297284 480 297312 564
rect 298480 480 298508 614
rect 299920 598 300256 614
rect 300596 598 300808 626
rect 299492 564 299704 592
rect 299492 490 299520 564
rect 296996 264 297048 270
rect 296996 206 297048 212
rect 297242 -960 297354 480
rect 297916 264 297968 270
rect 297620 212 297916 218
rect 297620 206 297968 212
rect 297620 190 297956 206
rect 298438 -960 298550 480
rect 299400 462 299520 490
rect 299676 480 299704 564
rect 300596 542 300624 598
rect 300584 536 300636 542
rect 299020 400 299072 406
rect 298724 348 299020 354
rect 298724 342 299072 348
rect 298724 326 299060 342
rect 299400 134 299428 462
rect 299388 128 299440 134
rect 299388 70 299440 76
rect 299634 -960 299746 480
rect 300584 478 300636 484
rect 300780 480 300808 598
rect 303160 604 303212 610
rect 301792 564 302004 592
rect 301320 536 301372 542
rect 301024 484 301320 490
rect 300738 -960 300850 480
rect 301024 478 301372 484
rect 301024 462 301360 478
rect 301792 474 301820 564
rect 301976 480 302004 564
rect 304428 598 304764 626
rect 305532 598 305826 626
rect 303160 546 303212 552
rect 303172 480 303200 546
rect 301780 468 301832 474
rect 301780 410 301832 416
rect 301934 -960 302046 480
rect 302128 202 302464 218
rect 302128 196 302476 202
rect 302128 190 302424 196
rect 302424 138 302476 144
rect 303130 -960 303242 480
rect 303324 474 303660 490
rect 303324 468 303672 474
rect 303324 462 303620 468
rect 303620 410 303672 416
rect 304326 354 304438 480
rect 304000 338 304438 354
rect 304736 338 304764 598
rect 306728 598 307064 626
rect 309968 672 310020 678
rect 307720 620 307832 626
rect 307668 614 307832 620
rect 315948 672 316000 678
rect 313830 640 313886 649
rect 310020 620 310132 626
rect 309968 614 310132 620
rect 307680 598 307832 614
rect 307944 604 307996 610
rect 305826 575 305882 584
rect 307036 513 307064 598
rect 307944 546 307996 552
rect 309048 604 309100 610
rect 309980 598 310132 614
rect 310244 604 310296 610
rect 309048 546 309100 552
rect 310244 546 310296 552
rect 311440 604 311492 610
rect 311440 546 311492 552
rect 312636 604 312688 610
rect 313830 575 313886 584
rect 315026 640 315082 649
rect 315836 620 315948 626
rect 318524 672 318576 678
rect 315836 614 316000 620
rect 316590 640 316646 649
rect 315836 598 315988 614
rect 316224 604 316276 610
rect 315026 575 315082 584
rect 312636 546 312688 552
rect 307022 504 307078 513
rect 303988 332 304438 338
rect 304040 326 304438 332
rect 303988 274 304040 280
rect 304326 -960 304438 326
rect 304724 332 304776 338
rect 304724 274 304776 280
rect 305522 218 305634 480
rect 306718 354 306830 480
rect 307956 480 307984 546
rect 309060 480 309088 546
rect 310256 480 310284 546
rect 311452 480 311480 546
rect 307022 439 307078 448
rect 306932 400 306984 406
rect 306718 348 306932 354
rect 306718 342 306984 348
rect 306718 326 306972 342
rect 305736 264 305788 270
rect 305522 212 305736 218
rect 305522 206 305788 212
rect 305522 190 305776 206
rect 305522 -960 305634 190
rect 306718 -960 306830 326
rect 307914 -960 308026 480
rect 308772 264 308824 270
rect 308824 212 308936 218
rect 308772 206 308936 212
rect 308784 190 308936 206
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311072 400 311124 406
rect 311124 348 311236 354
rect 311072 342 311236 348
rect 311084 326 311236 342
rect 311410 -960 311522 480
rect 312340 474 312492 490
rect 312648 480 312676 546
rect 313844 480 313872 575
rect 315040 480 315068 575
rect 317326 640 317382 649
rect 316940 610 317184 626
rect 316940 604 317196 610
rect 316940 598 317144 604
rect 316590 575 316646 584
rect 316224 546 316276 552
rect 316236 480 316264 546
rect 312340 468 312504 474
rect 312340 462 312452 468
rect 312452 410 312504 416
rect 312606 -960 312718 480
rect 313536 202 313688 218
rect 313536 196 313700 202
rect 313536 190 313648 196
rect 313648 138 313700 144
rect 313802 -960 313914 480
rect 314752 128 314804 134
rect 314640 76 314752 82
rect 314640 70 314804 76
rect 314640 54 314792 70
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 316604 270 316632 575
rect 324412 672 324464 678
rect 318524 614 318576 620
rect 317326 575 317382 584
rect 317144 546 317196 552
rect 317340 480 317368 575
rect 318536 480 318564 614
rect 319548 598 319760 626
rect 319352 536 319404 542
rect 319240 484 319352 490
rect 316592 264 316644 270
rect 316592 206 316644 212
rect 317298 -960 317410 480
rect 318044 338 318380 354
rect 318044 332 318392 338
rect 318044 326 318340 332
rect 318340 274 318392 280
rect 318494 -960 318606 480
rect 319240 478 319404 484
rect 319240 462 319392 478
rect 319548 406 319576 598
rect 319732 480 319760 598
rect 320744 598 320956 626
rect 325148 672 325200 678
rect 324412 614 324464 620
rect 324852 620 325148 626
rect 333612 672 333664 678
rect 328458 640 328514 649
rect 324852 614 325200 620
rect 319536 400 319588 406
rect 319536 342 319588 348
rect 319690 -960 319802 480
rect 320744 474 320772 598
rect 320928 480 320956 598
rect 321940 564 322152 592
rect 321940 490 321968 564
rect 320732 468 320784 474
rect 320732 410 320784 416
rect 320640 128 320692 134
rect 320344 76 320640 82
rect 320344 70 320692 76
rect 320344 54 320680 70
rect 320886 -960 320998 480
rect 321448 462 321600 490
rect 321572 406 321600 462
rect 321848 462 321968 490
rect 322124 480 322152 564
rect 323136 564 323348 592
rect 321560 400 321612 406
rect 321560 342 321612 348
rect 321848 202 321876 462
rect 321836 196 321888 202
rect 321836 138 321888 144
rect 322082 -960 322194 480
rect 322644 474 322888 490
rect 322644 468 322900 474
rect 322644 462 322848 468
rect 322848 410 322900 416
rect 323136 82 323164 564
rect 323320 480 323348 564
rect 324424 480 324452 614
rect 324852 598 325188 614
rect 325608 604 325660 610
rect 325608 546 325660 552
rect 326632 598 326844 626
rect 327152 610 327488 626
rect 327152 604 327500 610
rect 327152 598 327448 604
rect 325620 480 325648 546
rect 322860 66 323164 82
rect 322848 60 323164 66
rect 322900 54 323164 60
rect 322848 2 322900 8
rect 323278 -960 323390 480
rect 323748 66 324084 82
rect 323748 60 324096 66
rect 323748 54 324044 60
rect 324044 2 324096 8
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326632 338 326660 598
rect 326816 480 326844 598
rect 327448 546 327500 552
rect 327828 598 328040 626
rect 328256 598 328458 626
rect 327828 542 327856 598
rect 327816 536 327868 542
rect 326620 332 326672 338
rect 326620 274 326672 280
rect 326344 264 326396 270
rect 326048 212 326344 218
rect 326048 206 326396 212
rect 326048 190 326384 206
rect 326774 -960 326886 480
rect 327816 478 327868 484
rect 328012 480 328040 598
rect 328458 575 328514 584
rect 329024 598 329236 626
rect 327970 -960 328082 480
rect 329024 134 329052 598
rect 329208 480 329236 598
rect 330128 598 330432 626
rect 331660 598 331996 626
rect 329748 536 329800 542
rect 329452 484 329748 490
rect 329012 128 329064 134
rect 329012 70 329064 76
rect 329166 -960 329278 480
rect 329452 478 329800 484
rect 329452 462 329788 478
rect 330128 406 330156 598
rect 330404 480 330432 598
rect 330116 400 330168 406
rect 330116 342 330168 348
rect 330362 -960 330474 480
rect 331220 468 331272 474
rect 331220 410 331272 416
rect 331232 354 331260 410
rect 331558 354 331670 480
rect 331968 474 331996 598
rect 332520 598 332732 626
rect 335360 672 335412 678
rect 333612 614 333664 620
rect 331956 468 332008 474
rect 331956 410 332008 416
rect 331232 326 331670 354
rect 330852 128 330904 134
rect 330556 76 330852 82
rect 330556 70 330904 76
rect 330556 54 330892 70
rect 331558 -960 331670 326
rect 332520 66 332548 598
rect 332704 480 332732 598
rect 332508 60 332560 66
rect 332508 2 332560 8
rect 332662 -960 332774 480
rect 333624 354 333652 614
rect 333960 598 334296 626
rect 335064 620 335360 626
rect 338672 672 338724 678
rect 337474 640 337530 649
rect 335064 614 335412 620
rect 335064 598 335400 614
rect 336260 598 336596 626
rect 334268 513 334296 598
rect 334254 504 334310 513
rect 333858 354 333970 480
rect 335280 496 335400 524
rect 334254 439 334310 448
rect 333624 326 333970 354
rect 332856 202 333192 218
rect 332856 196 333204 202
rect 332856 190 333152 196
rect 333152 138 333204 144
rect 333858 -960 333970 326
rect 335054 354 335166 480
rect 335280 354 335308 496
rect 335054 326 335308 354
rect 335054 -960 335166 326
rect 335372 270 335400 496
rect 336250 354 336362 480
rect 336568 406 336596 598
rect 340880 672 340932 678
rect 338672 614 338724 620
rect 340768 620 340880 626
rect 344560 672 344612 678
rect 343362 640 343418 649
rect 340768 614 340932 620
rect 337474 575 337530 584
rect 337488 480 337516 575
rect 338684 480 338712 614
rect 339868 604 339920 610
rect 340768 598 340920 614
rect 340984 598 341196 626
rect 341964 610 342116 626
rect 341964 604 342128 610
rect 341964 598 342076 604
rect 339868 546 339920 552
rect 339880 480 339908 546
rect 340984 480 341012 598
rect 336464 400 336516 406
rect 336250 348 336464 354
rect 336250 342 336516 348
rect 336556 400 336608 406
rect 336556 342 336608 348
rect 336250 326 336504 342
rect 335360 264 335412 270
rect 335360 206 335412 212
rect 336250 -960 336362 326
rect 337212 66 337364 82
rect 337200 60 337364 66
rect 337252 54 337364 60
rect 337200 2 337252 8
rect 337446 -960 337558 480
rect 338302 368 338358 377
rect 338358 326 338468 354
rect 338302 303 338358 312
rect 338642 -960 338754 480
rect 339500 128 339552 134
rect 339552 76 339664 82
rect 339500 70 339664 76
rect 339512 54 339664 70
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 341168 474 341196 598
rect 342076 546 342128 552
rect 342180 598 342392 626
rect 342180 480 342208 598
rect 341156 468 341208 474
rect 341156 410 341208 416
rect 342138 -960 342250 480
rect 342364 202 342392 598
rect 347780 672 347832 678
rect 344560 614 344612 620
rect 345018 640 345074 649
rect 343362 575 343418 584
rect 343068 474 343220 490
rect 343376 480 343404 575
rect 344572 480 344600 614
rect 346950 640 347006 649
rect 345018 575 345074 584
rect 345584 598 345796 626
rect 343068 468 343232 474
rect 343068 462 343180 468
rect 343180 410 343232 416
rect 342352 196 342404 202
rect 342352 138 342404 144
rect 343334 -960 343446 480
rect 344172 338 344416 354
rect 344172 332 344428 338
rect 344172 326 344376 332
rect 344376 274 344428 280
rect 344530 -960 344642 480
rect 345032 66 345060 575
rect 345584 490 345612 598
rect 345492 462 345612 490
rect 345768 480 345796 598
rect 349252 672 349304 678
rect 349066 640 349122 649
rect 347780 614 347832 620
rect 346950 575 347006 584
rect 346964 480 346992 575
rect 345492 406 345520 462
rect 345480 400 345532 406
rect 345480 342 345532 348
rect 345572 264 345624 270
rect 345368 212 345572 218
rect 345368 206 345624 212
rect 345368 190 345612 206
rect 345020 60 345072 66
rect 345020 2 345072 8
rect 345726 -960 345838 480
rect 346472 202 346808 218
rect 346472 196 346820 202
rect 346472 190 346768 196
rect 346768 138 346820 144
rect 346922 -960 347034 480
rect 347792 134 347820 614
rect 347884 598 348096 626
rect 347884 513 347912 598
rect 347870 504 347926 513
rect 348068 480 348096 598
rect 360844 672 360896 678
rect 349252 614 349304 620
rect 350446 640 350502 649
rect 349066 575 349068 584
rect 349120 575 349122 584
rect 349068 546 349120 552
rect 349264 480 349292 614
rect 350446 575 350502 584
rect 350630 640 350686 649
rect 352838 640 352894 649
rect 350980 610 351316 626
rect 350980 604 351328 610
rect 350980 598 351276 604
rect 350630 575 350686 584
rect 350170 504 350226 513
rect 347870 439 347926 448
rect 347780 128 347832 134
rect 347576 66 347728 82
rect 347780 70 347832 76
rect 347576 60 347740 66
rect 347576 54 347688 60
rect 347688 2 347740 8
rect 348026 -960 348138 480
rect 349068 400 349120 406
rect 348772 348 349068 354
rect 348772 342 349120 348
rect 348772 326 349108 342
rect 349222 -960 349334 480
rect 349876 462 350170 490
rect 350460 480 350488 575
rect 350170 439 350226 448
rect 350418 -960 350530 480
rect 350644 474 350672 575
rect 351276 546 351328 552
rect 351472 598 351684 626
rect 351184 536 351236 542
rect 351472 490 351500 598
rect 351236 484 351500 490
rect 351184 478 351500 484
rect 351656 480 351684 598
rect 359922 640 359978 649
rect 352838 575 352894 584
rect 353864 598 354076 626
rect 355580 610 355916 626
rect 352472 536 352524 542
rect 352176 484 352472 490
rect 350632 468 350684 474
rect 351196 462 351500 478
rect 350632 410 350684 416
rect 351614 -960 351726 480
rect 352176 478 352524 484
rect 352852 480 352880 575
rect 352176 462 352512 478
rect 352810 -960 352922 480
rect 353280 474 353616 490
rect 353280 468 353628 474
rect 353280 462 353576 468
rect 353576 410 353628 416
rect 353864 338 353892 598
rect 354048 480 354076 598
rect 355232 604 355284 610
rect 355580 604 355928 610
rect 355580 598 355876 604
rect 355232 546 355284 552
rect 355876 546 355928 552
rect 356164 564 356376 592
rect 355244 480 355272 546
rect 356164 490 356192 564
rect 353852 332 353904 338
rect 353852 274 353904 280
rect 354006 -960 354118 480
rect 354384 338 354720 354
rect 354384 332 354732 338
rect 354384 326 354680 332
rect 354680 274 354732 280
rect 355202 -960 355314 480
rect 356072 462 356192 490
rect 356348 480 356376 564
rect 357360 564 357572 592
rect 356072 202 356100 462
rect 356060 196 356112 202
rect 356060 138 356112 144
rect 356306 -960 356418 480
rect 356684 202 357020 218
rect 356684 196 357032 202
rect 356684 190 356980 196
rect 356980 138 357032 144
rect 357360 66 357388 564
rect 357544 480 357572 564
rect 358464 564 358768 592
rect 369308 672 369360 678
rect 363786 640 363842 649
rect 360844 614 360896 620
rect 359922 575 359978 584
rect 357348 60 357400 66
rect 357348 2 357400 8
rect 357502 -960 357614 480
rect 358464 406 358492 564
rect 358740 480 358768 564
rect 358452 400 358504 406
rect 358452 342 358504 348
rect 358084 128 358136 134
rect 357788 76 358084 82
rect 357788 70 358136 76
rect 357788 54 358124 70
rect 358698 -960 358810 480
rect 358984 474 359320 490
rect 359936 480 359964 575
rect 358984 468 359332 474
rect 358984 462 359280 468
rect 359280 410 359332 416
rect 359894 -960 360006 480
rect 360856 218 360884 614
rect 361192 598 361528 626
rect 362388 598 362724 626
rect 363492 598 363786 626
rect 361090 218 361202 480
rect 361500 377 361528 598
rect 361948 536 362000 542
rect 362696 513 362724 598
rect 364596 598 364932 626
rect 365792 598 366128 626
rect 369196 620 369308 626
rect 371608 672 371660 678
rect 369196 614 369360 620
rect 371496 620 371608 626
rect 374276 672 374328 678
rect 371496 614 371660 620
rect 374090 640 374146 649
rect 363786 575 363842 584
rect 361948 478 362000 484
rect 362682 504 362738 513
rect 361486 368 361542 377
rect 361960 354 361988 478
rect 362286 354 362398 480
rect 362682 439 362738 448
rect 361960 326 362398 354
rect 361486 303 361542 312
rect 360856 190 361202 218
rect 360088 66 360424 82
rect 360088 60 360436 66
rect 360088 54 360384 60
rect 360384 2 360436 8
rect 361090 -960 361202 190
rect 362286 -960 362398 326
rect 363482 354 363594 480
rect 363482 338 363736 354
rect 363482 332 363748 338
rect 363482 326 363696 332
rect 363482 -960 363594 326
rect 363696 274 363748 280
rect 364586 218 364698 480
rect 364904 338 364932 598
rect 366100 542 366128 598
rect 367008 604 367060 610
rect 367008 546 367060 552
rect 368204 604 368256 610
rect 369196 598 369348 614
rect 369400 604 369452 610
rect 368204 546 368256 552
rect 369400 546 369452 552
rect 370596 604 370648 610
rect 371496 598 371648 614
rect 370596 546 370648 552
rect 371712 564 371924 592
rect 366088 536 366140 542
rect 365782 354 365894 480
rect 366088 478 366140 484
rect 366744 474 366896 490
rect 367020 480 367048 546
rect 366732 468 366896 474
rect 366784 462 366896 468
rect 366732 410 366784 416
rect 365996 400 366048 406
rect 365782 348 365996 354
rect 365782 342 366048 348
rect 364892 332 364944 338
rect 364892 274 364944 280
rect 365782 326 366036 342
rect 364800 264 364852 270
rect 364586 212 364800 218
rect 364586 206 364852 212
rect 364586 190 364840 206
rect 364586 -960 364698 190
rect 365782 -960 365894 326
rect 366978 -960 367090 480
rect 367848 474 368000 490
rect 368216 480 368244 546
rect 369412 480 369440 546
rect 370608 480 370636 546
rect 371712 480 371740 564
rect 371896 490 371924 564
rect 372724 564 372936 592
rect 374090 575 374146 584
rect 374274 640 374276 649
rect 375288 672 375340 678
rect 374328 640 374330 649
rect 377956 672 378008 678
rect 375288 614 375340 620
rect 377678 640 377734 649
rect 374274 575 374330 584
rect 372724 513 372752 564
rect 372710 504 372766 513
rect 367836 468 368000 474
rect 367888 462 368000 468
rect 367836 410 367888 416
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370412 128 370464 134
rect 370300 76 370412 82
rect 370300 70 370464 76
rect 370300 54 370452 70
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 371896 462 372016 490
rect 371988 377 372016 462
rect 372908 480 372936 564
rect 373816 536 373868 542
rect 373704 484 373816 490
rect 372710 439 372766 448
rect 371974 368 372030 377
rect 371974 303 372030 312
rect 372712 264 372764 270
rect 372600 212 372712 218
rect 372600 206 372764 212
rect 372600 190 372752 206
rect 372866 -960 372978 480
rect 373704 478 373868 484
rect 374104 480 374132 575
rect 375300 480 375328 614
rect 376484 604 376536 610
rect 377678 575 377734 584
rect 377954 640 377956 649
rect 379520 672 379572 678
rect 378008 640 378010 649
rect 377954 575 378010 584
rect 378704 598 378916 626
rect 379408 620 379520 626
rect 390284 672 390336 678
rect 379408 614 379572 620
rect 379978 640 380034 649
rect 379408 598 379560 614
rect 376484 546 376536 552
rect 375654 504 375710 513
rect 373704 462 373856 478
rect 374062 -960 374174 480
rect 374900 66 375144 82
rect 374900 60 375156 66
rect 374900 54 375104 60
rect 375104 2 375156 8
rect 375258 -960 375370 480
rect 376496 480 376524 546
rect 377692 480 377720 575
rect 378704 513 378732 598
rect 378690 504 378746 513
rect 375654 439 375656 448
rect 375708 439 375710 448
rect 375656 410 375708 416
rect 376300 400 376352 406
rect 376004 348 376300 354
rect 376004 342 376352 348
rect 376004 326 376340 342
rect 376454 -960 376566 480
rect 377108 202 377444 218
rect 377108 196 377456 202
rect 377108 190 377404 196
rect 377404 138 377456 144
rect 377650 -960 377762 480
rect 378304 474 378456 490
rect 378304 468 378468 474
rect 378304 462 378416 468
rect 378888 480 378916 598
rect 379978 575 380034 584
rect 380162 640 380218 649
rect 382370 640 382426 649
rect 380512 610 380848 626
rect 380512 604 380860 610
rect 380512 598 380808 604
rect 380162 575 380164 584
rect 379992 480 380020 575
rect 380216 575 380218 584
rect 380164 546 380216 552
rect 380808 546 380860 552
rect 381004 598 381216 626
rect 380900 536 380952 542
rect 380898 504 380900 513
rect 380952 504 380954 513
rect 378690 439 378746 448
rect 378416 410 378468 416
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 380898 439 380954 448
rect 381004 354 381032 598
rect 381188 480 381216 598
rect 384762 640 384818 649
rect 382812 610 383148 626
rect 382812 604 383160 610
rect 382812 598 383108 604
rect 382370 575 382426 584
rect 382384 480 382412 575
rect 383108 546 383160 552
rect 383396 564 383608 592
rect 385406 640 385462 649
rect 385112 598 385406 626
rect 384762 575 384818 584
rect 388088 598 388300 626
rect 389620 610 389956 626
rect 394240 672 394292 678
rect 390284 614 390336 620
rect 385406 575 385462 584
rect 383396 490 383424 564
rect 380912 326 381032 354
rect 380912 134 380940 326
rect 380900 128 380952 134
rect 380900 70 380952 76
rect 381146 -960 381258 480
rect 381708 338 382044 354
rect 381708 332 382056 338
rect 381708 326 382004 332
rect 382004 274 382056 280
rect 382342 -960 382454 480
rect 383304 462 383424 490
rect 383580 480 383608 564
rect 384776 480 384804 575
rect 385788 564 386000 592
rect 383304 270 383332 462
rect 383292 264 383344 270
rect 383292 206 383344 212
rect 383538 -960 383650 480
rect 384212 128 384264 134
rect 383916 76 384212 82
rect 383916 70 384264 76
rect 383916 54 384252 70
rect 384734 -960 384846 480
rect 385788 354 385816 564
rect 385972 480 386000 564
rect 386984 564 387196 592
rect 385696 326 385816 354
rect 385696 66 385724 326
rect 385684 60 385736 66
rect 385684 2 385736 8
rect 385930 -960 386042 480
rect 386984 406 387012 564
rect 387168 480 387196 564
rect 386972 400 387024 406
rect 386972 342 387024 348
rect 386512 128 386564 134
rect 386216 76 386512 82
rect 386216 70 386564 76
rect 386216 54 386552 70
rect 387126 -960 387238 480
rect 388088 270 388116 598
rect 388272 480 388300 598
rect 389456 604 389508 610
rect 389620 604 389968 610
rect 389620 598 389916 604
rect 389456 546 389508 552
rect 389916 546 389968 552
rect 389468 480 389496 546
rect 388076 264 388128 270
rect 387320 202 387656 218
rect 388076 206 388128 212
rect 387320 196 387668 202
rect 387320 190 387616 196
rect 387616 138 387668 144
rect 388230 -960 388342 480
rect 388812 400 388864 406
rect 388516 348 388812 354
rect 388516 342 388864 348
rect 388516 326 388852 342
rect 389426 -960 389538 480
rect 390296 354 390324 614
rect 390724 598 391060 626
rect 391920 598 392256 626
rect 393024 610 393360 626
rect 395620 672 395672 678
rect 394240 614 394292 620
rect 395324 620 395620 626
rect 401140 672 401192 678
rect 395324 614 395672 620
rect 396538 640 396594 649
rect 390622 354 390734 480
rect 391032 406 391060 598
rect 391572 536 391624 542
rect 391572 478 391624 484
rect 390296 326 390734 354
rect 391020 400 391072 406
rect 391020 342 391072 348
rect 390622 -960 390734 326
rect 391584 218 391612 478
rect 391818 218 391930 480
rect 392228 377 392256 598
rect 392400 604 392452 610
rect 393024 604 393372 610
rect 393024 598 393320 604
rect 392400 546 392452 552
rect 393320 546 393372 552
rect 392412 513 392440 546
rect 392398 504 392454 513
rect 394252 480 394280 614
rect 395324 598 395660 614
rect 396538 575 396594 584
rect 397748 598 397960 626
rect 398728 610 398880 626
rect 398728 604 398892 610
rect 398728 598 398840 604
rect 396552 480 396580 575
rect 397748 480 397776 598
rect 392398 439 392454 448
rect 392214 368 392270 377
rect 392214 303 392270 312
rect 393014 354 393126 480
rect 393014 338 393268 354
rect 393014 332 393280 338
rect 393014 326 393228 332
rect 391584 190 391930 218
rect 391818 -960 391930 190
rect 393014 -960 393126 326
rect 393228 274 393280 280
rect 393964 128 394016 134
rect 394016 76 394128 82
rect 393964 70 394128 76
rect 393976 54 394128 70
rect 394210 -960 394322 480
rect 395314 218 395426 480
rect 395314 190 395568 218
rect 395314 -960 395426 190
rect 395540 66 395568 190
rect 396276 66 396428 82
rect 395528 60 395580 66
rect 395528 2 395580 8
rect 396264 60 396428 66
rect 396316 54 396428 60
rect 396264 2 396316 8
rect 396510 -960 396622 480
rect 397460 128 397512 134
rect 397512 76 397624 82
rect 397460 70 397624 76
rect 397472 54 397624 70
rect 397706 -960 397818 480
rect 397932 270 397960 598
rect 398840 546 398892 552
rect 398944 598 399156 626
rect 398944 480 398972 598
rect 397920 264 397972 270
rect 397920 206 397972 212
rect 398902 -960 399014 480
rect 399128 354 399156 598
rect 399956 598 400168 626
rect 401028 620 401140 626
rect 404728 672 404780 678
rect 401414 640 401470 649
rect 401028 614 401192 620
rect 401028 598 401180 614
rect 401336 598 401414 626
rect 399956 542 399984 598
rect 399944 536 399996 542
rect 399944 478 399996 484
rect 400140 480 400168 598
rect 400312 536 400364 542
rect 399944 400 399996 406
rect 399128 326 399248 354
rect 399832 348 399944 354
rect 399832 342 399996 348
rect 399832 326 399984 342
rect 399220 202 399248 326
rect 399208 196 399260 202
rect 399208 138 399260 144
rect 400098 -960 400210 480
rect 400312 478 400364 484
rect 401336 480 401364 598
rect 403452 598 403664 626
rect 404432 620 404728 626
rect 404912 672 404964 678
rect 404432 614 404780 620
rect 404832 632 404912 660
rect 404432 598 404768 614
rect 401414 575 401470 584
rect 402256 564 402560 592
rect 400324 377 400352 478
rect 400310 368 400366 377
rect 400310 303 400366 312
rect 401294 -960 401406 480
rect 402256 338 402284 564
rect 402532 480 402560 564
rect 403452 542 403480 598
rect 403440 536 403492 542
rect 402244 332 402296 338
rect 402244 274 402296 280
rect 402132 202 402376 218
rect 402132 196 402388 202
rect 402132 190 402336 196
rect 402336 138 402388 144
rect 402490 -960 402602 480
rect 403440 478 403492 484
rect 403636 480 403664 598
rect 404832 480 404860 632
rect 407212 672 407264 678
rect 404912 614 404964 620
rect 405830 640 405886 649
rect 405830 575 405886 584
rect 406028 598 406240 626
rect 413744 672 413796 678
rect 409602 640 409658 649
rect 407212 614 407264 620
rect 403236 338 403480 354
rect 403236 332 403492 338
rect 403236 326 403440 332
rect 403440 274 403492 280
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405094 368 405150 377
rect 405094 303 405150 312
rect 405108 66 405136 303
rect 405536 202 405688 218
rect 405536 196 405700 202
rect 405536 190 405648 196
rect 405648 138 405700 144
rect 405844 134 405872 575
rect 406028 480 406056 598
rect 405832 128 405884 134
rect 405832 70 405884 76
rect 405096 60 405148 66
rect 405096 2 405148 8
rect 405986 -960 406098 480
rect 406212 474 406240 598
rect 407224 480 407252 614
rect 408236 598 408448 626
rect 406200 468 406252 474
rect 406200 410 406252 416
rect 406936 128 406988 134
rect 406640 76 406936 82
rect 406640 70 406988 76
rect 406640 54 406976 70
rect 407182 -960 407294 480
rect 407836 474 408172 490
rect 407836 468 408184 474
rect 407836 462 408132 468
rect 408132 410 408184 416
rect 408236 377 408264 598
rect 408420 480 408448 598
rect 412638 640 412694 649
rect 409602 575 409658 584
rect 410800 604 410852 610
rect 409616 480 409644 575
rect 412344 598 412638 626
rect 410800 546 410852 552
rect 411732 564 411944 592
rect 413448 620 413744 626
rect 413448 614 413796 620
rect 414296 672 414348 678
rect 414296 614 414348 620
rect 415492 672 415544 678
rect 415492 614 415544 620
rect 416688 672 416740 678
rect 417148 672 417200 678
rect 416688 614 416740 620
rect 416852 620 417148 626
rect 418344 672 418396 678
rect 416852 614 417200 620
rect 412638 575 412694 584
rect 413100 604 413152 610
rect 410812 480 410840 546
rect 408222 368 408278 377
rect 408222 303 408278 312
rect 408378 -960 408490 480
rect 408940 338 409276 354
rect 408940 332 409288 338
rect 408940 326 409236 332
rect 409236 274 409288 280
rect 409574 -960 409686 480
rect 410340 264 410392 270
rect 410044 212 410340 218
rect 410044 206 410392 212
rect 410044 190 410380 206
rect 410770 -960 410882 480
rect 411240 474 411576 490
rect 411240 468 411588 474
rect 411240 462 411536 468
rect 411536 410 411588 416
rect 411732 406 411760 564
rect 411916 480 411944 564
rect 413448 598 413784 614
rect 413100 546 413152 552
rect 413112 480 413140 546
rect 414308 480 414336 614
rect 414940 536 414992 542
rect 414644 484 414940 490
rect 411720 400 411772 406
rect 411720 342 411772 348
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 414644 478 414992 484
rect 415504 480 415532 614
rect 416700 480 416728 614
rect 416852 598 417188 614
rect 417712 598 417924 626
rect 418048 620 418344 626
rect 430856 672 430908 678
rect 421746 640 421802 649
rect 418048 614 418396 620
rect 418048 598 418384 614
rect 418816 598 419028 626
rect 414644 462 414980 478
rect 415462 -960 415574 480
rect 416044 400 416096 406
rect 415748 348 416044 354
rect 415748 342 416096 348
rect 415748 326 416084 342
rect 416658 -960 416770 480
rect 417712 134 417740 598
rect 417896 480 417924 598
rect 417700 128 417752 134
rect 417700 70 417752 76
rect 417854 -960 417966 480
rect 418816 66 418844 598
rect 419000 480 419028 598
rect 419908 604 419960 610
rect 420256 598 420592 626
rect 421452 610 421696 626
rect 421452 604 421708 610
rect 421452 598 421656 604
rect 419908 546 419960 552
rect 418804 60 418856 66
rect 418804 2 418856 8
rect 418958 -960 419070 480
rect 419448 264 419500 270
rect 419152 212 419448 218
rect 419152 206 419500 212
rect 419920 218 419948 546
rect 420154 218 420266 480
rect 420564 474 420592 598
rect 427266 640 427322 649
rect 422556 610 422892 626
rect 424704 610 424856 626
rect 422556 604 422904 610
rect 422556 598 422852 604
rect 421746 575 421802 584
rect 421656 546 421708 552
rect 421760 542 421788 575
rect 422852 546 422904 552
rect 423772 604 423824 610
rect 423772 546 423824 552
rect 424692 604 424856 610
rect 424744 598 424856 604
rect 424968 604 425020 610
rect 424692 546 424744 552
rect 424968 546 425020 552
rect 426176 598 426388 626
rect 421748 536 421800 542
rect 420552 468 420604 474
rect 420552 410 420604 416
rect 421350 354 421462 480
rect 421748 478 421800 484
rect 423784 480 423812 546
rect 424508 536 424560 542
rect 424506 504 424508 513
rect 424560 504 424562 513
rect 421024 338 421462 354
rect 421012 332 421462 338
rect 421064 326 421462 332
rect 421012 274 421064 280
rect 419152 190 419488 206
rect 419920 190 420266 218
rect 420154 -960 420266 190
rect 421350 -960 421462 326
rect 422546 218 422658 480
rect 423508 338 423660 354
rect 423496 332 423660 338
rect 423548 326 423660 332
rect 423496 274 423548 280
rect 422546 202 422800 218
rect 422546 196 422812 202
rect 422546 190 422760 196
rect 422546 -960 422658 190
rect 422760 138 422812 144
rect 423742 -960 423854 480
rect 424980 480 425008 546
rect 426176 480 426204 598
rect 426360 542 426388 598
rect 429014 640 429070 649
rect 427266 575 427322 584
rect 428476 598 428688 626
rect 426348 536 426400 542
rect 424506 439 424562 448
rect 424938 -960 425050 480
rect 425808 66 425960 82
rect 425796 60 425960 66
rect 425848 54 425960 60
rect 425796 2 425848 8
rect 426134 -960 426246 480
rect 426348 478 426400 484
rect 427280 480 427308 575
rect 428476 480 428504 598
rect 427004 202 427156 218
rect 426992 196 427156 202
rect 427044 190 427156 196
rect 426992 138 427044 144
rect 427238 -960 427350 480
rect 428096 128 428148 134
rect 428148 76 428260 82
rect 428096 70 428260 76
rect 428108 54 428260 70
rect 428434 -960 428546 480
rect 428660 406 428688 598
rect 429014 575 429070 584
rect 429658 640 429714 649
rect 434444 672 434496 678
rect 430856 614 430908 620
rect 429658 575 429714 584
rect 429028 542 429056 575
rect 429016 536 429068 542
rect 429476 536 429528 542
rect 429016 478 429068 484
rect 429364 484 429476 490
rect 429364 478 429528 484
rect 429672 480 429700 575
rect 429364 462 429516 478
rect 428648 400 428700 406
rect 428648 342 428700 348
rect 429630 -960 429742 480
rect 430408 474 430560 490
rect 430868 480 430896 614
rect 431880 598 432092 626
rect 435180 672 435232 678
rect 434444 614 434496 620
rect 435068 620 435180 626
rect 436468 672 436520 678
rect 435068 614 435232 620
rect 436172 620 436468 626
rect 437940 672 437992 678
rect 436172 614 436520 620
rect 430396 468 430560 474
rect 430448 462 430560 468
rect 430396 410 430448 416
rect 430826 -960 430938 480
rect 431880 354 431908 598
rect 432064 480 432092 598
rect 433248 604 433300 610
rect 433248 546 433300 552
rect 433260 480 433288 546
rect 431788 326 431908 354
rect 431788 270 431816 326
rect 431776 264 431828 270
rect 431776 206 431828 212
rect 431868 128 431920 134
rect 431664 76 431868 82
rect 431664 70 431920 76
rect 431664 54 431908 70
rect 432022 -960 432134 480
rect 432768 338 433104 354
rect 432768 332 433116 338
rect 432768 326 433064 332
rect 433064 274 433116 280
rect 433218 -960 433330 480
rect 433964 474 434300 490
rect 434456 480 434484 614
rect 435068 598 435220 614
rect 435548 604 435600 610
rect 436172 598 436508 614
rect 436572 598 436784 626
rect 442632 672 442684 678
rect 437940 614 437992 620
rect 435548 546 435600 552
rect 435560 480 435588 546
rect 433964 468 434312 474
rect 433964 462 434260 468
rect 434260 410 434312 416
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436468 400 436520 406
rect 436572 354 436600 598
rect 436756 480 436784 598
rect 437952 480 437980 614
rect 441876 610 442212 626
rect 448244 672 448296 678
rect 442632 614 442684 620
rect 441528 604 441580 610
rect 438964 564 439176 592
rect 436520 348 436600 354
rect 436468 342 436600 348
rect 436480 326 436600 342
rect 436714 -960 436826 480
rect 437480 400 437532 406
rect 437368 348 437480 354
rect 437368 342 437532 348
rect 437368 326 437520 342
rect 437910 -960 438022 480
rect 438964 354 438992 564
rect 439148 480 439176 564
rect 440160 564 440372 592
rect 438872 326 438992 354
rect 438768 264 438820 270
rect 438472 212 438768 218
rect 438472 206 438820 212
rect 438472 190 438808 206
rect 438872 66 438900 326
rect 438860 60 438912 66
rect 438860 2 438912 8
rect 439106 -960 439218 480
rect 440160 202 440188 564
rect 440344 480 440372 564
rect 441876 604 442224 610
rect 441876 598 442172 604
rect 441528 546 441580 552
rect 442172 546 442224 552
rect 441540 480 441568 546
rect 442644 480 442672 614
rect 444176 610 444512 626
rect 443828 604 443880 610
rect 444176 604 444524 610
rect 444176 598 444472 604
rect 443828 546 443880 552
rect 446048 598 446260 626
rect 444472 546 444524 552
rect 444852 564 445064 592
rect 443276 536 443328 542
rect 442980 484 443276 490
rect 440148 196 440200 202
rect 440148 138 440200 144
rect 439576 66 439912 82
rect 439576 60 439924 66
rect 439576 54 439872 60
rect 439872 2 439924 8
rect 440302 -960 440414 480
rect 440772 202 441108 218
rect 440772 196 441120 202
rect 440772 190 441068 196
rect 441068 138 441120 144
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 442980 478 443328 484
rect 443840 480 443868 546
rect 444852 490 444880 564
rect 442980 462 443316 478
rect 443798 -960 443910 480
rect 444760 462 444880 490
rect 445036 480 445064 564
rect 444760 134 444788 462
rect 444748 128 444800 134
rect 444748 70 444800 76
rect 444994 -960 445106 480
rect 446048 338 446076 598
rect 446232 480 446260 598
rect 447152 598 447456 626
rect 448980 672 449032 678
rect 448244 614 448296 620
rect 448684 620 448980 626
rect 456892 672 456944 678
rect 456062 640 456118 649
rect 448684 614 449032 620
rect 446036 332 446088 338
rect 446036 274 446088 280
rect 445576 128 445628 134
rect 445280 76 445576 82
rect 445280 70 445628 76
rect 445280 54 445616 70
rect 446190 -960 446302 480
rect 447152 474 447180 598
rect 447428 480 447456 598
rect 447140 468 447192 474
rect 447140 410 447192 416
rect 446678 368 446734 377
rect 446384 326 446678 354
rect 446678 303 446734 312
rect 447386 -960 447498 480
rect 448256 354 448284 614
rect 448684 598 449020 614
rect 449636 598 449788 626
rect 449866 610 450032 626
rect 450984 610 451320 626
rect 452088 610 452424 626
rect 449866 604 450044 610
rect 449866 598 449992 604
rect 448582 354 448694 480
rect 448256 326 448694 354
rect 447876 264 447928 270
rect 447580 212 447876 218
rect 447580 206 447928 212
rect 447580 190 447916 206
rect 448582 -960 448694 326
rect 449636 66 449664 598
rect 449866 480 449894 598
rect 450984 604 451332 610
rect 450984 598 451280 604
rect 449992 546 450044 552
rect 452088 604 452436 610
rect 452088 598 452384 604
rect 451280 546 451332 552
rect 453284 598 453620 626
rect 452384 546 452436 552
rect 453592 542 453620 598
rect 454500 604 454552 610
rect 454500 546 454552 552
rect 455696 604 455748 610
rect 457996 672 458048 678
rect 456892 614 456944 620
rect 457792 620 457996 626
rect 458180 672 458232 678
rect 457792 614 458048 620
rect 458100 620 458180 626
rect 460204 672 460256 678
rect 458100 614 458232 620
rect 460092 620 460204 626
rect 462780 672 462832 678
rect 460092 614 460256 620
rect 460478 640 460534 649
rect 456062 575 456118 584
rect 455696 546 455748 552
rect 453488 536 453540 542
rect 449778 326 449894 480
rect 450636 400 450688 406
rect 450882 354 450994 480
rect 450688 348 450994 354
rect 450636 342 450994 348
rect 450648 326 450994 342
rect 449624 60 449676 66
rect 449624 2 449676 8
rect 449778 -960 449890 326
rect 450882 -960 450994 326
rect 451922 368 451978 377
rect 451922 303 451924 312
rect 451976 303 451978 312
rect 452078 354 452190 480
rect 452292 400 452344 406
rect 452078 348 452292 354
rect 452078 342 452344 348
rect 453274 354 453386 480
rect 453488 478 453540 484
rect 453580 536 453632 542
rect 453580 478 453632 484
rect 454512 480 454540 546
rect 453500 354 453528 478
rect 452078 326 452332 342
rect 453274 326 453528 354
rect 454224 400 454276 406
rect 454276 348 454388 354
rect 454224 342 454388 348
rect 454236 326 454388 342
rect 451924 274 451976 280
rect 452078 -960 452190 326
rect 453274 -960 453386 326
rect 454470 -960 454582 480
rect 455340 474 455492 490
rect 455708 480 455736 546
rect 455328 468 455492 474
rect 455380 462 455492 468
rect 455328 410 455380 416
rect 455666 -960 455778 480
rect 456076 338 456104 575
rect 456536 474 456688 490
rect 456904 480 456932 614
rect 457792 598 458036 614
rect 458100 598 458220 614
rect 459192 604 459244 610
rect 458100 480 458128 598
rect 460092 598 460244 614
rect 459192 546 459244 552
rect 460400 584 460478 592
rect 462134 640 462190 649
rect 460400 575 460534 584
rect 461320 598 461624 626
rect 460400 564 460520 575
rect 459204 480 459232 546
rect 460400 480 460428 564
rect 456524 468 456688 474
rect 456576 462 456688 468
rect 456524 410 456576 416
rect 456064 332 456116 338
rect 456064 274 456116 280
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459008 128 459060 134
rect 458896 76 459008 82
rect 458896 70 459060 76
rect 458896 54 459048 70
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461044 338 461196 354
rect 461032 332 461196 338
rect 461084 326 461196 332
rect 461032 274 461084 280
rect 461320 270 461348 598
rect 461596 480 461624 598
rect 466276 672 466328 678
rect 462780 614 462832 620
rect 463974 640 464030 649
rect 462134 575 462190 584
rect 461308 264 461360 270
rect 461308 206 461360 212
rect 461554 -960 461666 480
rect 462148 66 462176 575
rect 462792 480 462820 614
rect 466090 640 466146 649
rect 463974 575 464030 584
rect 465172 604 465224 610
rect 463988 480 464016 575
rect 471060 672 471112 678
rect 466276 614 466328 620
rect 467470 640 467526 649
rect 466090 575 466146 584
rect 465172 546 465224 552
rect 465184 480 465212 546
rect 466104 542 466132 575
rect 466092 536 466144 542
rect 462300 202 462452 218
rect 462300 196 462464 202
rect 462300 190 462412 196
rect 462412 138 462464 144
rect 462136 60 462188 66
rect 462136 2 462188 8
rect 462750 -960 462862 480
rect 463608 264 463660 270
rect 463496 212 463608 218
rect 463496 206 463660 212
rect 463496 190 463648 206
rect 463946 -960 464058 480
rect 464600 66 464936 82
rect 464600 60 464948 66
rect 464600 54 464896 60
rect 464896 2 464948 8
rect 465142 -960 465254 480
rect 466092 478 466144 484
rect 466288 480 466316 614
rect 470598 640 470654 649
rect 469864 604 469916 610
rect 467470 575 467526 584
rect 467196 536 467248 542
rect 466900 484 467196 490
rect 466000 400 466052 406
rect 465704 348 466000 354
rect 465704 342 466052 348
rect 465704 326 466040 342
rect 466246 -960 466358 480
rect 466900 478 467248 484
rect 467484 480 467512 575
rect 468496 564 468708 592
rect 468298 504 468354 513
rect 466900 462 467236 478
rect 467442 -960 467554 480
rect 468004 462 468298 490
rect 468496 474 468524 564
rect 468680 480 468708 564
rect 470304 598 470598 626
rect 471704 672 471756 678
rect 471060 614 471112 620
rect 471408 620 471704 626
rect 471408 614 471756 620
rect 472256 672 472308 678
rect 472808 672 472860 678
rect 472256 614 472308 620
rect 472512 620 472808 626
rect 474556 672 474608 678
rect 472512 614 472860 620
rect 470598 575 470654 584
rect 469864 546 469916 552
rect 468298 439 468354 448
rect 468484 468 468536 474
rect 468484 410 468536 416
rect 468638 -960 468750 480
rect 469108 474 469260 490
rect 469876 480 469904 546
rect 471072 480 471100 614
rect 471408 598 471744 614
rect 472268 480 472296 614
rect 472512 598 472848 614
rect 473280 598 473492 626
rect 480720 672 480772 678
rect 477406 640 477462 649
rect 474556 614 474608 620
rect 469108 468 469272 474
rect 469108 462 469220 468
rect 469220 410 469272 416
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473280 134 473308 598
rect 473464 480 473492 598
rect 474568 480 474596 614
rect 474812 610 475148 626
rect 474812 604 475160 610
rect 474812 598 475108 604
rect 475108 546 475160 552
rect 475580 598 475792 626
rect 475916 610 476252 626
rect 475916 604 476264 610
rect 475916 598 476212 604
rect 475580 490 475608 598
rect 473268 128 473320 134
rect 473268 70 473320 76
rect 473422 -960 473534 480
rect 474004 128 474056 134
rect 473708 76 474004 82
rect 473708 70 474056 76
rect 473708 54 474044 70
rect 474526 -960 474638 480
rect 475488 462 475608 490
rect 475764 480 475792 598
rect 476212 546 476264 552
rect 476580 604 476632 610
rect 476580 546 476632 552
rect 476684 598 476988 626
rect 476592 513 476620 546
rect 476578 504 476634 513
rect 475488 270 475516 462
rect 475476 264 475528 270
rect 475476 206 475528 212
rect 475722 -960 475834 480
rect 476578 439 476634 448
rect 476684 202 476712 598
rect 476960 480 476988 598
rect 477406 575 477462 584
rect 477868 604 477920 610
rect 477420 542 477448 575
rect 478216 598 478552 626
rect 479320 598 479656 626
rect 480516 610 480668 626
rect 480720 614 480772 620
rect 481456 672 481508 678
rect 483756 672 483808 678
rect 483202 640 483258 649
rect 481508 620 481620 626
rect 481456 614 481620 620
rect 480516 604 480680 610
rect 480516 598 480628 604
rect 477868 546 477920 552
rect 477408 536 477460 542
rect 476672 196 476724 202
rect 476672 138 476724 144
rect 476918 -960 477030 480
rect 477408 478 477460 484
rect 477880 218 477908 546
rect 478114 218 478226 480
rect 478524 270 478552 598
rect 477112 202 477448 218
rect 477112 196 477460 202
rect 477112 190 477408 196
rect 477880 190 478226 218
rect 478512 264 478564 270
rect 478512 206 478564 212
rect 477408 138 477460 144
rect 478114 -960 478226 190
rect 479310 82 479422 480
rect 479628 406 479656 598
rect 480628 546 480680 552
rect 479616 400 479668 406
rect 479616 342 479668 348
rect 480506 354 480618 480
rect 480732 354 480760 614
rect 481468 598 481620 614
rect 481732 604 481784 610
rect 481732 546 481784 552
rect 482664 598 482816 626
rect 481744 480 481772 546
rect 480506 326 480760 354
rect 479310 66 479564 82
rect 479310 60 479576 66
rect 479310 54 479524 60
rect 479310 -960 479422 54
rect 479524 2 479576 8
rect 480506 -960 480618 326
rect 481702 -960 481814 480
rect 482664 66 482692 598
rect 485228 672 485280 678
rect 483808 620 483920 626
rect 483756 614 483920 620
rect 487712 672 487764 678
rect 485228 614 485280 620
rect 483768 598 483920 614
rect 484032 604 484084 610
rect 483202 575 483258 584
rect 482806 218 482918 480
rect 482974 332 483026 338
rect 482974 274 483026 280
rect 482986 218 483014 274
rect 482806 190 483014 218
rect 482652 60 482704 66
rect 482652 2 482704 8
rect 482806 -960 482918 190
rect 483216 134 483244 575
rect 484032 546 484084 552
rect 484044 480 484072 546
rect 485240 480 485268 614
rect 487324 610 487476 626
rect 487632 620 487712 626
rect 489920 672 489972 678
rect 487632 614 487764 620
rect 488814 640 488870 649
rect 486424 604 486476 610
rect 487324 604 487488 610
rect 487324 598 487436 604
rect 486424 546 486476 552
rect 487436 546 487488 552
rect 487632 598 487752 614
rect 486436 480 486464 546
rect 487632 480 487660 598
rect 489920 614 489972 620
rect 491116 672 491168 678
rect 491300 672 491352 678
rect 491116 614 491168 620
rect 491298 640 491300 649
rect 493324 672 493376 678
rect 491352 640 491354 649
rect 488814 575 488870 584
rect 488828 480 488856 575
rect 489736 536 489788 542
rect 489624 484 489736 490
rect 483662 232 483718 241
rect 483662 167 483664 176
rect 483716 167 483718 176
rect 483664 138 483716 144
rect 483204 128 483256 134
rect 483204 70 483256 76
rect 484002 -960 484114 480
rect 484872 338 485024 354
rect 484860 332 485024 338
rect 484912 326 485024 332
rect 484860 274 484912 280
rect 485198 -960 485310 480
rect 486068 202 486220 218
rect 486056 196 486220 202
rect 486108 190 486220 196
rect 486056 138 486108 144
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488540 128 488592 134
rect 488428 76 488540 82
rect 488428 70 488592 76
rect 488428 54 488580 70
rect 488786 -960 488898 480
rect 489624 478 489788 484
rect 489932 480 489960 614
rect 489624 462 489776 478
rect 489890 -960 490002 480
rect 490728 474 490972 490
rect 491128 480 491156 614
rect 491832 610 492168 626
rect 494428 672 494480 678
rect 493324 614 493376 620
rect 491832 604 492180 610
rect 491832 598 492128 604
rect 491298 575 491354 584
rect 492128 546 492180 552
rect 492324 564 492536 592
rect 492324 480 492352 564
rect 490728 468 490984 474
rect 490728 462 490932 468
rect 490932 410 490984 416
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 492508 241 492536 564
rect 493336 513 493364 614
rect 493520 598 493732 626
rect 494132 620 494428 626
rect 502984 672 503036 678
rect 495898 640 495954 649
rect 494132 614 494480 620
rect 494132 598 494468 614
rect 494532 598 494744 626
rect 495236 610 495388 626
rect 495236 604 495400 610
rect 495236 598 495348 604
rect 493322 504 493378 513
rect 493520 480 493548 598
rect 493704 490 493732 598
rect 494532 490 494560 598
rect 493322 439 493378 448
rect 493324 400 493376 406
rect 492678 368 492734 377
rect 493028 348 493324 354
rect 493028 342 493376 348
rect 493028 326 493364 342
rect 492678 303 492734 312
rect 492692 270 492720 303
rect 492680 264 492732 270
rect 492494 232 492550 241
rect 492680 206 492732 212
rect 492494 167 492550 176
rect 493478 -960 493590 480
rect 493704 462 493824 490
rect 493796 377 493824 462
rect 494440 462 494560 490
rect 494716 480 494744 598
rect 498014 640 498070 649
rect 496432 610 496768 626
rect 496432 604 496780 610
rect 496432 598 496728 604
rect 495898 575 495954 584
rect 495348 546 495400 552
rect 495912 480 495940 575
rect 496728 546 496780 552
rect 497094 606 497150 615
rect 500590 640 500646 649
rect 499836 610 500172 626
rect 498014 575 498070 584
rect 498200 604 498252 610
rect 497094 541 497150 550
rect 497108 480 497136 541
rect 493782 368 493838 377
rect 493782 303 493838 312
rect 494440 270 494468 462
rect 494428 264 494480 270
rect 494428 206 494480 212
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498028 338 498056 575
rect 498200 546 498252 552
rect 499396 604 499448 610
rect 499836 604 500184 610
rect 499836 598 500132 604
rect 499396 546 499448 552
rect 500590 575 500646 584
rect 501616 598 501828 626
rect 505744 672 505796 678
rect 502984 614 503036 620
rect 500132 546 500184 552
rect 498212 480 498240 546
rect 499408 480 499436 546
rect 500604 480 500632 575
rect 498016 332 498068 338
rect 498016 274 498068 280
rect 497832 264 497884 270
rect 497536 212 497832 218
rect 497536 206 497884 212
rect 497536 190 497872 206
rect 498170 -960 498282 480
rect 498640 66 498976 82
rect 498640 60 498988 66
rect 498640 54 498936 60
rect 498936 2 498988 8
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 500940 338 501276 354
rect 500940 332 501288 338
rect 500940 326 501236 332
rect 501236 274 501288 280
rect 501616 202 501644 598
rect 501800 480 501828 598
rect 501604 196 501656 202
rect 501604 138 501656 144
rect 501758 -960 501870 480
rect 502044 474 502380 490
rect 502996 480 503024 614
rect 504008 598 504220 626
rect 505448 620 505744 626
rect 505448 614 505796 620
rect 506480 672 506532 678
rect 506940 672 506992 678
rect 506480 614 506532 620
rect 506644 620 506940 626
rect 509240 672 509292 678
rect 506644 614 506992 620
rect 505448 598 505784 614
rect 502044 468 502392 474
rect 502044 462 502340 468
rect 502340 410 502392 416
rect 502954 -960 503066 480
rect 503240 474 503576 490
rect 503240 468 503588 474
rect 503240 462 503536 468
rect 503536 410 503588 416
rect 504008 134 504036 598
rect 504192 480 504220 598
rect 505100 536 505152 542
rect 503996 128 504048 134
rect 503996 70 504048 76
rect 504150 -960 504262 480
rect 505100 478 505152 484
rect 506492 480 506520 614
rect 506644 598 506980 614
rect 507748 598 507900 626
rect 508944 620 509240 626
rect 508944 614 509292 620
rect 509700 672 509752 678
rect 511264 672 511316 678
rect 509700 614 509752 620
rect 508944 598 509280 614
rect 507308 536 507360 542
rect 505112 218 505140 478
rect 505346 218 505458 480
rect 505112 190 505458 218
rect 504640 128 504692 134
rect 504344 76 504640 82
rect 504344 70 504692 76
rect 504344 54 504680 70
rect 505346 -960 505458 190
rect 506450 -960 506562 480
rect 507308 478 507360 484
rect 507320 354 507348 478
rect 507646 354 507758 480
rect 507320 326 507758 354
rect 507646 -960 507758 326
rect 507872 202 507900 598
rect 509712 513 509740 614
rect 510048 598 510384 626
rect 511264 614 511316 620
rect 512460 672 512512 678
rect 512460 614 512512 620
rect 513288 672 513340 678
rect 515864 672 515916 678
rect 514666 640 514722 649
rect 513340 620 513452 626
rect 513288 614 513452 620
rect 509698 504 509754 513
rect 508688 400 508740 406
rect 508594 368 508650 377
rect 508842 354 508954 480
rect 509698 439 509754 448
rect 508740 348 508954 354
rect 508688 342 508954 348
rect 508700 326 508954 342
rect 508594 303 508596 312
rect 508648 303 508650 312
rect 508596 274 508648 280
rect 507860 196 507912 202
rect 507860 138 507912 144
rect 508842 -960 508954 326
rect 510038 354 510150 480
rect 510252 400 510304 406
rect 510038 348 510252 354
rect 510038 342 510304 348
rect 510038 326 510292 342
rect 510356 338 510384 598
rect 511276 480 511304 614
rect 512184 536 512236 542
rect 512236 484 512348 490
rect 510988 400 511040 406
rect 511040 348 511152 354
rect 510988 342 511152 348
rect 510344 332 510396 338
rect 510038 -960 510150 326
rect 511000 326 511152 342
rect 510344 274 510396 280
rect 511234 -960 511346 480
rect 512184 478 512348 484
rect 512472 480 512500 614
rect 513300 598 513452 614
rect 513576 598 513788 626
rect 514556 598 514666 626
rect 513576 480 513604 598
rect 513760 524 513788 598
rect 514666 575 514722 584
rect 514772 598 514984 626
rect 515752 620 515864 626
rect 517060 672 517112 678
rect 515752 614 515916 620
rect 515752 598 515904 614
rect 515968 610 516180 626
rect 516856 620 517060 626
rect 519360 672 519412 678
rect 518346 640 518402 649
rect 516856 614 517112 620
rect 515968 604 516192 610
rect 515968 598 516140 604
rect 513760 496 513880 524
rect 512196 462 512348 478
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 513852 270 513880 496
rect 514772 480 514800 598
rect 513840 264 513892 270
rect 513840 206 513892 212
rect 514730 -960 514842 480
rect 514956 66 514984 598
rect 515968 480 515996 598
rect 516856 598 517100 614
rect 517960 610 518204 626
rect 517960 604 518216 610
rect 517960 598 518164 604
rect 516140 546 516192 552
rect 517164 564 517376 592
rect 517164 480 517192 564
rect 514944 60 514996 66
rect 514944 2 514996 8
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 517348 377 517376 564
rect 519156 620 519360 626
rect 521844 672 521896 678
rect 519156 614 519412 620
rect 519156 598 519400 614
rect 519556 598 519768 626
rect 518346 575 518402 584
rect 518164 546 518216 552
rect 518360 480 518388 575
rect 519556 480 519584 598
rect 517334 368 517390 377
rect 517334 303 517390 312
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 519740 474 519768 598
rect 520568 598 520780 626
rect 521844 614 521896 620
rect 523040 672 523092 678
rect 523960 672 524012 678
rect 523040 614 523092 620
rect 523664 620 523960 626
rect 532516 672 532568 678
rect 531318 640 531374 649
rect 523664 614 524012 620
rect 519728 468 519780 474
rect 519728 410 519780 416
rect 520260 338 520412 354
rect 520260 332 520424 338
rect 520260 326 520372 332
rect 520372 274 520424 280
rect 520568 134 520596 598
rect 520752 480 520780 598
rect 521856 480 521884 614
rect 523052 480 523080 614
rect 523664 598 524000 614
rect 524064 598 524276 626
rect 520556 128 520608 134
rect 520556 70 520608 76
rect 520710 -960 520822 480
rect 521364 66 521608 82
rect 521364 60 521620 66
rect 521364 54 521568 60
rect 521568 2 521620 8
rect 521814 -960 521926 480
rect 522856 128 522908 134
rect 522560 76 522856 82
rect 522560 70 522908 76
rect 522560 54 522896 70
rect 523010 -960 523122 480
rect 524064 202 524092 598
rect 524248 480 524276 598
rect 525168 598 525472 626
rect 524052 196 524104 202
rect 524052 138 524104 144
rect 524206 -960 524318 480
rect 524768 474 525104 490
rect 525168 474 525196 598
rect 525444 480 525472 598
rect 526456 598 526668 626
rect 524768 468 525116 474
rect 524768 462 525064 468
rect 525064 410 525116 416
rect 525156 468 525208 474
rect 525156 410 525208 416
rect 525402 -960 525514 480
rect 526456 270 526484 598
rect 526640 480 526668 598
rect 527652 598 527864 626
rect 526444 264 526496 270
rect 525964 202 526300 218
rect 526444 206 526496 212
rect 525964 196 526312 202
rect 525964 190 526260 196
rect 526260 138 526312 144
rect 526598 -960 526710 480
rect 527652 406 527680 598
rect 527836 480 527864 598
rect 529020 604 529072 610
rect 529020 546 529072 552
rect 530124 604 530176 610
rect 531576 610 531912 626
rect 533068 672 533120 678
rect 532516 614 532568 620
rect 532772 620 533068 626
rect 535828 672 535880 678
rect 532772 614 533120 620
rect 531576 604 531924 610
rect 531576 598 531872 604
rect 531318 575 531374 584
rect 530124 546 530176 552
rect 529032 480 529060 546
rect 529664 536 529716 542
rect 529368 484 529664 490
rect 527640 400 527692 406
rect 527178 368 527234 377
rect 527068 326 527178 354
rect 527640 342 527692 348
rect 527178 303 527234 312
rect 527794 -960 527906 480
rect 528468 400 528520 406
rect 528172 348 528468 354
rect 528172 342 528520 348
rect 528172 326 528508 342
rect 528990 -960 529102 480
rect 529368 478 529716 484
rect 530136 480 530164 546
rect 531332 480 531360 575
rect 531872 546 531924 552
rect 532528 480 532556 614
rect 532772 598 533108 614
rect 533712 604 533764 610
rect 534980 598 535316 626
rect 536472 672 536524 678
rect 535828 614 535880 620
rect 536176 620 536472 626
rect 540796 672 540848 678
rect 536176 614 536524 620
rect 533712 546 533764 552
rect 533724 480 533752 546
rect 529368 462 529704 478
rect 530094 -960 530206 480
rect 530766 96 530822 105
rect 530472 54 530766 82
rect 530766 31 530822 40
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534540 468 534592 474
rect 534540 410 534592 416
rect 534552 354 534580 410
rect 534878 354 534990 480
rect 534552 326 534990 354
rect 534170 232 534226 241
rect 533876 190 534170 218
rect 534170 167 534226 176
rect 534878 -960 534990 326
rect 535288 202 535316 598
rect 535840 218 535868 614
rect 536176 598 536512 614
rect 537280 598 537616 626
rect 538476 598 538812 626
rect 539580 598 539916 626
rect 542176 672 542228 678
rect 540796 614 540848 620
rect 541714 640 541770 649
rect 536074 218 536186 480
rect 537178 354 537290 480
rect 536944 338 537290 354
rect 537588 338 537616 598
rect 538784 542 538812 598
rect 538772 536 538824 542
rect 536932 332 537290 338
rect 536984 326 537290 332
rect 536932 274 536984 280
rect 535276 196 535328 202
rect 535840 190 536186 218
rect 535276 138 535328 144
rect 536074 -960 536186 190
rect 537178 -960 537290 326
rect 537576 332 537628 338
rect 537576 274 537628 280
rect 538374 82 538486 480
rect 538772 478 538824 484
rect 538048 66 538486 82
rect 538036 60 538486 66
rect 538088 54 538486 60
rect 538036 2 538088 8
rect 538374 -960 538486 54
rect 539570 82 539682 480
rect 539784 128 539836 134
rect 539570 76 539784 82
rect 539570 70 539836 76
rect 539570 54 539824 70
rect 539888 66 539916 598
rect 540518 504 540574 513
rect 540574 462 540684 490
rect 540808 480 540836 614
rect 541770 598 541880 626
rect 542004 620 542176 626
rect 543188 672 543240 678
rect 543094 640 543150 649
rect 542004 614 542228 620
rect 542004 598 542216 614
rect 542984 598 543094 626
rect 541714 575 541770 584
rect 542004 480 542032 598
rect 545488 672 545540 678
rect 543188 614 543240 620
rect 543462 640 543518 649
rect 543094 575 543150 584
rect 543200 480 543228 614
rect 543462 575 543518 584
rect 544396 598 544608 626
rect 553768 672 553820 678
rect 545488 614 545540 620
rect 540518 439 540574 448
rect 539876 60 539928 66
rect 539570 -960 539682 54
rect 539876 2 539928 8
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 543476 338 543504 575
rect 544396 480 544424 598
rect 543464 332 543516 338
rect 543464 274 543516 280
rect 544200 264 544252 270
rect 544088 212 544200 218
rect 544088 206 544252 212
rect 544088 190 544240 206
rect 544354 -960 544466 480
rect 544580 377 544608 598
rect 545500 480 545528 614
rect 546512 598 546724 626
rect 544566 368 544622 377
rect 545132 338 545284 354
rect 544566 303 544622 312
rect 545120 332 545284 338
rect 545172 326 545284 332
rect 545120 274 545172 280
rect 545458 -960 545570 480
rect 546512 474 546540 598
rect 546696 480 546724 598
rect 547892 598 548104 626
rect 546500 468 546552 474
rect 546500 410 546552 416
rect 546500 128 546552 134
rect 546388 76 546500 82
rect 546388 70 546552 76
rect 546388 54 546540 70
rect 546654 -960 546766 480
rect 547492 474 547736 490
rect 547892 480 547920 598
rect 547492 468 547748 474
rect 547492 462 547696 468
rect 547696 410 547748 416
rect 547850 -960 547962 480
rect 548076 105 548104 598
rect 549088 598 549300 626
rect 550896 610 551232 626
rect 548892 536 548944 542
rect 548688 484 548892 490
rect 548688 478 548944 484
rect 549088 480 549116 598
rect 549272 542 549300 598
rect 550272 604 550324 610
rect 550896 604 551244 610
rect 550896 598 551192 604
rect 550272 546 550324 552
rect 551192 546 551244 552
rect 551296 598 551508 626
rect 552092 610 552428 626
rect 552092 604 552440 610
rect 552092 598 552388 604
rect 549260 536 549312 542
rect 550088 536 550140 542
rect 548688 462 548932 478
rect 548062 96 548118 105
rect 548062 31 548118 40
rect 549046 -960 549158 480
rect 549260 478 549312 484
rect 549792 484 550088 490
rect 549792 478 550140 484
rect 550284 480 550312 546
rect 549792 462 550128 478
rect 550242 -960 550354 480
rect 551296 241 551324 598
rect 551480 480 551508 598
rect 552388 546 552440 552
rect 552492 598 552704 626
rect 555148 672 555200 678
rect 553768 614 553820 620
rect 554962 640 555018 649
rect 552492 490 552520 598
rect 551282 232 551338 241
rect 551282 167 551338 176
rect 551438 -960 551550 480
rect 552400 462 552520 490
rect 552676 480 552704 598
rect 553780 480 553808 614
rect 554962 575 555018 584
rect 555146 640 555148 649
rect 555792 672 555844 678
rect 555200 640 555202 649
rect 555496 620 555792 626
rect 556896 672 556948 678
rect 555496 614 555844 620
rect 556158 640 556214 649
rect 555496 598 555832 614
rect 555146 575 555202 584
rect 556600 620 556896 626
rect 560850 640 560906 649
rect 556600 614 556948 620
rect 556600 598 556936 614
rect 557184 598 557396 626
rect 556158 575 556214 584
rect 554976 480 555004 575
rect 556172 480 556200 575
rect 552400 202 552428 462
rect 552388 196 552440 202
rect 552388 138 552440 144
rect 552634 -960 552746 480
rect 553308 264 553360 270
rect 553196 212 553308 218
rect 553196 206 553360 212
rect 553196 190 553348 206
rect 553738 -960 553850 480
rect 554300 202 554636 218
rect 554300 196 554648 202
rect 554300 190 554596 196
rect 554596 138 554648 144
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557184 66 557212 598
rect 557368 480 557396 598
rect 558380 598 558592 626
rect 558000 536 558052 542
rect 557704 484 558000 490
rect 558380 513 558408 598
rect 557172 60 557224 66
rect 557172 2 557224 8
rect 557326 -960 557438 480
rect 557704 478 558052 484
rect 558366 504 558422 513
rect 557704 462 558040 478
rect 558564 480 558592 598
rect 559576 598 559788 626
rect 558736 536 558788 542
rect 559576 513 559604 598
rect 559562 504 559618 513
rect 558788 484 558900 490
rect 558366 439 558422 448
rect 558522 -960 558634 480
rect 558736 478 558900 484
rect 558748 462 558900 478
rect 559760 480 559788 598
rect 560850 575 560906 584
rect 561784 598 562088 626
rect 560208 536 560260 542
rect 560004 484 560208 490
rect 559562 439 559618 448
rect 559718 -960 559830 480
rect 560004 478 560260 484
rect 560864 480 560892 575
rect 560004 462 560248 478
rect 560822 -960 560934 480
rect 561784 338 561812 598
rect 562060 480 562088 598
rect 563072 598 563284 626
rect 561772 332 561824 338
rect 561772 274 561824 280
rect 561108 66 561444 82
rect 561108 60 561456 66
rect 561108 54 561404 60
rect 561404 2 561456 8
rect 562018 -960 562130 480
rect 562304 474 562640 490
rect 562304 468 562652 474
rect 562304 462 562600 468
rect 562600 410 562652 416
rect 563072 406 563100 598
rect 563256 480 563284 598
rect 564452 598 564664 626
rect 564452 480 564480 598
rect 563060 400 563112 406
rect 563060 342 563112 348
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 564636 134 564664 598
rect 565464 598 565676 626
rect 565832 610 565860 750
rect 565464 338 565492 598
rect 565648 480 565676 598
rect 565820 604 565872 610
rect 565820 546 565872 552
rect 566844 480 566872 1158
rect 568028 808 568080 814
rect 568028 750 568080 756
rect 568040 480 568068 750
rect 569144 480 569172 1362
rect 569880 1018 569908 3062
rect 573916 2984 573968 2990
rect 573916 2926 573968 2932
rect 569868 1012 569920 1018
rect 569868 954 569920 960
rect 570328 740 570380 746
rect 570328 682 570380 688
rect 570340 480 570368 682
rect 571352 598 571564 626
rect 565452 332 565504 338
rect 565452 274 565504 280
rect 564624 128 564676 134
rect 564624 70 564676 76
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571352 354 571380 598
rect 571536 480 571564 598
rect 572732 598 572944 626
rect 572732 480 572760 598
rect 571168 326 571380 354
rect 571168 270 571196 326
rect 571156 264 571208 270
rect 571156 206 571208 212
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 572916 202 572944 598
rect 573928 480 573956 2926
rect 575480 2916 575532 2922
rect 575480 2858 575532 2864
rect 575492 950 575520 2858
rect 576308 2848 576360 2854
rect 576308 2790 576360 2796
rect 575480 944 575532 950
rect 575480 886 575532 892
rect 575112 672 575164 678
rect 575112 614 575164 620
rect 575124 480 575152 614
rect 576320 480 576348 2790
rect 577424 480 577452 3062
rect 583392 3052 583444 3058
rect 583392 2994 583444 3000
rect 582196 2916 582248 2922
rect 582196 2858 582248 2864
rect 578608 604 578660 610
rect 578608 546 578660 552
rect 580828 598 581040 626
rect 578620 480 578648 546
rect 572904 196 572956 202
rect 572904 138 572956 144
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580828 218 580856 598
rect 581012 480 581040 598
rect 582208 480 582236 2858
rect 583404 480 583432 2994
rect 580736 190 580856 218
rect 580736 66 580764 190
rect 580724 60 580776 66
rect 580724 2 580776 8
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 110 701664 166 701720
rect 386 701936 442 701992
rect 1582 684256 1638 684312
rect 1030 658144 1086 658200
rect 1674 632032 1730 632088
rect 938 606056 994 606112
rect 1766 579944 1822 580000
rect 846 553832 902 553888
rect 2226 701800 2282 701856
rect 2042 701392 2098 701448
rect 1950 697992 2006 698048
rect 1858 527856 1914 527912
rect 754 501744 810 501800
rect 1950 475632 2006 475688
rect 662 449520 718 449576
rect 570 293120 626 293176
rect 570 267144 626 267200
rect 570 254088 626 254144
rect 570 162832 626 162888
rect 202 111152 258 111208
rect 110 85176 166 85232
rect 18 71848 74 71904
rect 2134 697584 2190 697640
rect 2134 214920 2190 214976
rect 2318 697856 2374 697912
rect 2686 698128 2742 698184
rect 3054 671200 3110 671256
rect 2962 619112 3018 619168
rect 3238 700440 3294 700496
rect 3146 566888 3202 566944
rect 3054 462576 3110 462632
rect 2686 423544 2742 423600
rect 2594 397432 2650 397488
rect 2502 371320 2558 371376
rect 2410 358400 2466 358456
rect 2318 319232 2374 319288
rect 3238 410488 3294 410544
rect 3606 699896 3662 699952
rect 3514 698400 3570 698456
rect 3330 345344 3386 345400
rect 3146 306176 3202 306232
rect 2226 188808 2282 188864
rect 2042 58520 2098 58576
rect 3882 700168 3938 700224
rect 4066 514800 4122 514856
rect 4434 701256 4490 701312
rect 16302 702344 16358 702400
rect 31206 701528 31262 701584
rect 60646 700032 60702 700088
rect 90178 700304 90234 700360
rect 26146 699760 26202 699816
rect 163870 700576 163926 700632
rect 207018 702072 207074 702128
rect 252282 701120 252338 701176
rect 286690 701120 286746 701176
rect 298006 701120 298062 701176
rect 443274 700440 443330 700496
rect 487434 701936 487490 701992
rect 497278 701800 497334 701856
rect 502476 700168 502532 700224
rect 516966 702072 517022 702128
rect 526718 701664 526774 701720
rect 546498 701392 546554 701448
rect 531686 699896 531742 699952
rect 551282 701256 551338 701312
rect 561126 702208 561182 702264
rect 386234 699508 386290 699544
rect 386234 699488 386236 699508
rect 386236 699488 386288 699508
rect 386288 699488 386290 699508
rect 11610 699352 11666 699408
rect 41050 699352 41106 699408
rect 46018 699352 46074 699408
rect 50894 699352 50950 699408
rect 55770 699352 55826 699408
rect 95146 699352 95202 699408
rect 124586 699352 124642 699408
rect 418710 699352 418766 699408
rect 433430 699352 433486 699408
rect 462870 699352 462926 699408
rect 492586 699352 492642 699408
rect 541530 699352 541586 699408
rect 3974 241032 4030 241088
rect 3882 201864 3938 201920
rect 3790 149776 3846 149832
rect 3698 136720 3754 136776
rect 3606 97552 3662 97608
rect 3514 45464 3570 45520
rect 4066 32408 4122 32464
rect 3422 19352 3478 19408
rect 2962 6432 3018 6488
rect 565082 699760 565138 699816
rect 565174 698808 565230 698864
rect 565266 697720 565322 697776
rect 566646 698536 566702 698592
rect 566462 698264 566518 698320
rect 569222 701528 569278 701584
rect 570694 700032 570750 700088
rect 569314 698944 569370 699000
rect 570602 698672 570658 698728
rect 570786 697992 570842 698048
rect 573362 700304 573418 700360
rect 576306 700576 576362 700632
rect 577502 702344 577558 702400
rect 580262 699080 580318 699136
rect 580170 697176 580226 697232
rect 579066 683848 579122 683904
rect 579618 670656 579674 670712
rect 580170 644000 580226 644056
rect 580170 630808 580226 630864
rect 580170 617480 580226 617536
rect 580170 590960 580226 591016
rect 578974 577632 579030 577688
rect 580170 564340 580172 564360
rect 580172 564340 580224 564360
rect 580224 564340 580226 564360
rect 580170 564304 580226 564340
rect 580170 537784 580226 537840
rect 580170 511264 580226 511320
rect 578882 484608 578938 484664
rect 579802 471416 579858 471472
rect 579710 431568 579766 431624
rect 580170 418240 580226 418296
rect 580170 404912 580226 404968
rect 579618 378392 579674 378448
rect 580170 365064 580226 365120
rect 580170 351872 580226 351928
rect 579710 312024 579766 312080
rect 579802 298696 579858 298752
rect 580170 272176 580226 272232
rect 580170 245556 580172 245576
rect 580172 245556 580224 245576
rect 580224 245556 580226 245576
rect 580170 245520 580226 245556
rect 580170 232328 580226 232384
rect 580170 219000 580226 219056
rect 579894 205672 579950 205728
rect 580170 192480 580226 192536
rect 580170 165824 580226 165880
rect 579802 152632 579858 152688
rect 580170 139340 580172 139360
rect 580172 139340 580224 139360
rect 580224 139340 580226 139360
rect 580170 139304 580226 139340
rect 580170 125976 580226 126032
rect 580170 112784 580226 112840
rect 580170 99456 580226 99512
rect 580170 86128 580226 86184
rect 579986 72936 580042 72992
rect 580170 59608 580226 59664
rect 580170 46280 580226 46336
rect 580170 33108 580226 33144
rect 580170 33088 580172 33108
rect 580172 33088 580224 33108
rect 580224 33088 580226 33108
rect 579710 19760 579766 19816
rect 580722 524456 580778 524512
rect 580630 458088 580686 458144
rect 580538 325216 580594 325272
rect 580446 258848 580502 258904
rect 580354 179152 580410 179208
rect 580262 6568 580318 6624
rect 8758 584 8814 640
rect 9954 584 10010 640
rect 13266 584 13322 640
rect 12622 448 12678 504
rect 20626 584 20682 640
rect 23478 584 23534 640
rect 26514 584 26570 640
rect 28722 604 28778 640
rect 28722 584 28724 604
rect 28724 584 28776 604
rect 28776 584 28778 604
rect 27894 448 27950 504
rect 30286 584 30342 640
rect 34794 584 34850 640
rect 35990 584 36046 640
rect 37370 448 37426 504
rect 38474 584 38530 640
rect 52550 584 52606 640
rect 53562 448 53618 504
rect 54206 584 54262 640
rect 56046 584 56102 640
rect 55310 448 55366 504
rect 57610 584 57666 640
rect 58438 584 58494 640
rect 57426 448 57482 504
rect 59818 584 59874 640
rect 60830 584 60886 640
rect 58806 448 58862 504
rect 59450 448 59506 504
rect 62118 584 62174 640
rect 61106 448 61162 504
rect 142066 584 142122 640
rect 143446 584 143502 640
rect 144734 584 144790 640
rect 145746 584 145802 640
rect 143722 448 143778 504
rect 147126 584 147182 640
rect 148966 584 149022 640
rect 147770 448 147826 504
rect 149334 448 149390 504
rect 150622 584 150678 640
rect 151818 584 151874 640
rect 150254 448 150310 504
rect 164790 584 164846 640
rect 167366 584 167422 640
rect 169482 584 169538 640
rect 168194 312 168250 368
rect 171966 584 172022 640
rect 172978 584 173034 640
rect 170954 312 171010 368
rect 171690 312 171746 368
rect 173898 448 173954 504
rect 175462 584 175518 640
rect 176382 584 176438 640
rect 173990 312 174046 368
rect 175186 312 175242 368
rect 176842 448 176898 504
rect 177486 448 177542 504
rect 179050 584 179106 640
rect 180246 584 180302 640
rect 177670 312 177726 368
rect 178682 312 178738 368
rect 182086 584 182142 640
rect 184938 584 184994 640
rect 181258 312 181314 368
rect 186594 448 186650 504
rect 192298 584 192354 640
rect 189906 448 189962 504
rect 194046 448 194102 504
rect 195610 584 195666 640
rect 197910 584 197966 640
rect 200026 584 200082 640
rect 196622 312 196678 368
rect 197726 40 197782 96
rect 198922 448 198978 504
rect 200118 312 200174 368
rect 201314 448 201370 504
rect 203890 584 203946 640
rect 204166 604 204222 640
rect 204166 584 204168 604
rect 204168 584 204220 604
rect 204220 584 204222 604
rect 202510 312 202566 368
rect 202418 176 202474 232
rect 201682 40 201738 96
rect 204902 448 204958 504
rect 207386 584 207442 640
rect 208214 584 208270 640
rect 208398 584 208454 640
rect 204810 312 204866 368
rect 206006 176 206062 232
rect 206926 448 206982 504
rect 209318 584 209374 640
rect 208766 312 208822 368
rect 210790 448 210846 504
rect 213366 584 213422 640
rect 216126 584 216182 640
rect 220726 584 220782 640
rect 221830 584 221886 640
rect 223578 448 223634 504
rect 226338 584 226394 640
rect 228730 584 228786 640
rect 230938 584 230994 640
rect 235814 584 235870 640
rect 237746 584 237802 640
rect 242898 584 242954 640
rect 242254 448 242310 504
rect 249706 584 249762 640
rect 247314 448 247370 504
rect 255870 584 255926 640
rect 267278 584 267334 640
rect 273626 584 273682 640
rect 275190 584 275246 640
rect 282090 584 282146 640
rect 285678 584 285734 640
rect 285218 448 285274 504
rect 287794 584 287850 640
rect 286414 312 286470 368
rect 292578 584 292634 640
rect 293406 312 293462 368
rect 294602 584 294658 640
rect 296074 584 296130 640
rect 305826 584 305882 640
rect 313830 584 313886 640
rect 315026 584 315082 640
rect 307022 448 307078 504
rect 316590 584 316646 640
rect 317326 584 317382 640
rect 328458 584 328514 640
rect 334254 448 334310 504
rect 337474 584 337530 640
rect 338302 312 338358 368
rect 343362 584 343418 640
rect 345018 584 345074 640
rect 346950 584 347006 640
rect 347870 448 347926 504
rect 349066 604 349122 640
rect 349066 584 349068 604
rect 349068 584 349120 604
rect 349120 584 349122 604
rect 350446 584 350502 640
rect 350630 584 350686 640
rect 350170 448 350226 504
rect 352838 584 352894 640
rect 359922 584 359978 640
rect 363786 584 363842 640
rect 361486 312 361542 368
rect 362682 448 362738 504
rect 374090 584 374146 640
rect 374274 620 374276 640
rect 374276 620 374328 640
rect 374328 620 374330 640
rect 374274 584 374330 620
rect 372710 448 372766 504
rect 371974 312 372030 368
rect 377678 584 377734 640
rect 377954 620 377956 640
rect 377956 620 378008 640
rect 378008 620 378010 640
rect 377954 584 378010 620
rect 375654 468 375710 504
rect 375654 448 375656 468
rect 375656 448 375708 468
rect 375708 448 375710 468
rect 378690 448 378746 504
rect 379978 584 380034 640
rect 380162 604 380218 640
rect 380162 584 380164 604
rect 380164 584 380216 604
rect 380216 584 380218 604
rect 380898 484 380900 504
rect 380900 484 380952 504
rect 380952 484 380954 504
rect 380898 448 380954 484
rect 382370 584 382426 640
rect 384762 584 384818 640
rect 385406 584 385462 640
rect 392398 448 392454 504
rect 396538 584 396594 640
rect 392214 312 392270 368
rect 401414 584 401470 640
rect 400310 312 400366 368
rect 405830 584 405886 640
rect 405094 312 405150 368
rect 409602 584 409658 640
rect 412638 584 412694 640
rect 408222 312 408278 368
rect 421746 584 421802 640
rect 424506 484 424508 504
rect 424508 484 424560 504
rect 424560 484 424562 504
rect 424506 448 424562 484
rect 427266 584 427322 640
rect 429014 584 429070 640
rect 429658 584 429714 640
rect 446678 312 446734 368
rect 456062 584 456118 640
rect 451922 332 451978 368
rect 451922 312 451924 332
rect 451924 312 451976 332
rect 451976 312 451978 332
rect 460478 584 460534 640
rect 462134 584 462190 640
rect 463974 584 464030 640
rect 466090 584 466146 640
rect 467470 584 467526 640
rect 468298 448 468354 504
rect 470598 584 470654 640
rect 476578 448 476634 504
rect 477406 584 477462 640
rect 483202 584 483258 640
rect 488814 584 488870 640
rect 491298 620 491300 640
rect 491300 620 491352 640
rect 491352 620 491354 640
rect 483662 196 483718 232
rect 483662 176 483664 196
rect 483664 176 483716 196
rect 483716 176 483718 196
rect 491298 584 491354 620
rect 493322 448 493378 504
rect 492678 312 492734 368
rect 492494 176 492550 232
rect 495898 584 495954 640
rect 497094 550 497150 606
rect 498014 584 498070 640
rect 493782 312 493838 368
rect 500590 584 500646 640
rect 508594 332 508650 368
rect 509698 448 509754 504
rect 508594 312 508596 332
rect 508596 312 508648 332
rect 508648 312 508650 332
rect 514666 584 514722 640
rect 518346 584 518402 640
rect 517334 312 517390 368
rect 531318 584 531374 640
rect 527178 312 527234 368
rect 530766 40 530822 96
rect 534170 176 534226 232
rect 540518 448 540574 504
rect 541714 584 541770 640
rect 543094 584 543150 640
rect 543462 584 543518 640
rect 544566 312 544622 368
rect 548062 40 548118 96
rect 551282 176 551338 232
rect 554962 584 555018 640
rect 555146 620 555148 640
rect 555148 620 555200 640
rect 555200 620 555202 640
rect 555146 584 555202 620
rect 556158 584 556214 640
rect 558366 448 558422 504
rect 559562 448 559618 504
rect 560850 584 560906 640
<< metal3 >>
rect 16297 702402 16363 702405
rect 577497 702402 577563 702405
rect 16297 702400 577563 702402
rect 16297 702344 16302 702400
rect 16358 702344 577502 702400
rect 577558 702344 577563 702400
rect 16297 702342 577563 702344
rect 16297 702339 16363 702342
rect 577497 702339 577563 702342
rect 386270 702204 386276 702268
rect 386340 702266 386346 702268
rect 561121 702266 561187 702269
rect 386340 702264 561187 702266
rect 386340 702208 561126 702264
rect 561182 702208 561187 702264
rect 386340 702206 561187 702208
rect 386340 702204 386346 702206
rect 561121 702203 561187 702206
rect 207013 702130 207079 702133
rect 516961 702130 517027 702133
rect 207013 702128 517027 702130
rect 207013 702072 207018 702128
rect 207074 702072 516966 702128
rect 517022 702072 517027 702128
rect 207013 702070 517027 702072
rect 207013 702067 207079 702070
rect 516961 702067 517027 702070
rect 381 701994 447 701997
rect 487429 701994 487495 701997
rect 381 701992 487495 701994
rect 381 701936 386 701992
rect 442 701936 487434 701992
rect 487490 701936 487495 701992
rect 381 701934 487495 701936
rect 381 701931 447 701934
rect 487429 701931 487495 701934
rect 2221 701858 2287 701861
rect 497273 701858 497339 701861
rect 2221 701856 497339 701858
rect 2221 701800 2226 701856
rect 2282 701800 497278 701856
rect 497334 701800 497339 701856
rect 2221 701798 497339 701800
rect 2221 701795 2287 701798
rect 497273 701795 497339 701798
rect 105 701722 171 701725
rect 526713 701722 526779 701725
rect 105 701720 526779 701722
rect 105 701664 110 701720
rect 166 701664 526718 701720
rect 526774 701664 526779 701720
rect 105 701662 526779 701664
rect 105 701659 171 701662
rect 526713 701659 526779 701662
rect 31201 701586 31267 701589
rect 569217 701586 569283 701589
rect 31201 701584 569283 701586
rect 31201 701528 31206 701584
rect 31262 701528 569222 701584
rect 569278 701528 569283 701584
rect 31201 701526 569283 701528
rect 31201 701523 31267 701526
rect 569217 701523 569283 701526
rect 2037 701450 2103 701453
rect 546493 701450 546559 701453
rect 2037 701448 546559 701450
rect 2037 701392 2042 701448
rect 2098 701392 546498 701448
rect 546554 701392 546559 701448
rect 2037 701390 546559 701392
rect 2037 701387 2103 701390
rect 546493 701387 546559 701390
rect 4429 701314 4495 701317
rect 551277 701314 551343 701317
rect 4429 701312 551343 701314
rect 4429 701256 4434 701312
rect 4490 701256 551282 701312
rect 551338 701256 551343 701312
rect 4429 701254 551343 701256
rect 4429 701251 4495 701254
rect 551277 701251 551343 701254
rect 252277 701178 252343 701181
rect 259126 701178 259132 701180
rect 252277 701176 259132 701178
rect 252277 701120 252282 701176
rect 252338 701120 259132 701176
rect 252277 701118 259132 701120
rect 252277 701115 252343 701118
rect 259126 701116 259132 701118
rect 259196 701116 259202 701180
rect 286685 701178 286751 701181
rect 298001 701178 298067 701181
rect 286685 701176 298067 701178
rect 286685 701120 286690 701176
rect 286746 701120 298006 701176
rect 298062 701120 298067 701176
rect 286685 701118 298067 701120
rect 286685 701115 286751 701118
rect 298001 701115 298067 701118
rect 163865 700634 163931 700637
rect 576301 700634 576367 700637
rect 163865 700632 576367 700634
rect 163865 700576 163870 700632
rect 163926 700576 576306 700632
rect 576362 700576 576367 700632
rect 163865 700574 576367 700576
rect 163865 700571 163931 700574
rect 576301 700571 576367 700574
rect 3233 700498 3299 700501
rect 443269 700498 443335 700501
rect 3233 700496 443335 700498
rect 3233 700440 3238 700496
rect 3294 700440 443274 700496
rect 443330 700440 443335 700496
rect 3233 700438 443335 700440
rect 3233 700435 3299 700438
rect 443269 700435 443335 700438
rect 90173 700362 90239 700365
rect 573357 700362 573423 700365
rect 90173 700360 573423 700362
rect 90173 700304 90178 700360
rect 90234 700304 573362 700360
rect 573418 700304 573423 700360
rect 90173 700302 573423 700304
rect 90173 700299 90239 700302
rect 573357 700299 573423 700302
rect 3877 700226 3943 700229
rect 502471 700226 502537 700229
rect 3877 700224 502537 700226
rect 3877 700168 3882 700224
rect 3938 700168 502476 700224
rect 502532 700168 502537 700224
rect 3877 700166 502537 700168
rect 3877 700163 3943 700166
rect 502471 700163 502537 700166
rect 60641 700090 60707 700093
rect 570689 700090 570755 700093
rect 60641 700088 570755 700090
rect 60641 700032 60646 700088
rect 60702 700032 570694 700088
rect 570750 700032 570755 700088
rect 60641 700030 570755 700032
rect 60641 700027 60707 700030
rect 570689 700027 570755 700030
rect 3601 699954 3667 699957
rect 531681 699954 531747 699957
rect 3601 699952 531747 699954
rect 3601 699896 3606 699952
rect 3662 699896 531686 699952
rect 531742 699896 531747 699952
rect 3601 699894 531747 699896
rect 3601 699891 3667 699894
rect 531681 699891 531747 699894
rect 26141 699818 26207 699821
rect 565077 699818 565143 699821
rect 26141 699816 565143 699818
rect 26141 699760 26146 699816
rect 26202 699760 565082 699816
rect 565138 699760 565143 699816
rect 26141 699758 565143 699760
rect 26141 699755 26207 699758
rect 565077 699755 565143 699758
rect 386229 699548 386295 699549
rect 386229 699546 386276 699548
rect 386184 699544 386276 699546
rect 386184 699488 386234 699544
rect 386184 699486 386276 699488
rect 386229 699484 386276 699486
rect 386340 699484 386346 699548
rect 386229 699483 386295 699484
rect 11605 699410 11671 699413
rect 13854 699410 13860 699412
rect 11605 699408 13860 699410
rect 11605 699352 11610 699408
rect 11666 699352 13860 699408
rect 11605 699350 13860 699352
rect 11605 699347 11671 699350
rect 13854 699348 13860 699350
rect 13924 699348 13930 699412
rect 41045 699410 41111 699413
rect 46013 699410 46079 699413
rect 50889 699410 50955 699413
rect 55765 699410 55831 699413
rect 95141 699412 95207 699413
rect 41045 699408 45570 699410
rect 41045 699352 41050 699408
rect 41106 699352 45570 699408
rect 41045 699350 45570 699352
rect 41045 699347 41111 699350
rect 45510 698594 45570 699350
rect 46013 699408 50538 699410
rect 46013 699352 46018 699408
rect 46074 699352 50538 699408
rect 46013 699350 50538 699352
rect 46013 699347 46079 699350
rect 50478 698730 50538 699350
rect 50889 699408 55230 699410
rect 50889 699352 50894 699408
rect 50950 699352 55230 699408
rect 50889 699350 55230 699352
rect 50889 699347 50955 699350
rect 55170 698866 55230 699350
rect 55765 699408 64890 699410
rect 55765 699352 55770 699408
rect 55826 699352 64890 699408
rect 55765 699350 64890 699352
rect 55765 699347 55831 699350
rect 64830 699002 64890 699350
rect 95141 699408 95188 699412
rect 95252 699410 95258 699412
rect 124581 699410 124647 699413
rect 418705 699412 418771 699413
rect 433425 699412 433491 699413
rect 462865 699412 462931 699413
rect 418654 699410 418660 699412
rect 95141 699352 95146 699408
rect 95141 699348 95188 699352
rect 95252 699350 95298 699410
rect 124581 699408 132510 699410
rect 124581 699352 124586 699408
rect 124642 699352 132510 699408
rect 124581 699350 132510 699352
rect 95252 699348 95258 699350
rect 95141 699347 95207 699348
rect 124581 699347 124647 699350
rect 132450 699138 132510 699350
rect 251130 699350 260850 699410
rect 418614 699350 418660 699410
rect 418724 699408 418771 699412
rect 433374 699410 433380 699412
rect 418766 699352 418771 699408
rect 251130 699138 251190 699350
rect 260790 699274 260850 699350
rect 418654 699348 418660 699350
rect 418724 699348 418771 699352
rect 433334 699350 433380 699410
rect 433444 699408 433491 699412
rect 462814 699410 462820 699412
rect 433486 699352 433491 699408
rect 433374 699348 433380 699350
rect 433444 699348 433491 699352
rect 462774 699350 462820 699410
rect 462884 699408 462931 699412
rect 462926 699352 462931 699408
rect 462814 699348 462820 699350
rect 462884 699348 462931 699352
rect 418705 699347 418771 699348
rect 433425 699347 433491 699348
rect 462865 699347 462931 699348
rect 492581 699412 492647 699413
rect 492581 699408 492628 699412
rect 492692 699410 492698 699412
rect 492581 699352 492586 699408
rect 492581 699348 492628 699352
rect 492692 699350 492738 699410
rect 492692 699348 492698 699350
rect 539910 699348 539916 699412
rect 539980 699410 539986 699412
rect 541525 699410 541591 699413
rect 539980 699408 541591 699410
rect 539980 699352 541530 699408
rect 541586 699352 541591 699408
rect 539980 699350 541591 699352
rect 539980 699348 539986 699350
rect 492581 699347 492647 699348
rect 541525 699347 541591 699350
rect 418838 699274 418844 699276
rect 260790 699214 418844 699274
rect 418838 699212 418844 699214
rect 418908 699212 418914 699276
rect 132450 699078 251190 699138
rect 259126 699076 259132 699140
rect 259196 699138 259202 699140
rect 580257 699138 580323 699141
rect 259196 699136 580323 699138
rect 259196 699080 580262 699136
rect 580318 699080 580323 699136
rect 259196 699078 580323 699080
rect 259196 699076 259202 699078
rect 580257 699075 580323 699078
rect 569309 699002 569375 699005
rect 64830 699000 569375 699002
rect 64830 698944 569314 699000
rect 569370 698944 569375 699000
rect 64830 698942 569375 698944
rect 569309 698939 569375 698942
rect 565169 698866 565235 698869
rect 55170 698864 565235 698866
rect 55170 698808 565174 698864
rect 565230 698808 565235 698864
rect 55170 698806 565235 698808
rect 565169 698803 565235 698806
rect 570597 698730 570663 698733
rect 50478 698728 570663 698730
rect 50478 698672 570602 698728
rect 570658 698672 570663 698728
rect 50478 698670 570663 698672
rect 570597 698667 570663 698670
rect 566641 698594 566707 698597
rect 45510 698592 566707 698594
rect 45510 698536 566646 698592
rect 566702 698536 566707 698592
rect 45510 698534 566707 698536
rect 566641 698531 566707 698534
rect 3509 698458 3575 698461
rect 539910 698458 539916 698460
rect 3509 698456 539916 698458
rect 3509 698400 3514 698456
rect 3570 698400 539916 698456
rect 3509 698398 539916 698400
rect 3509 698395 3575 698398
rect 539910 698396 539916 698398
rect 539980 698396 539986 698460
rect 13854 698260 13860 698324
rect 13924 698322 13930 698324
rect 566457 698322 566523 698325
rect 13924 698320 566523 698322
rect 13924 698264 566462 698320
rect 566518 698264 566523 698320
rect 13924 698262 566523 698264
rect 13924 698260 13930 698262
rect 566457 698259 566523 698262
rect 2681 698186 2747 698189
rect 433374 698186 433380 698188
rect 2681 698184 433380 698186
rect 2681 698128 2686 698184
rect 2742 698128 433380 698184
rect 2681 698126 433380 698128
rect 2681 698123 2747 698126
rect 433374 698124 433380 698126
rect 433444 698124 433450 698188
rect 1945 698050 2011 698053
rect 418654 698050 418660 698052
rect 1945 698048 418660 698050
rect 1945 697992 1950 698048
rect 2006 697992 418660 698048
rect 1945 697990 418660 697992
rect 1945 697987 2011 697990
rect 418654 697988 418660 697990
rect 418724 697988 418730 698052
rect 418838 697988 418844 698052
rect 418908 698050 418914 698052
rect 570781 698050 570847 698053
rect 418908 698048 570847 698050
rect 418908 697992 570786 698048
rect 570842 697992 570847 698048
rect 418908 697990 570847 697992
rect 418908 697988 418914 697990
rect 570781 697987 570847 697990
rect 2313 697914 2379 697917
rect 462814 697914 462820 697916
rect 2313 697912 462820 697914
rect 2313 697856 2318 697912
rect 2374 697856 462820 697912
rect 2313 697854 462820 697856
rect 2313 697851 2379 697854
rect 462814 697852 462820 697854
rect 462884 697852 462890 697916
rect 95182 697716 95188 697780
rect 95252 697778 95258 697780
rect 565261 697778 565327 697781
rect 95252 697776 565327 697778
rect 95252 697720 565266 697776
rect 565322 697720 565327 697776
rect 95252 697718 565327 697720
rect 95252 697716 95258 697718
rect 565261 697715 565327 697718
rect 2129 697642 2195 697645
rect 492622 697642 492628 697644
rect 2129 697640 492628 697642
rect 2129 697584 2134 697640
rect 2190 697584 492628 697640
rect 2129 697582 492628 697584
rect 2129 697579 2195 697582
rect 492622 697580 492628 697582
rect 492692 697580 492698 697644
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 1577 684314 1643 684317
rect -960 684312 1643 684314
rect -960 684256 1582 684312
rect 1638 684256 1643 684312
rect -960 684254 1643 684256
rect -960 684164 480 684254
rect 1577 684251 1643 684254
rect 579061 683906 579127 683909
rect 583520 683906 584960 683996
rect 579061 683904 584960 683906
rect 579061 683848 579066 683904
rect 579122 683848 584960 683904
rect 579061 683846 584960 683848
rect 579061 683843 579127 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3049 671258 3115 671261
rect -960 671256 3115 671258
rect -960 671200 3054 671256
rect 3110 671200 3115 671256
rect -960 671198 3115 671200
rect -960 671108 480 671198
rect 3049 671195 3115 671198
rect 579613 670714 579679 670717
rect 583520 670714 584960 670804
rect 579613 670712 584960 670714
rect 579613 670656 579618 670712
rect 579674 670656 584960 670712
rect 579613 670654 584960 670656
rect 579613 670651 579679 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 1025 658202 1091 658205
rect -960 658200 1091 658202
rect -960 658144 1030 658200
rect 1086 658144 1091 658200
rect -960 658142 1091 658144
rect -960 658052 480 658142
rect 1025 658139 1091 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 1669 632090 1735 632093
rect -960 632088 1735 632090
rect -960 632032 1674 632088
rect 1730 632032 1735 632088
rect -960 632030 1735 632032
rect -960 631940 480 632030
rect 1669 632027 1735 632030
rect 580165 630866 580231 630869
rect 583520 630866 584960 630956
rect 580165 630864 584960 630866
rect 580165 630808 580170 630864
rect 580226 630808 584960 630864
rect 580165 630806 584960 630808
rect 580165 630803 580231 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 2957 619170 3023 619173
rect -960 619168 3023 619170
rect -960 619112 2962 619168
rect 3018 619112 3023 619168
rect -960 619110 3023 619112
rect -960 619020 480 619110
rect 2957 619107 3023 619110
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 933 606114 999 606117
rect -960 606112 999 606114
rect -960 606056 938 606112
rect 994 606056 999 606112
rect -960 606054 999 606056
rect -960 605964 480 606054
rect 933 606051 999 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 580165 591018 580231 591021
rect 583520 591018 584960 591108
rect 580165 591016 584960 591018
rect 580165 590960 580170 591016
rect 580226 590960 584960 591016
rect 580165 590958 584960 590960
rect 580165 590955 580231 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 1761 580002 1827 580005
rect -960 580000 1827 580002
rect -960 579944 1766 580000
rect 1822 579944 1827 580000
rect -960 579942 1827 579944
rect -960 579852 480 579942
rect 1761 579939 1827 579942
rect 578969 577690 579035 577693
rect 583520 577690 584960 577780
rect 578969 577688 584960 577690
rect 578969 577632 578974 577688
rect 579030 577632 584960 577688
rect 578969 577630 584960 577632
rect 578969 577627 579035 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3141 566946 3207 566949
rect -960 566944 3207 566946
rect -960 566888 3146 566944
rect 3202 566888 3207 566944
rect -960 566886 3207 566888
rect -960 566796 480 566886
rect 3141 566883 3207 566886
rect 580165 564362 580231 564365
rect 583520 564362 584960 564452
rect 580165 564360 584960 564362
rect 580165 564304 580170 564360
rect 580226 564304 584960 564360
rect 580165 564302 584960 564304
rect 580165 564299 580231 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 841 553890 907 553893
rect -960 553888 907 553890
rect -960 553832 846 553888
rect 902 553832 907 553888
rect -960 553830 907 553832
rect -960 553740 480 553830
rect 841 553827 907 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 580165 537842 580231 537845
rect 583520 537842 584960 537932
rect 580165 537840 584960 537842
rect 580165 537784 580170 537840
rect 580226 537784 584960 537840
rect 580165 537782 584960 537784
rect 580165 537779 580231 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 1853 527914 1919 527917
rect -960 527912 1919 527914
rect -960 527856 1858 527912
rect 1914 527856 1919 527912
rect -960 527854 1919 527856
rect -960 527764 480 527854
rect 1853 527851 1919 527854
rect 580717 524514 580783 524517
rect 583520 524514 584960 524604
rect 580717 524512 584960 524514
rect 580717 524456 580722 524512
rect 580778 524456 584960 524512
rect 580717 524454 584960 524456
rect 580717 524451 580783 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 4061 514858 4127 514861
rect -960 514856 4127 514858
rect -960 514800 4066 514856
rect 4122 514800 4127 514856
rect -960 514798 4127 514800
rect -960 514708 480 514798
rect 4061 514795 4127 514798
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 749 501802 815 501805
rect -960 501800 815 501802
rect -960 501744 754 501800
rect 810 501744 815 501800
rect -960 501742 815 501744
rect -960 501652 480 501742
rect 749 501739 815 501742
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 578877 484666 578943 484669
rect 583520 484666 584960 484756
rect 578877 484664 584960 484666
rect 578877 484608 578882 484664
rect 578938 484608 584960 484664
rect 578877 484606 584960 484608
rect 578877 484603 578943 484606
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect 1945 475690 2011 475693
rect -960 475688 2011 475690
rect -960 475632 1950 475688
rect 2006 475632 2011 475688
rect -960 475630 2011 475632
rect -960 475540 480 475630
rect 1945 475627 2011 475630
rect 579797 471474 579863 471477
rect 583520 471474 584960 471564
rect 579797 471472 584960 471474
rect 579797 471416 579802 471472
rect 579858 471416 584960 471472
rect 579797 471414 584960 471416
rect 579797 471411 579863 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 3049 462634 3115 462637
rect -960 462632 3115 462634
rect -960 462576 3054 462632
rect 3110 462576 3115 462632
rect -960 462574 3115 462576
rect -960 462484 480 462574
rect 3049 462571 3115 462574
rect 580625 458146 580691 458149
rect 583520 458146 584960 458236
rect 580625 458144 584960 458146
rect 580625 458088 580630 458144
rect 580686 458088 584960 458144
rect 580625 458086 584960 458088
rect 580625 458083 580691 458086
rect 583520 457996 584960 458086
rect -960 449578 480 449668
rect 657 449578 723 449581
rect -960 449576 723 449578
rect -960 449520 662 449576
rect 718 449520 723 449576
rect -960 449518 723 449520
rect -960 449428 480 449518
rect 657 449515 723 449518
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 579705 431626 579771 431629
rect 583520 431626 584960 431716
rect 579705 431624 584960 431626
rect 579705 431568 579710 431624
rect 579766 431568 584960 431624
rect 579705 431566 584960 431568
rect 579705 431563 579771 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 2681 423602 2747 423605
rect -960 423600 2747 423602
rect -960 423544 2686 423600
rect 2742 423544 2747 423600
rect -960 423542 2747 423544
rect -960 423452 480 423542
rect 2681 423539 2747 423542
rect 580165 418298 580231 418301
rect 583520 418298 584960 418388
rect 580165 418296 584960 418298
rect 580165 418240 580170 418296
rect 580226 418240 584960 418296
rect 580165 418238 584960 418240
rect 580165 418235 580231 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 3233 410546 3299 410549
rect -960 410544 3299 410546
rect -960 410488 3238 410544
rect 3294 410488 3299 410544
rect -960 410486 3299 410488
rect -960 410396 480 410486
rect 3233 410483 3299 410486
rect 580165 404970 580231 404973
rect 583520 404970 584960 405060
rect 580165 404968 584960 404970
rect 580165 404912 580170 404968
rect 580226 404912 584960 404968
rect 580165 404910 584960 404912
rect 580165 404907 580231 404910
rect 583520 404820 584960 404910
rect -960 397490 480 397580
rect 2589 397490 2655 397493
rect -960 397488 2655 397490
rect -960 397432 2594 397488
rect 2650 397432 2655 397488
rect -960 397430 2655 397432
rect -960 397340 480 397430
rect 2589 397427 2655 397430
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 579613 378450 579679 378453
rect 583520 378450 584960 378540
rect 579613 378448 584960 378450
rect 579613 378392 579618 378448
rect 579674 378392 584960 378448
rect 579613 378390 584960 378392
rect 579613 378387 579679 378390
rect 583520 378300 584960 378390
rect -960 371378 480 371468
rect 2497 371378 2563 371381
rect -960 371376 2563 371378
rect -960 371320 2502 371376
rect 2558 371320 2563 371376
rect -960 371318 2563 371320
rect -960 371228 480 371318
rect 2497 371315 2563 371318
rect 580165 365122 580231 365125
rect 583520 365122 584960 365212
rect 580165 365120 584960 365122
rect 580165 365064 580170 365120
rect 580226 365064 584960 365120
rect 580165 365062 584960 365064
rect 580165 365059 580231 365062
rect 583520 364972 584960 365062
rect -960 358458 480 358548
rect 2405 358458 2471 358461
rect -960 358456 2471 358458
rect -960 358400 2410 358456
rect 2466 358400 2471 358456
rect -960 358398 2471 358400
rect -960 358308 480 358398
rect 2405 358395 2471 358398
rect 580165 351930 580231 351933
rect 583520 351930 584960 352020
rect 580165 351928 584960 351930
rect 580165 351872 580170 351928
rect 580226 351872 584960 351928
rect 580165 351870 584960 351872
rect 580165 351867 580231 351870
rect 583520 351780 584960 351870
rect -960 345402 480 345492
rect 3325 345402 3391 345405
rect -960 345400 3391 345402
rect -960 345344 3330 345400
rect 3386 345344 3391 345400
rect -960 345342 3391 345344
rect -960 345252 480 345342
rect 3325 345339 3391 345342
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 580533 325274 580599 325277
rect 583520 325274 584960 325364
rect 580533 325272 584960 325274
rect 580533 325216 580538 325272
rect 580594 325216 584960 325272
rect 580533 325214 584960 325216
rect 580533 325211 580599 325214
rect 583520 325124 584960 325214
rect -960 319290 480 319380
rect 2313 319290 2379 319293
rect -960 319288 2379 319290
rect -960 319232 2318 319288
rect 2374 319232 2379 319288
rect -960 319230 2379 319232
rect -960 319140 480 319230
rect 2313 319227 2379 319230
rect 579705 312082 579771 312085
rect 583520 312082 584960 312172
rect 579705 312080 584960 312082
rect 579705 312024 579710 312080
rect 579766 312024 584960 312080
rect 579705 312022 584960 312024
rect 579705 312019 579771 312022
rect 583520 311932 584960 312022
rect -960 306234 480 306324
rect 3141 306234 3207 306237
rect -960 306232 3207 306234
rect -960 306176 3146 306232
rect 3202 306176 3207 306232
rect -960 306174 3207 306176
rect -960 306084 480 306174
rect 3141 306171 3207 306174
rect 579797 298754 579863 298757
rect 583520 298754 584960 298844
rect 579797 298752 584960 298754
rect 579797 298696 579802 298752
rect 579858 298696 584960 298752
rect 579797 298694 584960 298696
rect 579797 298691 579863 298694
rect 583520 298604 584960 298694
rect -960 293178 480 293268
rect 565 293178 631 293181
rect -960 293176 631 293178
rect -960 293120 570 293176
rect 626 293120 631 293176
rect -960 293118 631 293120
rect -960 293028 480 293118
rect 565 293115 631 293118
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 580165 272234 580231 272237
rect 583520 272234 584960 272324
rect 580165 272232 584960 272234
rect 580165 272176 580170 272232
rect 580226 272176 584960 272232
rect 580165 272174 584960 272176
rect 580165 272171 580231 272174
rect 583520 272084 584960 272174
rect -960 267202 480 267292
rect 565 267202 631 267205
rect -960 267200 631 267202
rect -960 267144 570 267200
rect 626 267144 631 267200
rect -960 267142 631 267144
rect -960 267052 480 267142
rect 565 267139 631 267142
rect 580441 258906 580507 258909
rect 583520 258906 584960 258996
rect 580441 258904 584960 258906
rect 580441 258848 580446 258904
rect 580502 258848 584960 258904
rect 580441 258846 584960 258848
rect 580441 258843 580507 258846
rect 583520 258756 584960 258846
rect -960 254146 480 254236
rect 565 254146 631 254149
rect -960 254144 631 254146
rect -960 254088 570 254144
rect 626 254088 631 254144
rect -960 254086 631 254088
rect -960 253996 480 254086
rect 565 254083 631 254086
rect 580165 245578 580231 245581
rect 583520 245578 584960 245668
rect 580165 245576 584960 245578
rect 580165 245520 580170 245576
rect 580226 245520 584960 245576
rect 580165 245518 584960 245520
rect 580165 245515 580231 245518
rect 583520 245428 584960 245518
rect -960 241090 480 241180
rect 3969 241090 4035 241093
rect -960 241088 4035 241090
rect -960 241032 3974 241088
rect 4030 241032 4035 241088
rect -960 241030 4035 241032
rect -960 240940 480 241030
rect 3969 241027 4035 241030
rect 580165 232386 580231 232389
rect 583520 232386 584960 232476
rect 580165 232384 584960 232386
rect 580165 232328 580170 232384
rect 580226 232328 584960 232384
rect 580165 232326 584960 232328
rect 580165 232323 580231 232326
rect 583520 232236 584960 232326
rect -960 227884 480 228124
rect 580165 219058 580231 219061
rect 583520 219058 584960 219148
rect 580165 219056 584960 219058
rect 580165 219000 580170 219056
rect 580226 219000 584960 219056
rect 580165 218998 584960 219000
rect 580165 218995 580231 218998
rect 583520 218908 584960 218998
rect -960 214978 480 215068
rect 2129 214978 2195 214981
rect -960 214976 2195 214978
rect -960 214920 2134 214976
rect 2190 214920 2195 214976
rect -960 214918 2195 214920
rect -960 214828 480 214918
rect 2129 214915 2195 214918
rect 579889 205730 579955 205733
rect 583520 205730 584960 205820
rect 579889 205728 584960 205730
rect 579889 205672 579894 205728
rect 579950 205672 584960 205728
rect 579889 205670 584960 205672
rect 579889 205667 579955 205670
rect 583520 205580 584960 205670
rect -960 201922 480 202012
rect 3877 201922 3943 201925
rect -960 201920 3943 201922
rect -960 201864 3882 201920
rect 3938 201864 3943 201920
rect -960 201862 3943 201864
rect -960 201772 480 201862
rect 3877 201859 3943 201862
rect 580165 192538 580231 192541
rect 583520 192538 584960 192628
rect 580165 192536 584960 192538
rect 580165 192480 580170 192536
rect 580226 192480 584960 192536
rect 580165 192478 584960 192480
rect 580165 192475 580231 192478
rect 583520 192388 584960 192478
rect -960 188866 480 188956
rect 2221 188866 2287 188869
rect -960 188864 2287 188866
rect -960 188808 2226 188864
rect 2282 188808 2287 188864
rect -960 188806 2287 188808
rect -960 188716 480 188806
rect 2221 188803 2287 188806
rect 580349 179210 580415 179213
rect 583520 179210 584960 179300
rect 580349 179208 584960 179210
rect 580349 179152 580354 179208
rect 580410 179152 584960 179208
rect 580349 179150 584960 179152
rect 580349 179147 580415 179150
rect 583520 179060 584960 179150
rect -960 175796 480 176036
rect 580165 165882 580231 165885
rect 583520 165882 584960 165972
rect 580165 165880 584960 165882
rect 580165 165824 580170 165880
rect 580226 165824 584960 165880
rect 580165 165822 584960 165824
rect 580165 165819 580231 165822
rect 583520 165732 584960 165822
rect -960 162890 480 162980
rect 565 162890 631 162893
rect -960 162888 631 162890
rect -960 162832 570 162888
rect 626 162832 631 162888
rect -960 162830 631 162832
rect -960 162740 480 162830
rect 565 162827 631 162830
rect 579797 152690 579863 152693
rect 583520 152690 584960 152780
rect 579797 152688 584960 152690
rect 579797 152632 579802 152688
rect 579858 152632 584960 152688
rect 579797 152630 584960 152632
rect 579797 152627 579863 152630
rect 583520 152540 584960 152630
rect -960 149834 480 149924
rect 3785 149834 3851 149837
rect -960 149832 3851 149834
rect -960 149776 3790 149832
rect 3846 149776 3851 149832
rect -960 149774 3851 149776
rect -960 149684 480 149774
rect 3785 149771 3851 149774
rect 580165 139362 580231 139365
rect 583520 139362 584960 139452
rect 580165 139360 584960 139362
rect 580165 139304 580170 139360
rect 580226 139304 584960 139360
rect 580165 139302 584960 139304
rect 580165 139299 580231 139302
rect 583520 139212 584960 139302
rect -960 136778 480 136868
rect 3693 136778 3759 136781
rect -960 136776 3759 136778
rect -960 136720 3698 136776
rect 3754 136720 3759 136776
rect -960 136718 3759 136720
rect -960 136628 480 136718
rect 3693 136715 3759 136718
rect 580165 126034 580231 126037
rect 583520 126034 584960 126124
rect 580165 126032 584960 126034
rect 580165 125976 580170 126032
rect 580226 125976 584960 126032
rect 580165 125974 584960 125976
rect 580165 125971 580231 125974
rect 583520 125884 584960 125974
rect -960 123572 480 123812
rect 580165 112842 580231 112845
rect 583520 112842 584960 112932
rect 580165 112840 584960 112842
rect 580165 112784 580170 112840
rect 580226 112784 584960 112840
rect 580165 112782 584960 112784
rect 580165 112779 580231 112782
rect 583520 112692 584960 112782
rect 197 111210 263 111213
rect 197 111208 306 111210
rect 197 111152 202 111208
rect 258 111152 306 111208
rect 197 111147 306 111152
rect 246 110802 306 111147
rect 246 110756 674 110802
rect -960 110742 674 110756
rect -960 110666 480 110742
rect 614 110666 674 110742
rect -960 110606 674 110666
rect -960 110516 480 110606
rect 580165 99514 580231 99517
rect 583520 99514 584960 99604
rect 580165 99512 584960 99514
rect 580165 99456 580170 99512
rect 580226 99456 584960 99512
rect 580165 99454 584960 99456
rect 580165 99451 580231 99454
rect 583520 99364 584960 99454
rect -960 97610 480 97700
rect 3601 97610 3667 97613
rect -960 97608 3667 97610
rect -960 97552 3606 97608
rect 3662 97552 3667 97608
rect -960 97550 3667 97552
rect -960 97460 480 97550
rect 3601 97547 3667 97550
rect 580165 86186 580231 86189
rect 583520 86186 584960 86276
rect 580165 86184 584960 86186
rect 580165 86128 580170 86184
rect 580226 86128 584960 86184
rect 580165 86126 584960 86128
rect 580165 86123 580231 86126
rect 583520 86036 584960 86126
rect 105 85234 171 85237
rect 105 85232 306 85234
rect 105 85176 110 85232
rect 166 85176 306 85232
rect 105 85174 306 85176
rect 105 85171 171 85174
rect 246 84826 306 85174
rect 246 84780 674 84826
rect -960 84766 674 84780
rect -960 84690 480 84766
rect 614 84690 674 84766
rect -960 84630 674 84690
rect -960 84540 480 84630
rect 579981 72994 580047 72997
rect 583520 72994 584960 73084
rect 579981 72992 584960 72994
rect 579981 72936 579986 72992
rect 580042 72936 584960 72992
rect 579981 72934 584960 72936
rect 579981 72931 580047 72934
rect 583520 72844 584960 72934
rect 13 71906 79 71909
rect 13 71904 122 71906
rect 13 71848 18 71904
rect 74 71848 122 71904
rect 13 71843 122 71848
rect 62 71770 122 71843
rect 62 71724 674 71770
rect -960 71710 674 71724
rect -960 71634 480 71710
rect 614 71634 674 71710
rect -960 71574 674 71634
rect -960 71484 480 71574
rect 580165 59666 580231 59669
rect 583520 59666 584960 59756
rect 580165 59664 584960 59666
rect 580165 59608 580170 59664
rect 580226 59608 584960 59664
rect 580165 59606 584960 59608
rect 580165 59603 580231 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 2037 58578 2103 58581
rect -960 58576 2103 58578
rect -960 58520 2042 58576
rect 2098 58520 2103 58576
rect -960 58518 2103 58520
rect -960 58428 480 58518
rect 2037 58515 2103 58518
rect 580165 46338 580231 46341
rect 583520 46338 584960 46428
rect 580165 46336 584960 46338
rect 580165 46280 580170 46336
rect 580226 46280 584960 46336
rect 580165 46278 584960 46280
rect 580165 46275 580231 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3509 45522 3575 45525
rect -960 45520 3575 45522
rect -960 45464 3514 45520
rect 3570 45464 3575 45520
rect -960 45462 3575 45464
rect -960 45372 480 45462
rect 3509 45459 3575 45462
rect 580165 33146 580231 33149
rect 583520 33146 584960 33236
rect 580165 33144 584960 33146
rect 580165 33088 580170 33144
rect 580226 33088 584960 33144
rect 580165 33086 584960 33088
rect 580165 33083 580231 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 4061 32466 4127 32469
rect -960 32464 4127 32466
rect -960 32408 4066 32464
rect 4122 32408 4127 32464
rect -960 32406 4127 32408
rect -960 32316 480 32406
rect 4061 32403 4127 32406
rect 579705 19818 579771 19821
rect 583520 19818 584960 19908
rect 579705 19816 584960 19818
rect 579705 19760 579710 19816
rect 579766 19760 584960 19816
rect 579705 19758 584960 19760
rect 579705 19755 579771 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 580257 6626 580323 6629
rect 583520 6626 584960 6716
rect 580257 6624 584960 6626
rect -960 6490 480 6580
rect 580257 6568 580262 6624
rect 580318 6568 584960 6624
rect 580257 6566 584960 6568
rect 580257 6563 580323 6566
rect 2957 6490 3023 6493
rect -960 6488 3023 6490
rect -960 6432 2962 6488
rect 3018 6432 3023 6488
rect 583520 6476 584960 6566
rect -960 6430 3023 6432
rect -960 6340 480 6430
rect 2957 6427 3023 6430
rect 531262 1458 531268 1460
rect 514710 1398 531268 1458
rect 514710 645 514770 1398
rect 531262 1396 531268 1398
rect 531332 1396 531338 1460
rect 559414 914 559420 916
rect 542310 854 559420 914
rect 8753 642 8819 645
rect 9949 642 10015 645
rect 13261 642 13327 645
rect 8753 640 8954 642
rect 8753 584 8758 640
rect 8814 584 8954 640
rect 8753 582 8954 584
rect 8753 579 8819 582
rect 8894 506 8954 582
rect 9949 640 13327 642
rect 9949 584 9954 640
rect 10010 584 13266 640
rect 13322 584 13327 640
rect 9949 582 13327 584
rect 9949 579 10015 582
rect 13261 579 13327 582
rect 20621 642 20687 645
rect 23473 642 23539 645
rect 20621 640 23539 642
rect 20621 584 20626 640
rect 20682 584 23478 640
rect 23534 584 23539 640
rect 20621 582 23539 584
rect 20621 579 20687 582
rect 23473 579 23539 582
rect 26509 642 26575 645
rect 28717 642 28783 645
rect 30281 642 30347 645
rect 26509 640 28783 642
rect 26509 584 26514 640
rect 26570 584 28722 640
rect 28778 584 28783 640
rect 26509 582 28783 584
rect 26509 579 26575 582
rect 28717 579 28783 582
rect 29134 640 30347 642
rect 29134 584 30286 640
rect 30342 584 30347 640
rect 29134 582 30347 584
rect 12617 506 12683 509
rect 8894 504 12683 506
rect 8894 448 12622 504
rect 12678 448 12683 504
rect 8894 446 12683 448
rect 12617 443 12683 446
rect 27889 506 27955 509
rect 29134 506 29194 582
rect 30281 579 30347 582
rect 34789 642 34855 645
rect 35985 642 36051 645
rect 38469 642 38535 645
rect 34789 640 34898 642
rect 34789 584 34794 640
rect 34850 584 34898 640
rect 34789 579 34898 584
rect 35985 640 38535 642
rect 35985 584 35990 640
rect 36046 584 38474 640
rect 38530 584 38535 640
rect 35985 582 38535 584
rect 35985 579 36051 582
rect 38469 579 38535 582
rect 52545 642 52611 645
rect 54201 642 54267 645
rect 52545 640 54267 642
rect 52545 584 52550 640
rect 52606 584 54206 640
rect 54262 584 54267 640
rect 52545 582 54267 584
rect 52545 579 52611 582
rect 54201 579 54267 582
rect 56041 642 56107 645
rect 57605 642 57671 645
rect 56041 640 57671 642
rect 56041 584 56046 640
rect 56102 584 57610 640
rect 57666 584 57671 640
rect 56041 582 57671 584
rect 56041 579 56107 582
rect 57605 579 57671 582
rect 58433 642 58499 645
rect 59813 642 59879 645
rect 58433 640 59879 642
rect 58433 584 58438 640
rect 58494 584 59818 640
rect 59874 584 59879 640
rect 58433 582 59879 584
rect 58433 579 58499 582
rect 59813 579 59879 582
rect 60825 642 60891 645
rect 62113 642 62179 645
rect 60825 640 62179 642
rect 60825 584 60830 640
rect 60886 584 62118 640
rect 62174 584 62179 640
rect 60825 582 62179 584
rect 60825 579 60891 582
rect 62113 579 62179 582
rect 142061 642 142127 645
rect 143441 642 143507 645
rect 144729 642 144795 645
rect 142061 640 142170 642
rect 142061 584 142066 640
rect 142122 584 142170 640
rect 142061 579 142170 584
rect 143441 640 144795 642
rect 143441 584 143446 640
rect 143502 584 144734 640
rect 144790 584 144795 640
rect 143441 582 144795 584
rect 143441 579 143507 582
rect 144729 579 144795 582
rect 145741 642 145807 645
rect 147121 642 147187 645
rect 145741 640 147187 642
rect 145741 584 145746 640
rect 145802 584 147126 640
rect 147182 584 147187 640
rect 145741 582 147187 584
rect 145741 579 145807 582
rect 147121 579 147187 582
rect 148961 642 149027 645
rect 150617 642 150683 645
rect 151813 642 151879 645
rect 148961 640 150683 642
rect 148961 584 148966 640
rect 149022 584 150622 640
rect 150678 584 150683 640
rect 148961 582 150683 584
rect 148961 579 149027 582
rect 150617 579 150683 582
rect 151678 640 151879 642
rect 151678 584 151818 640
rect 151874 584 151879 640
rect 151678 582 151879 584
rect 27889 504 29194 506
rect 27889 448 27894 504
rect 27950 448 29194 504
rect 27889 446 29194 448
rect 34838 506 34898 579
rect 37365 506 37431 509
rect 34838 504 37431 506
rect 34838 448 37370 504
rect 37426 448 37431 504
rect 34838 446 37431 448
rect 27889 443 27955 446
rect 37365 443 37431 446
rect 53557 506 53623 509
rect 55305 506 55371 509
rect 53557 504 55371 506
rect 53557 448 53562 504
rect 53618 448 55310 504
rect 55366 448 55371 504
rect 53557 446 55371 448
rect 53557 443 53623 446
rect 55305 443 55371 446
rect 57421 506 57487 509
rect 58801 506 58867 509
rect 57421 504 58867 506
rect 57421 448 57426 504
rect 57482 448 58806 504
rect 58862 448 58867 504
rect 57421 446 58867 448
rect 57421 443 57487 446
rect 58801 443 58867 446
rect 59445 506 59511 509
rect 61101 506 61167 509
rect 59445 504 61167 506
rect 59445 448 59450 504
rect 59506 448 61106 504
rect 61162 448 61167 504
rect 59445 446 61167 448
rect 142110 506 142170 579
rect 143717 506 143783 509
rect 142110 504 143783 506
rect 142110 448 143722 504
rect 143778 448 143783 504
rect 142110 446 143783 448
rect 59445 443 59511 446
rect 61101 443 61167 446
rect 143717 443 143783 446
rect 147765 506 147831 509
rect 149329 506 149395 509
rect 147765 504 149395 506
rect 147765 448 147770 504
rect 147826 448 149334 504
rect 149390 448 149395 504
rect 147765 446 149395 448
rect 147765 443 147831 446
rect 149329 443 149395 446
rect 150249 506 150315 509
rect 151678 506 151738 582
rect 151813 579 151879 582
rect 164785 642 164851 645
rect 167361 642 167427 645
rect 164785 640 167427 642
rect 164785 584 164790 640
rect 164846 584 167366 640
rect 167422 584 167427 640
rect 164785 582 167427 584
rect 164785 579 164851 582
rect 167361 579 167427 582
rect 169477 642 169543 645
rect 171961 642 172027 645
rect 169477 640 172027 642
rect 169477 584 169482 640
rect 169538 584 171966 640
rect 172022 584 172027 640
rect 169477 582 172027 584
rect 169477 579 169543 582
rect 171961 579 172027 582
rect 172973 642 173039 645
rect 175457 642 175523 645
rect 172973 640 175523 642
rect 172973 584 172978 640
rect 173034 584 175462 640
rect 175518 584 175523 640
rect 172973 582 175523 584
rect 172973 579 173039 582
rect 175457 579 175523 582
rect 176377 642 176443 645
rect 179045 642 179111 645
rect 180241 642 180307 645
rect 176377 640 179111 642
rect 176377 584 176382 640
rect 176438 584 179050 640
rect 179106 584 179111 640
rect 176377 582 179111 584
rect 176377 579 176443 582
rect 179045 579 179111 582
rect 179370 640 180307 642
rect 179370 584 180246 640
rect 180302 584 180307 640
rect 179370 582 180307 584
rect 150249 504 151738 506
rect 150249 448 150254 504
rect 150310 448 151738 504
rect 150249 446 151738 448
rect 173893 506 173959 509
rect 176837 506 176903 509
rect 173893 504 176903 506
rect 173893 448 173898 504
rect 173954 448 176842 504
rect 176898 448 176903 504
rect 173893 446 176903 448
rect 150249 443 150315 446
rect 173893 443 173959 446
rect 176837 443 176903 446
rect 177481 506 177547 509
rect 179370 506 179430 582
rect 180241 579 180307 582
rect 182081 642 182147 645
rect 184933 642 184999 645
rect 182081 640 184999 642
rect 182081 584 182086 640
rect 182142 584 184938 640
rect 184994 584 184999 640
rect 182081 582 184999 584
rect 182081 579 182147 582
rect 184933 579 184999 582
rect 192293 642 192359 645
rect 195605 642 195671 645
rect 197905 642 197971 645
rect 192293 640 195671 642
rect 192293 584 192298 640
rect 192354 584 195610 640
rect 195666 584 195671 640
rect 192293 582 195671 584
rect 192293 579 192359 582
rect 195605 579 195671 582
rect 197310 640 197971 642
rect 197310 584 197910 640
rect 197966 584 197971 640
rect 197310 582 197971 584
rect 177481 504 179430 506
rect 177481 448 177486 504
rect 177542 448 179430 504
rect 177481 446 179430 448
rect 186589 506 186655 509
rect 189901 506 189967 509
rect 186589 504 189967 506
rect 186589 448 186594 504
rect 186650 448 189906 504
rect 189962 448 189967 504
rect 186589 446 189967 448
rect 177481 443 177547 446
rect 186589 443 186655 446
rect 189901 443 189967 446
rect 194041 506 194107 509
rect 197310 506 197370 582
rect 197905 579 197971 582
rect 200021 642 200087 645
rect 203885 642 203951 645
rect 200021 640 203951 642
rect 200021 584 200026 640
rect 200082 584 203890 640
rect 203946 584 203951 640
rect 200021 582 203951 584
rect 200021 579 200087 582
rect 203885 579 203951 582
rect 204161 642 204227 645
rect 207381 642 207447 645
rect 204161 640 207447 642
rect 204161 584 204166 640
rect 204222 584 207386 640
rect 207442 584 207447 640
rect 204161 582 207447 584
rect 204161 579 204227 582
rect 207381 579 207447 582
rect 208209 642 208275 645
rect 208393 642 208459 645
rect 208209 640 208459 642
rect 208209 584 208214 640
rect 208270 584 208398 640
rect 208454 584 208459 640
rect 208209 582 208459 584
rect 208209 579 208275 582
rect 208393 579 208459 582
rect 209313 642 209379 645
rect 213361 642 213427 645
rect 209313 640 213427 642
rect 209313 584 209318 640
rect 209374 584 213366 640
rect 213422 584 213427 640
rect 209313 582 213427 584
rect 209313 579 209379 582
rect 213361 579 213427 582
rect 216121 642 216187 645
rect 220721 642 220787 645
rect 216121 640 220787 642
rect 216121 584 216126 640
rect 216182 584 220726 640
rect 220782 584 220787 640
rect 216121 582 220787 584
rect 216121 579 216187 582
rect 220721 579 220787 582
rect 221825 642 221891 645
rect 226333 642 226399 645
rect 228725 642 228791 645
rect 221825 640 226399 642
rect 221825 584 221830 640
rect 221886 584 226338 640
rect 226394 584 226399 640
rect 221825 582 226399 584
rect 221825 579 221891 582
rect 226333 579 226399 582
rect 227670 640 228791 642
rect 227670 584 228730 640
rect 228786 584 228791 640
rect 227670 582 228791 584
rect 194041 504 197370 506
rect 194041 448 194046 504
rect 194102 448 197370 504
rect 194041 446 197370 448
rect 198917 506 198983 509
rect 201309 506 201375 509
rect 204897 506 204963 509
rect 198917 504 200866 506
rect 198917 448 198922 504
rect 198978 448 200866 504
rect 198917 446 200866 448
rect 194041 443 194107 446
rect 198917 443 198983 446
rect 168189 370 168255 373
rect 170949 370 171015 373
rect 168189 368 171015 370
rect 168189 312 168194 368
rect 168250 312 170954 368
rect 171010 312 171015 368
rect 168189 310 171015 312
rect 168189 307 168255 310
rect 170949 307 171015 310
rect 171685 370 171751 373
rect 173985 370 174051 373
rect 171685 368 174051 370
rect 171685 312 171690 368
rect 171746 312 173990 368
rect 174046 312 174051 368
rect 171685 310 174051 312
rect 171685 307 171751 310
rect 173985 307 174051 310
rect 175181 370 175247 373
rect 177665 370 177731 373
rect 175181 368 177731 370
rect 175181 312 175186 368
rect 175242 312 177670 368
rect 177726 312 177731 368
rect 175181 310 177731 312
rect 175181 307 175247 310
rect 177665 307 177731 310
rect 178677 370 178743 373
rect 181253 370 181319 373
rect 178677 368 181319 370
rect 178677 312 178682 368
rect 178738 312 181258 368
rect 181314 312 181319 368
rect 178677 310 181319 312
rect 178677 307 178743 310
rect 181253 307 181319 310
rect 196617 370 196683 373
rect 200113 370 200179 373
rect 196617 368 200179 370
rect 196617 312 196622 368
rect 196678 312 200118 368
rect 200174 312 200179 368
rect 196617 310 200179 312
rect 200806 370 200866 446
rect 201309 504 204963 506
rect 201309 448 201314 504
rect 201370 448 204902 504
rect 204958 448 204963 504
rect 201309 446 204963 448
rect 201309 443 201375 446
rect 204897 443 204963 446
rect 206921 506 206987 509
rect 210785 506 210851 509
rect 206921 504 210851 506
rect 206921 448 206926 504
rect 206982 448 210790 504
rect 210846 448 210851 504
rect 206921 446 210851 448
rect 206921 443 206987 446
rect 210785 443 210851 446
rect 223573 506 223639 509
rect 227670 506 227730 582
rect 228725 579 228791 582
rect 230933 642 230999 645
rect 235809 642 235875 645
rect 230933 640 235875 642
rect 230933 584 230938 640
rect 230994 584 235814 640
rect 235870 584 235875 640
rect 230933 582 235875 584
rect 230933 579 230999 582
rect 235809 579 235875 582
rect 237741 642 237807 645
rect 242893 642 242959 645
rect 237741 640 242959 642
rect 237741 584 237746 640
rect 237802 584 242898 640
rect 242954 584 242959 640
rect 237741 582 242959 584
rect 237741 579 237807 582
rect 242893 579 242959 582
rect 249701 642 249767 645
rect 255865 642 255931 645
rect 249701 640 255931 642
rect 249701 584 249706 640
rect 249762 584 255870 640
rect 255926 584 255931 640
rect 249701 582 255931 584
rect 249701 579 249767 582
rect 255865 579 255931 582
rect 267273 642 267339 645
rect 273621 642 273687 645
rect 267273 640 273687 642
rect 267273 584 267278 640
rect 267334 584 273626 640
rect 273682 584 273687 640
rect 267273 582 273687 584
rect 267273 579 267339 582
rect 273621 579 273687 582
rect 275185 642 275251 645
rect 282085 642 282151 645
rect 275185 640 282151 642
rect 275185 584 275190 640
rect 275246 584 282090 640
rect 282146 584 282151 640
rect 275185 582 282151 584
rect 275185 579 275251 582
rect 282085 579 282151 582
rect 285673 642 285739 645
rect 287789 642 287855 645
rect 292573 642 292639 645
rect 285673 640 287855 642
rect 285673 584 285678 640
rect 285734 584 287794 640
rect 287850 584 287855 640
rect 285673 582 287855 584
rect 285673 579 285739 582
rect 287789 579 287855 582
rect 288758 640 292639 642
rect 288758 584 292578 640
rect 292634 584 292639 640
rect 288758 582 292639 584
rect 223573 504 227730 506
rect 223573 448 223578 504
rect 223634 448 227730 504
rect 223573 446 227730 448
rect 242249 506 242315 509
rect 247309 506 247375 509
rect 242249 504 247375 506
rect 242249 448 242254 504
rect 242310 448 247314 504
rect 247370 448 247375 504
rect 242249 446 247375 448
rect 223573 443 223639 446
rect 242249 443 242315 446
rect 247309 443 247375 446
rect 285213 506 285279 509
rect 288758 506 288818 582
rect 292573 579 292639 582
rect 294597 642 294663 645
rect 296069 642 296135 645
rect 294597 640 296135 642
rect 294597 584 294602 640
rect 294658 584 296074 640
rect 296130 584 296135 640
rect 294597 582 296135 584
rect 294597 579 294663 582
rect 296069 579 296135 582
rect 305821 642 305887 645
rect 313825 642 313891 645
rect 305821 640 313891 642
rect 305821 584 305826 640
rect 305882 584 313830 640
rect 313886 584 313891 640
rect 305821 582 313891 584
rect 305821 579 305887 582
rect 313825 579 313891 582
rect 315021 640 315087 645
rect 315021 584 315026 640
rect 315082 584 315087 640
rect 315021 579 315087 584
rect 316585 642 316651 645
rect 317321 642 317387 645
rect 316585 640 317387 642
rect 316585 584 316590 640
rect 316646 584 317326 640
rect 317382 584 317387 640
rect 316585 582 317387 584
rect 316585 579 316651 582
rect 317321 579 317387 582
rect 328453 642 328519 645
rect 337469 642 337535 645
rect 343357 642 343423 645
rect 328453 640 337535 642
rect 328453 584 328458 640
rect 328514 584 337474 640
rect 337530 584 337535 640
rect 328453 582 337535 584
rect 328453 579 328519 582
rect 337469 579 337535 582
rect 340830 640 343423 642
rect 340830 584 343362 640
rect 343418 584 343423 640
rect 340830 582 343423 584
rect 285213 504 288818 506
rect 285213 448 285218 504
rect 285274 448 288818 504
rect 285213 446 288818 448
rect 307017 506 307083 509
rect 315024 506 315084 579
rect 307017 504 315084 506
rect 307017 448 307022 504
rect 307078 448 315084 504
rect 307017 446 315084 448
rect 334249 506 334315 509
rect 340830 506 340890 582
rect 343357 579 343423 582
rect 345013 642 345079 645
rect 346945 642 347011 645
rect 345013 640 347011 642
rect 345013 584 345018 640
rect 345074 584 346950 640
rect 347006 584 347011 640
rect 345013 582 347011 584
rect 345013 579 345079 582
rect 346945 579 347011 582
rect 349061 642 349127 645
rect 350441 642 350507 645
rect 349061 640 350507 642
rect 349061 584 349066 640
rect 349122 584 350446 640
rect 350502 584 350507 640
rect 349061 582 350507 584
rect 349061 579 349127 582
rect 350441 579 350507 582
rect 350625 642 350691 645
rect 352833 642 352899 645
rect 359917 642 359983 645
rect 350625 640 352899 642
rect 350625 584 350630 640
rect 350686 584 352838 640
rect 352894 584 352899 640
rect 350625 582 352899 584
rect 350625 579 350691 582
rect 352833 579 352899 582
rect 353250 640 359983 642
rect 353250 584 359922 640
rect 359978 584 359983 640
rect 353250 582 359983 584
rect 347865 506 347931 509
rect 334249 504 340890 506
rect 334249 448 334254 504
rect 334310 448 340890 504
rect 334249 446 340890 448
rect 342210 504 347931 506
rect 342210 448 347870 504
rect 347926 448 347931 504
rect 342210 446 347931 448
rect 285213 443 285279 446
rect 307017 443 307083 446
rect 334249 443 334315 446
rect 202505 370 202571 373
rect 200806 368 202571 370
rect 200806 312 202510 368
rect 202566 312 202571 368
rect 200806 310 202571 312
rect 196617 307 196683 310
rect 200113 307 200179 310
rect 202505 307 202571 310
rect 204805 370 204871 373
rect 208761 370 208827 373
rect 204805 368 208827 370
rect 204805 312 204810 368
rect 204866 312 208766 368
rect 208822 312 208827 368
rect 204805 310 208827 312
rect 204805 307 204871 310
rect 208761 307 208827 310
rect 286409 370 286475 373
rect 293401 370 293467 373
rect 286409 368 293467 370
rect 286409 312 286414 368
rect 286470 312 293406 368
rect 293462 312 293467 368
rect 286409 310 293467 312
rect 286409 307 286475 310
rect 293401 307 293467 310
rect 338297 370 338363 373
rect 342210 370 342270 446
rect 347865 443 347931 446
rect 350165 506 350231 509
rect 353250 506 353310 582
rect 359917 579 359983 582
rect 363781 642 363847 645
rect 374085 642 374151 645
rect 363781 640 374151 642
rect 363781 584 363786 640
rect 363842 584 374090 640
rect 374146 584 374151 640
rect 363781 582 374151 584
rect 363781 579 363847 582
rect 374085 579 374151 582
rect 374269 642 374335 645
rect 377673 642 377739 645
rect 374269 640 377739 642
rect 374269 584 374274 640
rect 374330 584 377678 640
rect 377734 584 377739 640
rect 374269 582 377739 584
rect 374269 579 374335 582
rect 377673 579 377739 582
rect 377949 642 378015 645
rect 379973 642 380039 645
rect 377949 640 380039 642
rect 377949 584 377954 640
rect 378010 584 379978 640
rect 380034 584 380039 640
rect 377949 582 380039 584
rect 377949 579 378015 582
rect 379973 579 380039 582
rect 380157 642 380223 645
rect 382365 642 382431 645
rect 384757 642 384823 645
rect 380157 640 382431 642
rect 380157 584 380162 640
rect 380218 584 382370 640
rect 382426 584 382431 640
rect 380157 582 382431 584
rect 380157 579 380223 582
rect 382365 579 382431 582
rect 383610 640 384823 642
rect 383610 584 384762 640
rect 384818 584 384823 640
rect 383610 582 384823 584
rect 350165 504 353310 506
rect 350165 448 350170 504
rect 350226 448 353310 504
rect 350165 446 353310 448
rect 362677 506 362743 509
rect 372705 506 372771 509
rect 362677 504 372771 506
rect 362677 448 362682 504
rect 362738 448 372710 504
rect 372766 448 372771 504
rect 362677 446 372771 448
rect 350165 443 350231 446
rect 362677 443 362743 446
rect 372705 443 372771 446
rect 375649 506 375715 509
rect 378685 506 378751 509
rect 375649 504 378751 506
rect 375649 448 375654 504
rect 375710 448 378690 504
rect 378746 448 378751 504
rect 375649 446 378751 448
rect 375649 443 375715 446
rect 378685 443 378751 446
rect 380893 506 380959 509
rect 383610 506 383670 582
rect 384757 579 384823 582
rect 385401 642 385467 645
rect 396533 642 396599 645
rect 401409 642 401475 645
rect 385401 640 396599 642
rect 385401 584 385406 640
rect 385462 584 396538 640
rect 396594 584 396599 640
rect 385401 582 396599 584
rect 385401 579 385467 582
rect 396533 579 396599 582
rect 401366 640 401475 642
rect 401366 584 401414 640
rect 401470 584 401475 640
rect 401366 579 401475 584
rect 405825 642 405891 645
rect 409597 642 409663 645
rect 405825 640 409663 642
rect 405825 584 405830 640
rect 405886 584 409602 640
rect 409658 584 409663 640
rect 405825 582 409663 584
rect 405825 579 405891 582
rect 409597 579 409663 582
rect 412633 642 412699 645
rect 421741 642 421807 645
rect 427261 642 427327 645
rect 412633 640 416790 642
rect 412633 584 412638 640
rect 412694 584 416790 640
rect 412633 582 416790 584
rect 412633 579 412699 582
rect 380893 504 383670 506
rect 380893 448 380898 504
rect 380954 448 383670 504
rect 380893 446 383670 448
rect 392393 506 392459 509
rect 401366 506 401426 579
rect 392393 504 401426 506
rect 392393 448 392398 504
rect 392454 448 401426 504
rect 392393 446 401426 448
rect 416730 506 416790 582
rect 421741 640 427327 642
rect 421741 584 421746 640
rect 421802 584 427266 640
rect 427322 584 427327 640
rect 421741 582 427327 584
rect 421741 579 421807 582
rect 427261 579 427327 582
rect 429009 642 429075 645
rect 429653 642 429719 645
rect 429009 640 429719 642
rect 429009 584 429014 640
rect 429070 584 429658 640
rect 429714 584 429719 640
rect 429009 582 429719 584
rect 429009 579 429075 582
rect 429653 579 429719 582
rect 456057 642 456123 645
rect 460473 642 460539 645
rect 456057 640 460539 642
rect 456057 584 456062 640
rect 456118 584 460478 640
rect 460534 584 460539 640
rect 456057 582 460539 584
rect 456057 579 456123 582
rect 460473 579 460539 582
rect 462129 642 462195 645
rect 463969 642 464035 645
rect 462129 640 464035 642
rect 462129 584 462134 640
rect 462190 584 463974 640
rect 464030 584 464035 640
rect 462129 582 464035 584
rect 462129 579 462195 582
rect 463969 579 464035 582
rect 466085 642 466151 645
rect 467465 642 467531 645
rect 466085 640 467531 642
rect 466085 584 466090 640
rect 466146 584 467470 640
rect 467526 584 467531 640
rect 466085 582 467531 584
rect 466085 579 466151 582
rect 467465 579 467531 582
rect 470593 642 470659 645
rect 477401 642 477467 645
rect 470593 640 477467 642
rect 470593 584 470598 640
rect 470654 584 477406 640
rect 477462 584 477467 640
rect 470593 582 477467 584
rect 470593 579 470659 582
rect 477401 579 477467 582
rect 483197 642 483263 645
rect 488809 642 488875 645
rect 483197 640 488875 642
rect 483197 584 483202 640
rect 483258 584 488814 640
rect 488870 584 488875 640
rect 483197 582 488875 584
rect 483197 579 483263 582
rect 488809 579 488875 582
rect 491293 642 491359 645
rect 495893 642 495959 645
rect 491293 640 495959 642
rect 491293 584 491298 640
rect 491354 584 495898 640
rect 495954 584 495959 640
rect 498009 642 498075 645
rect 500585 642 500651 645
rect 498009 640 500651 642
rect 497089 608 497155 611
rect 491293 582 495959 584
rect 491293 579 491359 582
rect 495893 579 495959 582
rect 497046 606 497155 608
rect 497046 550 497094 606
rect 497150 550 497155 606
rect 498009 584 498014 640
rect 498070 584 500590 640
rect 500646 584 500651 640
rect 498009 582 500651 584
rect 498009 579 498075 582
rect 500585 579 500651 582
rect 514661 640 514770 645
rect 518341 642 518407 645
rect 531313 644 531379 645
rect 514661 584 514666 640
rect 514722 584 514770 640
rect 514661 582 514770 584
rect 518206 640 518407 642
rect 518206 584 518346 640
rect 518402 584 518407 640
rect 518206 582 518407 584
rect 514661 579 514727 582
rect 497046 545 497155 550
rect 424501 506 424567 509
rect 416730 504 424567 506
rect 416730 448 424506 504
rect 424562 448 424567 504
rect 416730 446 424567 448
rect 380893 443 380959 446
rect 392393 443 392459 446
rect 424501 443 424567 446
rect 468293 506 468359 509
rect 476573 506 476639 509
rect 468293 504 476639 506
rect 468293 448 468298 504
rect 468354 448 476578 504
rect 476634 448 476639 504
rect 468293 446 476639 448
rect 468293 443 468359 446
rect 476573 443 476639 446
rect 493317 506 493383 509
rect 497046 506 497106 545
rect 493317 504 497106 506
rect 493317 448 493322 504
rect 493378 448 497106 504
rect 493317 446 497106 448
rect 509693 506 509759 509
rect 518206 506 518266 582
rect 518341 579 518407 582
rect 531262 580 531268 644
rect 531332 642 531379 644
rect 541709 642 541775 645
rect 542310 642 542370 854
rect 559414 852 559420 854
rect 559484 852 559490 916
rect 543230 718 557550 778
rect 531332 640 531424 642
rect 531374 584 531424 640
rect 531332 582 531424 584
rect 541709 640 542370 642
rect 541709 584 541714 640
rect 541770 584 542370 640
rect 541709 582 542370 584
rect 543089 642 543155 645
rect 543230 642 543290 718
rect 543089 640 543290 642
rect 543089 584 543094 640
rect 543150 584 543290 640
rect 543089 582 543290 584
rect 543457 642 543523 645
rect 554957 642 555023 645
rect 543457 640 555023 642
rect 543457 584 543462 640
rect 543518 584 554962 640
rect 555018 584 555023 640
rect 543457 582 555023 584
rect 531332 580 531379 582
rect 531313 579 531379 580
rect 541709 579 541775 582
rect 543089 579 543155 582
rect 543457 579 543523 582
rect 554957 579 555023 582
rect 555141 642 555207 645
rect 556153 642 556219 645
rect 555141 640 556219 642
rect 555141 584 555146 640
rect 555202 584 556158 640
rect 556214 584 556219 640
rect 555141 582 556219 584
rect 557490 642 557550 718
rect 560845 642 560911 645
rect 557490 640 560911 642
rect 557490 584 560850 640
rect 560906 584 560911 640
rect 557490 582 560911 584
rect 555141 579 555207 582
rect 556153 579 556219 582
rect 560845 579 560911 582
rect 509693 504 518266 506
rect 509693 448 509698 504
rect 509754 448 518266 504
rect 509693 446 518266 448
rect 540513 506 540579 509
rect 558361 506 558427 509
rect 540513 504 558427 506
rect 540513 448 540518 504
rect 540574 448 558366 504
rect 558422 448 558427 504
rect 540513 446 558427 448
rect 493317 443 493383 446
rect 509693 443 509759 446
rect 540513 443 540579 446
rect 558361 443 558427 446
rect 559414 444 559420 508
rect 559484 506 559490 508
rect 559557 506 559623 509
rect 559484 504 559623 506
rect 559484 448 559562 504
rect 559618 448 559623 504
rect 559484 446 559623 448
rect 559484 444 559490 446
rect 559557 443 559623 446
rect 338297 368 342270 370
rect 338297 312 338302 368
rect 338358 312 342270 368
rect 338297 310 342270 312
rect 361481 370 361547 373
rect 371969 370 372035 373
rect 361481 368 372035 370
rect 361481 312 361486 368
rect 361542 312 371974 368
rect 372030 312 372035 368
rect 361481 310 372035 312
rect 338297 307 338363 310
rect 361481 307 361547 310
rect 371969 307 372035 310
rect 392209 370 392275 373
rect 400305 370 400371 373
rect 392209 368 400371 370
rect 392209 312 392214 368
rect 392270 312 400310 368
rect 400366 312 400371 368
rect 392209 310 400371 312
rect 392209 307 392275 310
rect 400305 307 400371 310
rect 405089 370 405155 373
rect 408217 370 408283 373
rect 405089 368 408283 370
rect 405089 312 405094 368
rect 405150 312 408222 368
rect 408278 312 408283 368
rect 405089 310 408283 312
rect 405089 307 405155 310
rect 408217 307 408283 310
rect 446673 370 446739 373
rect 451917 370 451983 373
rect 446673 368 451983 370
rect 446673 312 446678 368
rect 446734 312 451922 368
rect 451978 312 451983 368
rect 446673 310 451983 312
rect 446673 307 446739 310
rect 451917 307 451983 310
rect 492673 370 492739 373
rect 493777 370 493843 373
rect 492673 368 493843 370
rect 492673 312 492678 368
rect 492734 312 493782 368
rect 493838 312 493843 368
rect 492673 310 493843 312
rect 492673 307 492739 310
rect 493777 307 493843 310
rect 508589 370 508655 373
rect 517329 370 517395 373
rect 508589 368 517395 370
rect 508589 312 508594 368
rect 508650 312 517334 368
rect 517390 312 517395 368
rect 508589 310 517395 312
rect 508589 307 508655 310
rect 517329 307 517395 310
rect 527173 370 527239 373
rect 544561 370 544627 373
rect 527173 368 544627 370
rect 527173 312 527178 368
rect 527234 312 544566 368
rect 544622 312 544627 368
rect 527173 310 544627 312
rect 527173 307 527239 310
rect 544561 307 544627 310
rect 202413 234 202479 237
rect 206001 234 206067 237
rect 202413 232 206067 234
rect 202413 176 202418 232
rect 202474 176 206006 232
rect 206062 176 206067 232
rect 202413 174 206067 176
rect 202413 171 202479 174
rect 206001 171 206067 174
rect 483657 234 483723 237
rect 492489 234 492555 237
rect 483657 232 492555 234
rect 483657 176 483662 232
rect 483718 176 492494 232
rect 492550 176 492555 232
rect 483657 174 492555 176
rect 483657 171 483723 174
rect 492489 171 492555 174
rect 534165 234 534231 237
rect 551277 234 551343 237
rect 534165 232 551343 234
rect 534165 176 534170 232
rect 534226 176 551282 232
rect 551338 176 551343 232
rect 534165 174 551343 176
rect 534165 171 534231 174
rect 551277 171 551343 174
rect 197721 98 197787 101
rect 201677 98 201743 101
rect 197721 96 201743 98
rect 197721 40 197726 96
rect 197782 40 201682 96
rect 201738 40 201743 96
rect 197721 38 201743 40
rect 197721 35 197787 38
rect 201677 35 201743 38
rect 530761 98 530827 101
rect 548057 98 548123 101
rect 530761 96 548123 98
rect 530761 40 530766 96
rect 530822 40 548062 96
rect 548118 40 548123 96
rect 530761 38 548123 40
rect 530761 35 530827 38
rect 548057 35 548123 38
<< via3 >>
rect 386276 702204 386340 702268
rect 259132 701116 259196 701180
rect 386276 699544 386340 699548
rect 386276 699488 386290 699544
rect 386290 699488 386340 699544
rect 386276 699484 386340 699488
rect 13860 699348 13924 699412
rect 95188 699408 95252 699412
rect 95188 699352 95202 699408
rect 95202 699352 95252 699408
rect 95188 699348 95252 699352
rect 418660 699408 418724 699412
rect 418660 699352 418710 699408
rect 418710 699352 418724 699408
rect 418660 699348 418724 699352
rect 433380 699408 433444 699412
rect 433380 699352 433430 699408
rect 433430 699352 433444 699408
rect 433380 699348 433444 699352
rect 462820 699408 462884 699412
rect 462820 699352 462870 699408
rect 462870 699352 462884 699408
rect 462820 699348 462884 699352
rect 492628 699408 492692 699412
rect 492628 699352 492642 699408
rect 492642 699352 492692 699408
rect 492628 699348 492692 699352
rect 539916 699348 539980 699412
rect 418844 699212 418908 699276
rect 259132 699076 259196 699140
rect 539916 698396 539980 698460
rect 13860 698260 13924 698324
rect 433380 698124 433444 698188
rect 418660 697988 418724 698052
rect 418844 697988 418908 698052
rect 462820 697852 462884 697916
rect 95188 697716 95252 697780
rect 492628 697580 492692 697644
rect 531268 1396 531332 1460
rect 531268 640 531332 644
rect 559420 852 559484 916
rect 531268 584 531318 640
rect 531318 584 531332 640
rect 531268 580 531332 584
rect 559420 444 559484 508
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 680614 -8106 711002
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 -8106 680614
rect -8726 680294 -8106 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 -8106 680294
rect -8726 644614 -8106 680058
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 -8106 644614
rect -8726 644294 -8106 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 -8106 644294
rect -8726 608614 -8106 644058
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 -8106 608614
rect -8726 608294 -8106 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 -8106 608294
rect -8726 572614 -8106 608058
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 -8106 572614
rect -8726 572294 -8106 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 -8106 572294
rect -8726 536614 -8106 572058
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 -8106 536614
rect -8726 536294 -8106 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 -8106 536294
rect -8726 500614 -8106 536058
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 -8106 500614
rect -8726 500294 -8106 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 -8106 500294
rect -8726 464614 -8106 500058
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 -8106 464614
rect -8726 464294 -8106 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 -8106 464294
rect -8726 428614 -8106 464058
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 -8106 428614
rect -8726 428294 -8106 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 -8106 428294
rect -8726 392614 -8106 428058
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 -8106 392614
rect -8726 392294 -8106 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 -8106 392294
rect -8726 356614 -8106 392058
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 -8106 356614
rect -8726 356294 -8106 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 -8106 356294
rect -8726 320614 -8106 356058
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 -8106 320614
rect -8726 320294 -8106 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 -8106 320294
rect -8726 284614 -8106 320058
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 -8106 284614
rect -8726 284294 -8106 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 -8106 284294
rect -8726 248614 -8106 284058
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 -8106 248614
rect -8726 248294 -8106 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 -8106 248294
rect -8726 212614 -8106 248058
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 -8106 212614
rect -8726 212294 -8106 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 -8106 212294
rect -8726 176614 -8106 212058
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 -8106 176614
rect -8726 176294 -8106 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 -8106 176294
rect -8726 140614 -8106 176058
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 -8106 140614
rect -8726 140294 -8106 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 -8106 140294
rect -8726 104614 -8106 140058
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 -8106 104614
rect -8726 104294 -8106 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 -8106 104294
rect -8726 68614 -8106 104058
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 -8106 68614
rect -8726 68294 -8106 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 -8106 68294
rect -8726 32614 -8106 68058
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 -8106 32614
rect -8726 32294 -8106 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 -8106 32294
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 13574 710598
rect 12954 710278 13574 710362
rect 12954 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 13574 710278
rect -7766 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 -7146 698614
rect -7766 698294 -7146 698378
rect -7766 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 -7146 698294
rect -7766 662614 -7146 698058
rect -7766 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 -7146 662614
rect -7766 662294 -7146 662378
rect -7766 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 -7146 662294
rect -7766 626614 -7146 662058
rect -7766 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 -7146 626614
rect -7766 626294 -7146 626378
rect -7766 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 -7146 626294
rect -7766 590614 -7146 626058
rect -7766 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 -7146 590614
rect -7766 590294 -7146 590378
rect -7766 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 -7146 590294
rect -7766 554614 -7146 590058
rect -7766 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 -7146 554614
rect -7766 554294 -7146 554378
rect -7766 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 -7146 554294
rect -7766 518614 -7146 554058
rect -7766 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 -7146 518614
rect -7766 518294 -7146 518378
rect -7766 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 -7146 518294
rect -7766 482614 -7146 518058
rect -7766 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 -7146 482614
rect -7766 482294 -7146 482378
rect -7766 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 -7146 482294
rect -7766 446614 -7146 482058
rect -7766 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 -7146 446614
rect -7766 446294 -7146 446378
rect -7766 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 -7146 446294
rect -7766 410614 -7146 446058
rect -7766 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 -7146 410614
rect -7766 410294 -7146 410378
rect -7766 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 -7146 410294
rect -7766 374614 -7146 410058
rect -7766 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 -7146 374614
rect -7766 374294 -7146 374378
rect -7766 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 -7146 374294
rect -7766 338614 -7146 374058
rect -7766 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 -7146 338614
rect -7766 338294 -7146 338378
rect -7766 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 -7146 338294
rect -7766 302614 -7146 338058
rect -7766 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 -7146 302614
rect -7766 302294 -7146 302378
rect -7766 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 -7146 302294
rect -7766 266614 -7146 302058
rect -7766 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 -7146 266614
rect -7766 266294 -7146 266378
rect -7766 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 -7146 266294
rect -7766 230614 -7146 266058
rect -7766 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 -7146 230614
rect -7766 230294 -7146 230378
rect -7766 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 -7146 230294
rect -7766 194614 -7146 230058
rect -7766 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 -7146 194614
rect -7766 194294 -7146 194378
rect -7766 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 -7146 194294
rect -7766 158614 -7146 194058
rect -7766 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 -7146 158614
rect -7766 158294 -7146 158378
rect -7766 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 -7146 158294
rect -7766 122614 -7146 158058
rect -7766 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 -7146 122614
rect -7766 122294 -7146 122378
rect -7766 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 -7146 122294
rect -7766 86614 -7146 122058
rect -7766 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 -7146 86614
rect -7766 86294 -7146 86378
rect -7766 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 -7146 86294
rect -7766 50614 -7146 86058
rect -7766 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 -7146 50614
rect -7766 50294 -7146 50378
rect -7766 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 -7146 50294
rect -7766 14614 -7146 50058
rect -7766 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 -7146 14614
rect -7766 14294 -7146 14378
rect -7766 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 -7146 14294
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 676894 -6186 709082
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 -6186 676894
rect -6806 676574 -6186 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 -6186 676574
rect -6806 640894 -6186 676338
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 -6186 640894
rect -6806 640574 -6186 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 -6186 640574
rect -6806 604894 -6186 640338
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 -6186 604894
rect -6806 604574 -6186 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 -6186 604574
rect -6806 568894 -6186 604338
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 -6186 568894
rect -6806 568574 -6186 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 -6186 568574
rect -6806 532894 -6186 568338
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 -6186 532894
rect -6806 532574 -6186 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 -6186 532574
rect -6806 496894 -6186 532338
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 -6186 496894
rect -6806 496574 -6186 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 -6186 496574
rect -6806 460894 -6186 496338
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 -6186 460894
rect -6806 460574 -6186 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 -6186 460574
rect -6806 424894 -6186 460338
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 -6186 424894
rect -6806 424574 -6186 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 -6186 424574
rect -6806 388894 -6186 424338
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 -6186 388894
rect -6806 388574 -6186 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 -6186 388574
rect -6806 352894 -6186 388338
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 -6186 352894
rect -6806 352574 -6186 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 -6186 352574
rect -6806 316894 -6186 352338
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 -6186 316894
rect -6806 316574 -6186 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 -6186 316574
rect -6806 280894 -6186 316338
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 -6186 280894
rect -6806 280574 -6186 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 -6186 280574
rect -6806 244894 -6186 280338
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 -6186 244894
rect -6806 244574 -6186 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 -6186 244574
rect -6806 208894 -6186 244338
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 -6186 208894
rect -6806 208574 -6186 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 -6186 208574
rect -6806 172894 -6186 208338
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 -6186 172894
rect -6806 172574 -6186 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 -6186 172574
rect -6806 136894 -6186 172338
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 -6186 136894
rect -6806 136574 -6186 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 -6186 136574
rect -6806 100894 -6186 136338
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 -6186 100894
rect -6806 100574 -6186 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 -6186 100574
rect -6806 64894 -6186 100338
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 -6186 64894
rect -6806 64574 -6186 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 -6186 64574
rect -6806 28894 -6186 64338
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 -6186 28894
rect -6806 28574 -6186 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 -6186 28574
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 9854 708678
rect 9234 708358 9854 708442
rect 9234 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 9854 708358
rect -5846 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 -5226 694894
rect -5846 694574 -5226 694658
rect -5846 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 -5226 694574
rect -5846 658894 -5226 694338
rect -5846 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 -5226 658894
rect -5846 658574 -5226 658658
rect -5846 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 -5226 658574
rect -5846 622894 -5226 658338
rect -5846 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 -5226 622894
rect -5846 622574 -5226 622658
rect -5846 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 -5226 622574
rect -5846 586894 -5226 622338
rect -5846 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 -5226 586894
rect -5846 586574 -5226 586658
rect -5846 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 -5226 586574
rect -5846 550894 -5226 586338
rect -5846 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 -5226 550894
rect -5846 550574 -5226 550658
rect -5846 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 -5226 550574
rect -5846 514894 -5226 550338
rect -5846 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 -5226 514894
rect -5846 514574 -5226 514658
rect -5846 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 -5226 514574
rect -5846 478894 -5226 514338
rect -5846 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 -5226 478894
rect -5846 478574 -5226 478658
rect -5846 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 -5226 478574
rect -5846 442894 -5226 478338
rect -5846 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 -5226 442894
rect -5846 442574 -5226 442658
rect -5846 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 -5226 442574
rect -5846 406894 -5226 442338
rect -5846 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 -5226 406894
rect -5846 406574 -5226 406658
rect -5846 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 -5226 406574
rect -5846 370894 -5226 406338
rect -5846 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 -5226 370894
rect -5846 370574 -5226 370658
rect -5846 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 -5226 370574
rect -5846 334894 -5226 370338
rect -5846 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 -5226 334894
rect -5846 334574 -5226 334658
rect -5846 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 -5226 334574
rect -5846 298894 -5226 334338
rect -5846 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 -5226 298894
rect -5846 298574 -5226 298658
rect -5846 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 -5226 298574
rect -5846 262894 -5226 298338
rect -5846 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 -5226 262894
rect -5846 262574 -5226 262658
rect -5846 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 -5226 262574
rect -5846 226894 -5226 262338
rect -5846 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 -5226 226894
rect -5846 226574 -5226 226658
rect -5846 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 -5226 226574
rect -5846 190894 -5226 226338
rect -5846 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 -5226 190894
rect -5846 190574 -5226 190658
rect -5846 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 -5226 190574
rect -5846 154894 -5226 190338
rect -5846 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 -5226 154894
rect -5846 154574 -5226 154658
rect -5846 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 -5226 154574
rect -5846 118894 -5226 154338
rect -5846 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 -5226 118894
rect -5846 118574 -5226 118658
rect -5846 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 -5226 118574
rect -5846 82894 -5226 118338
rect -5846 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 -5226 82894
rect -5846 82574 -5226 82658
rect -5846 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 -5226 82574
rect -5846 46894 -5226 82338
rect -5846 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 -5226 46894
rect -5846 46574 -5226 46658
rect -5846 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 -5226 46574
rect -5846 10894 -5226 46338
rect -5846 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 -5226 10894
rect -5846 10574 -5226 10658
rect -5846 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 -5226 10574
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 673174 -4266 707162
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 -4266 673174
rect -4886 672854 -4266 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 -4266 672854
rect -4886 637174 -4266 672618
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 -4266 637174
rect -4886 636854 -4266 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 -4266 636854
rect -4886 601174 -4266 636618
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 -4266 601174
rect -4886 600854 -4266 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 -4266 600854
rect -4886 565174 -4266 600618
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 -4266 565174
rect -4886 564854 -4266 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 -4266 564854
rect -4886 529174 -4266 564618
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 -4266 529174
rect -4886 528854 -4266 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 -4266 528854
rect -4886 493174 -4266 528618
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 -4266 493174
rect -4886 492854 -4266 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 -4266 492854
rect -4886 457174 -4266 492618
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 -4266 457174
rect -4886 456854 -4266 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 -4266 456854
rect -4886 421174 -4266 456618
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 -4266 421174
rect -4886 420854 -4266 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 -4266 420854
rect -4886 385174 -4266 420618
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 -4266 385174
rect -4886 384854 -4266 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 -4266 384854
rect -4886 349174 -4266 384618
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 -4266 349174
rect -4886 348854 -4266 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 -4266 348854
rect -4886 313174 -4266 348618
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 -4266 313174
rect -4886 312854 -4266 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 -4266 312854
rect -4886 277174 -4266 312618
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 -4266 277174
rect -4886 276854 -4266 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 -4266 276854
rect -4886 241174 -4266 276618
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 -4266 241174
rect -4886 240854 -4266 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 -4266 240854
rect -4886 205174 -4266 240618
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 -4266 205174
rect -4886 204854 -4266 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 -4266 204854
rect -4886 169174 -4266 204618
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 -4266 169174
rect -4886 168854 -4266 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 -4266 168854
rect -4886 133174 -4266 168618
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 -4266 133174
rect -4886 132854 -4266 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 -4266 132854
rect -4886 97174 -4266 132618
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 -4266 97174
rect -4886 96854 -4266 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 -4266 96854
rect -4886 61174 -4266 96618
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 -4266 61174
rect -4886 60854 -4266 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 -4266 60854
rect -4886 25174 -4266 60618
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 -4266 25174
rect -4886 24854 -4266 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 -4266 24854
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 6134 706758
rect 5514 706438 6134 706522
rect 5514 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 6134 706438
rect -3926 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 -3306 691174
rect -3926 690854 -3306 690938
rect -3926 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 -3306 690854
rect -3926 655174 -3306 690618
rect -3926 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 -3306 655174
rect -3926 654854 -3306 654938
rect -3926 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 -3306 654854
rect -3926 619174 -3306 654618
rect -3926 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 -3306 619174
rect -3926 618854 -3306 618938
rect -3926 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 -3306 618854
rect -3926 583174 -3306 618618
rect -3926 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 -3306 583174
rect -3926 582854 -3306 582938
rect -3926 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 -3306 582854
rect -3926 547174 -3306 582618
rect -3926 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 -3306 547174
rect -3926 546854 -3306 546938
rect -3926 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 -3306 546854
rect -3926 511174 -3306 546618
rect -3926 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 -3306 511174
rect -3926 510854 -3306 510938
rect -3926 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 -3306 510854
rect -3926 475174 -3306 510618
rect -3926 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 -3306 475174
rect -3926 474854 -3306 474938
rect -3926 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 -3306 474854
rect -3926 439174 -3306 474618
rect -3926 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 -3306 439174
rect -3926 438854 -3306 438938
rect -3926 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 -3306 438854
rect -3926 403174 -3306 438618
rect -3926 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 -3306 403174
rect -3926 402854 -3306 402938
rect -3926 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 -3306 402854
rect -3926 367174 -3306 402618
rect -3926 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 -3306 367174
rect -3926 366854 -3306 366938
rect -3926 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 -3306 366854
rect -3926 331174 -3306 366618
rect -3926 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 -3306 331174
rect -3926 330854 -3306 330938
rect -3926 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 -3306 330854
rect -3926 295174 -3306 330618
rect -3926 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 -3306 295174
rect -3926 294854 -3306 294938
rect -3926 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 -3306 294854
rect -3926 259174 -3306 294618
rect -3926 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 -3306 259174
rect -3926 258854 -3306 258938
rect -3926 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 -3306 258854
rect -3926 223174 -3306 258618
rect -3926 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 -3306 223174
rect -3926 222854 -3306 222938
rect -3926 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 -3306 222854
rect -3926 187174 -3306 222618
rect -3926 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 -3306 187174
rect -3926 186854 -3306 186938
rect -3926 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 -3306 186854
rect -3926 151174 -3306 186618
rect -3926 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 -3306 151174
rect -3926 150854 -3306 150938
rect -3926 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 -3306 150854
rect -3926 115174 -3306 150618
rect -3926 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 -3306 115174
rect -3926 114854 -3306 114938
rect -3926 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 -3306 114854
rect -3926 79174 -3306 114618
rect -3926 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 -3306 79174
rect -3926 78854 -3306 78938
rect -3926 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 -3306 78854
rect -3926 43174 -3306 78618
rect -3926 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 -3306 43174
rect -3926 42854 -3306 42938
rect -3926 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 -3306 42854
rect -3926 7174 -3306 42618
rect -3926 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 -3306 7174
rect -3926 6854 -3306 6938
rect -3926 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 -3306 6854
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 702000 2414 704282
rect 5514 702000 6134 706202
rect 9234 702000 9854 708122
rect 12954 702000 13574 710042
rect 30954 711558 31574 711590
rect 30954 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 31574 711558
rect 30954 711238 31574 711322
rect 30954 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 31574 711238
rect 27234 709638 27854 709670
rect 27234 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 27854 709638
rect 27234 709318 27854 709402
rect 27234 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 27854 709318
rect 23514 707718 24134 707750
rect 23514 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 24134 707718
rect 23514 707398 24134 707482
rect 23514 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 24134 707398
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 19794 702000 20414 705242
rect 23514 702000 24134 707162
rect 27234 702000 27854 709082
rect 30954 702000 31574 711002
rect 48954 710598 49574 711590
rect 48954 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 49574 710598
rect 48954 710278 49574 710362
rect 48954 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 49574 710278
rect 45234 708678 45854 709670
rect 45234 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 45854 708678
rect 45234 708358 45854 708442
rect 45234 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 45854 708358
rect 41514 706758 42134 707750
rect 41514 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 42134 706758
rect 41514 706438 42134 706522
rect 41514 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 42134 706438
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 702000 38414 704282
rect 41514 702000 42134 706202
rect 45234 702000 45854 708122
rect 48954 702000 49574 710042
rect 66954 711558 67574 711590
rect 66954 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 67574 711558
rect 66954 711238 67574 711322
rect 66954 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 67574 711238
rect 63234 709638 63854 709670
rect 63234 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 63854 709638
rect 63234 709318 63854 709402
rect 63234 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 63854 709318
rect 59514 707718 60134 707750
rect 59514 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 60134 707718
rect 59514 707398 60134 707482
rect 59514 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 60134 707398
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 702000 56414 705242
rect 59514 702000 60134 707162
rect 63234 702000 63854 709082
rect 66954 702000 67574 711002
rect 84954 710598 85574 711590
rect 84954 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 85574 710598
rect 84954 710278 85574 710362
rect 84954 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 85574 710278
rect 81234 708678 81854 709670
rect 81234 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 81854 708678
rect 81234 708358 81854 708442
rect 81234 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 81854 708358
rect 77514 706758 78134 707750
rect 77514 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 78134 706758
rect 77514 706438 78134 706522
rect 77514 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 78134 706438
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 702000 74414 704282
rect 77514 702000 78134 706202
rect 81234 702000 81854 708122
rect 84954 702000 85574 710042
rect 102954 711558 103574 711590
rect 102954 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 103574 711558
rect 102954 711238 103574 711322
rect 102954 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 103574 711238
rect 99234 709638 99854 709670
rect 99234 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 99854 709638
rect 99234 709318 99854 709402
rect 99234 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 99854 709318
rect 95514 707718 96134 707750
rect 95514 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 96134 707718
rect 95514 707398 96134 707482
rect 95514 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 96134 707398
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 702000 92414 705242
rect 95514 702000 96134 707162
rect 99234 702000 99854 709082
rect 102954 702000 103574 711002
rect 120954 710598 121574 711590
rect 120954 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 121574 710598
rect 120954 710278 121574 710362
rect 120954 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 121574 710278
rect 117234 708678 117854 709670
rect 117234 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 117854 708678
rect 117234 708358 117854 708442
rect 117234 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 117854 708358
rect 113514 706758 114134 707750
rect 113514 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 114134 706758
rect 113514 706438 114134 706522
rect 113514 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 114134 706438
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 702000 110414 704282
rect 113514 702000 114134 706202
rect 117234 702000 117854 708122
rect 120954 702000 121574 710042
rect 138954 711558 139574 711590
rect 138954 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 139574 711558
rect 138954 711238 139574 711322
rect 138954 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 139574 711238
rect 135234 709638 135854 709670
rect 135234 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 135854 709638
rect 135234 709318 135854 709402
rect 135234 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 135854 709318
rect 131514 707718 132134 707750
rect 131514 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 132134 707718
rect 131514 707398 132134 707482
rect 131514 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 132134 707398
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 127794 702000 128414 705242
rect 131514 702000 132134 707162
rect 135234 702000 135854 709082
rect 138954 702000 139574 711002
rect 156954 710598 157574 711590
rect 156954 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 157574 710598
rect 156954 710278 157574 710362
rect 156954 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 157574 710278
rect 153234 708678 153854 709670
rect 153234 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 153854 708678
rect 153234 708358 153854 708442
rect 153234 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 153854 708358
rect 149514 706758 150134 707750
rect 149514 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 150134 706758
rect 149514 706438 150134 706522
rect 149514 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 150134 706438
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 702000 146414 704282
rect 149514 702000 150134 706202
rect 153234 702000 153854 708122
rect 156954 702000 157574 710042
rect 174954 711558 175574 711590
rect 174954 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 175574 711558
rect 174954 711238 175574 711322
rect 174954 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 175574 711238
rect 171234 709638 171854 709670
rect 171234 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 171854 709638
rect 171234 709318 171854 709402
rect 171234 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 171854 709318
rect 167514 707718 168134 707750
rect 167514 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 168134 707718
rect 167514 707398 168134 707482
rect 167514 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 168134 707398
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 702000 164414 705242
rect 167514 702000 168134 707162
rect 171234 702000 171854 709082
rect 174954 702000 175574 711002
rect 192954 710598 193574 711590
rect 192954 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 193574 710598
rect 192954 710278 193574 710362
rect 192954 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 193574 710278
rect 189234 708678 189854 709670
rect 189234 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 189854 708678
rect 189234 708358 189854 708442
rect 189234 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 189854 708358
rect 185514 706758 186134 707750
rect 185514 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 186134 706758
rect 185514 706438 186134 706522
rect 185514 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 186134 706438
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 702000 182414 704282
rect 185514 702000 186134 706202
rect 189234 702000 189854 708122
rect 192954 702000 193574 710042
rect 210954 711558 211574 711590
rect 210954 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 211574 711558
rect 210954 711238 211574 711322
rect 210954 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 211574 711238
rect 207234 709638 207854 709670
rect 207234 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 207854 709638
rect 207234 709318 207854 709402
rect 207234 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 207854 709318
rect 203514 707718 204134 707750
rect 203514 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 204134 707718
rect 203514 707398 204134 707482
rect 203514 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 204134 707398
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 702000 200414 705242
rect 203514 702000 204134 707162
rect 207234 702000 207854 709082
rect 210954 702000 211574 711002
rect 228954 710598 229574 711590
rect 228954 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 229574 710598
rect 228954 710278 229574 710362
rect 228954 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 229574 710278
rect 225234 708678 225854 709670
rect 225234 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 225854 708678
rect 225234 708358 225854 708442
rect 225234 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 225854 708358
rect 221514 706758 222134 707750
rect 221514 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 222134 706758
rect 221514 706438 222134 706522
rect 221514 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 222134 706438
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 702000 218414 704282
rect 221514 702000 222134 706202
rect 225234 702000 225854 708122
rect 228954 702000 229574 710042
rect 246954 711558 247574 711590
rect 246954 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 247574 711558
rect 246954 711238 247574 711322
rect 246954 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 247574 711238
rect 243234 709638 243854 709670
rect 243234 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 243854 709638
rect 243234 709318 243854 709402
rect 243234 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 243854 709318
rect 239514 707718 240134 707750
rect 239514 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 240134 707718
rect 239514 707398 240134 707482
rect 239514 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 240134 707398
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 235794 702000 236414 705242
rect 239514 702000 240134 707162
rect 243234 702000 243854 709082
rect 246954 702000 247574 711002
rect 264954 710598 265574 711590
rect 264954 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 265574 710598
rect 264954 710278 265574 710362
rect 264954 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 265574 710278
rect 261234 708678 261854 709670
rect 261234 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 261854 708678
rect 261234 708358 261854 708442
rect 261234 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 261854 708358
rect 257514 706758 258134 707750
rect 257514 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 258134 706758
rect 257514 706438 258134 706522
rect 257514 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 258134 706438
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 702000 254414 704282
rect 257514 702000 258134 706202
rect 261234 702000 261854 708122
rect 264954 702000 265574 710042
rect 282954 711558 283574 711590
rect 282954 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 283574 711558
rect 282954 711238 283574 711322
rect 282954 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 283574 711238
rect 279234 709638 279854 709670
rect 279234 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 279854 709638
rect 279234 709318 279854 709402
rect 279234 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 279854 709318
rect 275514 707718 276134 707750
rect 275514 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 276134 707718
rect 275514 707398 276134 707482
rect 275514 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 276134 707398
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 271794 702000 272414 705242
rect 275514 702000 276134 707162
rect 279234 702000 279854 709082
rect 282954 702000 283574 711002
rect 300954 710598 301574 711590
rect 300954 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 301574 710598
rect 300954 710278 301574 710362
rect 300954 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 301574 710278
rect 297234 708678 297854 709670
rect 297234 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 297854 708678
rect 297234 708358 297854 708442
rect 297234 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 297854 708358
rect 293514 706758 294134 707750
rect 293514 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 294134 706758
rect 293514 706438 294134 706522
rect 293514 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 294134 706438
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 702000 290414 704282
rect 293514 702000 294134 706202
rect 297234 702000 297854 708122
rect 300954 702000 301574 710042
rect 318954 711558 319574 711590
rect 318954 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 319574 711558
rect 318954 711238 319574 711322
rect 318954 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 319574 711238
rect 315234 709638 315854 709670
rect 315234 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 315854 709638
rect 315234 709318 315854 709402
rect 315234 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 315854 709318
rect 311514 707718 312134 707750
rect 311514 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 312134 707718
rect 311514 707398 312134 707482
rect 311514 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 312134 707398
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 702000 308414 705242
rect 311514 702000 312134 707162
rect 315234 702000 315854 709082
rect 318954 702000 319574 711002
rect 336954 710598 337574 711590
rect 336954 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 337574 710598
rect 336954 710278 337574 710362
rect 336954 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 337574 710278
rect 333234 708678 333854 709670
rect 333234 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 333854 708678
rect 333234 708358 333854 708442
rect 333234 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 333854 708358
rect 329514 706758 330134 707750
rect 329514 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 330134 706758
rect 329514 706438 330134 706522
rect 329514 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 330134 706438
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 702000 326414 704282
rect 329514 702000 330134 706202
rect 333234 702000 333854 708122
rect 336954 702000 337574 710042
rect 354954 711558 355574 711590
rect 354954 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 355574 711558
rect 354954 711238 355574 711322
rect 354954 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 355574 711238
rect 351234 709638 351854 709670
rect 351234 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 351854 709638
rect 351234 709318 351854 709402
rect 351234 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 351854 709318
rect 347514 707718 348134 707750
rect 347514 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 348134 707718
rect 347514 707398 348134 707482
rect 347514 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 348134 707398
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 343794 702000 344414 705242
rect 347514 702000 348134 707162
rect 351234 702000 351854 709082
rect 354954 702000 355574 711002
rect 372954 710598 373574 711590
rect 372954 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 373574 710598
rect 372954 710278 373574 710362
rect 372954 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 373574 710278
rect 369234 708678 369854 709670
rect 369234 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 369854 708678
rect 369234 708358 369854 708442
rect 369234 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 369854 708358
rect 365514 706758 366134 707750
rect 365514 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 366134 706758
rect 365514 706438 366134 706522
rect 365514 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 366134 706438
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 702000 362414 704282
rect 365514 702000 366134 706202
rect 369234 702000 369854 708122
rect 372954 702000 373574 710042
rect 390954 711558 391574 711590
rect 390954 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 391574 711558
rect 390954 711238 391574 711322
rect 390954 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 391574 711238
rect 387234 709638 387854 709670
rect 387234 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 387854 709638
rect 387234 709318 387854 709402
rect 387234 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 387854 709318
rect 383514 707718 384134 707750
rect 383514 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 384134 707718
rect 383514 707398 384134 707482
rect 383514 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 384134 707398
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 379794 702000 380414 705242
rect 383514 702000 384134 707162
rect 386275 702268 386341 702269
rect 386275 702204 386276 702268
rect 386340 702204 386341 702268
rect 386275 702203 386341 702204
rect 259131 701180 259197 701181
rect 259131 701116 259132 701180
rect 259196 701116 259197 701180
rect 259131 701115 259197 701116
rect 13859 699412 13925 699413
rect 13859 699348 13860 699412
rect 13924 699348 13925 699412
rect 13859 699347 13925 699348
rect 95187 699412 95253 699413
rect 95187 699348 95188 699412
rect 95252 699348 95253 699412
rect 95187 699347 95253 699348
rect 13862 698325 13922 699347
rect 13859 698324 13925 698325
rect 13859 698260 13860 698324
rect 13924 698260 13925 698324
rect 13859 698259 13925 698260
rect 95190 697781 95250 699347
rect 259134 699141 259194 701115
rect 386278 699549 386338 702203
rect 387234 702000 387854 709082
rect 390954 702000 391574 711002
rect 408954 710598 409574 711590
rect 408954 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 409574 710598
rect 408954 710278 409574 710362
rect 408954 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 409574 710278
rect 405234 708678 405854 709670
rect 405234 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 405854 708678
rect 405234 708358 405854 708442
rect 405234 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 405854 708358
rect 401514 706758 402134 707750
rect 401514 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 402134 706758
rect 401514 706438 402134 706522
rect 401514 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 402134 706438
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 702000 398414 704282
rect 401514 702000 402134 706202
rect 405234 702000 405854 708122
rect 408954 702000 409574 710042
rect 426954 711558 427574 711590
rect 426954 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 427574 711558
rect 426954 711238 427574 711322
rect 426954 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 427574 711238
rect 423234 709638 423854 709670
rect 423234 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 423854 709638
rect 423234 709318 423854 709402
rect 423234 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 423854 709318
rect 419514 707718 420134 707750
rect 419514 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 420134 707718
rect 419514 707398 420134 707482
rect 419514 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 420134 707398
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 415794 702000 416414 705242
rect 419514 702000 420134 707162
rect 423234 702000 423854 709082
rect 426954 702000 427574 711002
rect 444954 710598 445574 711590
rect 444954 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 445574 710598
rect 444954 710278 445574 710362
rect 444954 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 445574 710278
rect 441234 708678 441854 709670
rect 441234 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 441854 708678
rect 441234 708358 441854 708442
rect 441234 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 441854 708358
rect 437514 706758 438134 707750
rect 437514 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 438134 706758
rect 437514 706438 438134 706522
rect 437514 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 438134 706438
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 702000 434414 704282
rect 437514 702000 438134 706202
rect 441234 702000 441854 708122
rect 444954 702000 445574 710042
rect 462954 711558 463574 711590
rect 462954 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 463574 711558
rect 462954 711238 463574 711322
rect 462954 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 463574 711238
rect 459234 709638 459854 709670
rect 459234 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 459854 709638
rect 459234 709318 459854 709402
rect 459234 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 459854 709318
rect 455514 707718 456134 707750
rect 455514 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 456134 707718
rect 455514 707398 456134 707482
rect 455514 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 456134 707398
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 702000 452414 705242
rect 455514 702000 456134 707162
rect 459234 702000 459854 709082
rect 462954 702000 463574 711002
rect 480954 710598 481574 711590
rect 480954 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 481574 710598
rect 480954 710278 481574 710362
rect 480954 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 481574 710278
rect 477234 708678 477854 709670
rect 477234 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 477854 708678
rect 477234 708358 477854 708442
rect 477234 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 477854 708358
rect 473514 706758 474134 707750
rect 473514 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 474134 706758
rect 473514 706438 474134 706522
rect 473514 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 474134 706438
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 702000 470414 704282
rect 473514 702000 474134 706202
rect 477234 702000 477854 708122
rect 480954 702000 481574 710042
rect 498954 711558 499574 711590
rect 498954 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 499574 711558
rect 498954 711238 499574 711322
rect 498954 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 499574 711238
rect 495234 709638 495854 709670
rect 495234 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 495854 709638
rect 495234 709318 495854 709402
rect 495234 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 495854 709318
rect 491514 707718 492134 707750
rect 491514 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 492134 707718
rect 491514 707398 492134 707482
rect 491514 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 492134 707398
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 487794 702000 488414 705242
rect 491514 702000 492134 707162
rect 495234 702000 495854 709082
rect 498954 702000 499574 711002
rect 516954 710598 517574 711590
rect 516954 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 517574 710598
rect 516954 710278 517574 710362
rect 516954 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 517574 710278
rect 513234 708678 513854 709670
rect 513234 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 513854 708678
rect 513234 708358 513854 708442
rect 513234 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 513854 708358
rect 509514 706758 510134 707750
rect 509514 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 510134 706758
rect 509514 706438 510134 706522
rect 509514 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 510134 706438
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 702000 506414 704282
rect 509514 702000 510134 706202
rect 513234 702000 513854 708122
rect 516954 702000 517574 710042
rect 534954 711558 535574 711590
rect 534954 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 535574 711558
rect 534954 711238 535574 711322
rect 534954 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 535574 711238
rect 531234 709638 531854 709670
rect 531234 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 531854 709638
rect 531234 709318 531854 709402
rect 531234 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 531854 709318
rect 527514 707718 528134 707750
rect 527514 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 528134 707718
rect 527514 707398 528134 707482
rect 527514 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 528134 707398
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 702000 524414 705242
rect 527514 702000 528134 707162
rect 531234 702000 531854 709082
rect 534954 702000 535574 711002
rect 552954 710598 553574 711590
rect 552954 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 553574 710598
rect 552954 710278 553574 710362
rect 552954 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 553574 710278
rect 549234 708678 549854 709670
rect 549234 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 549854 708678
rect 549234 708358 549854 708442
rect 549234 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 549854 708358
rect 545514 706758 546134 707750
rect 545514 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 546134 706758
rect 545514 706438 546134 706522
rect 545514 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 546134 706438
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 702000 542414 704282
rect 545514 702000 546134 706202
rect 549234 702000 549854 708122
rect 552954 702000 553574 710042
rect 570954 711558 571574 711590
rect 570954 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 571574 711558
rect 570954 711238 571574 711322
rect 570954 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 571574 711238
rect 567234 709638 567854 709670
rect 567234 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 567854 709638
rect 567234 709318 567854 709402
rect 567234 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 567854 709318
rect 563514 707718 564134 707750
rect 563514 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 564134 707718
rect 563514 707398 564134 707482
rect 563514 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 564134 707398
rect 559794 705798 560414 705830
rect 559794 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 560414 705798
rect 559794 705478 560414 705562
rect 559794 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 560414 705478
rect 559794 702000 560414 705242
rect 563514 702000 564134 707162
rect 386275 699548 386341 699549
rect 386275 699484 386276 699548
rect 386340 699484 386341 699548
rect 386275 699483 386341 699484
rect 418659 699412 418725 699413
rect 418659 699348 418660 699412
rect 418724 699348 418725 699412
rect 418659 699347 418725 699348
rect 433379 699412 433445 699413
rect 433379 699348 433380 699412
rect 433444 699348 433445 699412
rect 433379 699347 433445 699348
rect 462819 699412 462885 699413
rect 462819 699348 462820 699412
rect 462884 699348 462885 699412
rect 462819 699347 462885 699348
rect 492627 699412 492693 699413
rect 492627 699348 492628 699412
rect 492692 699348 492693 699412
rect 492627 699347 492693 699348
rect 539915 699412 539981 699413
rect 539915 699348 539916 699412
rect 539980 699348 539981 699412
rect 539915 699347 539981 699348
rect 259131 699140 259197 699141
rect 259131 699076 259132 699140
rect 259196 699076 259197 699140
rect 259131 699075 259197 699076
rect 418662 698053 418722 699347
rect 418843 699276 418909 699277
rect 418843 699212 418844 699276
rect 418908 699212 418909 699276
rect 418843 699211 418909 699212
rect 418846 698053 418906 699211
rect 433382 698189 433442 699347
rect 433379 698188 433445 698189
rect 433379 698124 433380 698188
rect 433444 698124 433445 698188
rect 433379 698123 433445 698124
rect 418659 698052 418725 698053
rect 418659 697988 418660 698052
rect 418724 697988 418725 698052
rect 418659 697987 418725 697988
rect 418843 698052 418909 698053
rect 418843 697988 418844 698052
rect 418908 697988 418909 698052
rect 418843 697987 418909 697988
rect 462822 697917 462882 699347
rect 462819 697916 462885 697917
rect 462819 697852 462820 697916
rect 462884 697852 462885 697916
rect 462819 697851 462885 697852
rect 95187 697780 95253 697781
rect 95187 697716 95188 697780
rect 95252 697716 95253 697780
rect 95187 697715 95253 697716
rect 492630 697645 492690 699347
rect 539918 698461 539978 699347
rect 539915 698460 539981 698461
rect 539915 698396 539916 698460
rect 539980 698396 539981 698460
rect 539915 698395 539981 698396
rect 492627 697644 492693 697645
rect 492627 697580 492628 697644
rect 492692 697580 492693 697644
rect 492627 697579 492693 697580
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect 8208 687454 8528 687486
rect 8208 687218 8250 687454
rect 8486 687218 8528 687454
rect 8208 687134 8528 687218
rect 8208 686898 8250 687134
rect 8486 686898 8528 687134
rect 8208 686866 8528 686898
rect 38928 687454 39248 687486
rect 38928 687218 38970 687454
rect 39206 687218 39248 687454
rect 38928 687134 39248 687218
rect 38928 686898 38970 687134
rect 39206 686898 39248 687134
rect 38928 686866 39248 686898
rect 69648 687454 69968 687486
rect 69648 687218 69690 687454
rect 69926 687218 69968 687454
rect 69648 687134 69968 687218
rect 69648 686898 69690 687134
rect 69926 686898 69968 687134
rect 69648 686866 69968 686898
rect 100368 687454 100688 687486
rect 100368 687218 100410 687454
rect 100646 687218 100688 687454
rect 100368 687134 100688 687218
rect 100368 686898 100410 687134
rect 100646 686898 100688 687134
rect 100368 686866 100688 686898
rect 131088 687454 131408 687486
rect 131088 687218 131130 687454
rect 131366 687218 131408 687454
rect 131088 687134 131408 687218
rect 131088 686898 131130 687134
rect 131366 686898 131408 687134
rect 131088 686866 131408 686898
rect 161808 687454 162128 687486
rect 161808 687218 161850 687454
rect 162086 687218 162128 687454
rect 161808 687134 162128 687218
rect 161808 686898 161850 687134
rect 162086 686898 162128 687134
rect 161808 686866 162128 686898
rect 192528 687454 192848 687486
rect 192528 687218 192570 687454
rect 192806 687218 192848 687454
rect 192528 687134 192848 687218
rect 192528 686898 192570 687134
rect 192806 686898 192848 687134
rect 192528 686866 192848 686898
rect 223248 687454 223568 687486
rect 223248 687218 223290 687454
rect 223526 687218 223568 687454
rect 223248 687134 223568 687218
rect 223248 686898 223290 687134
rect 223526 686898 223568 687134
rect 223248 686866 223568 686898
rect 253968 687454 254288 687486
rect 253968 687218 254010 687454
rect 254246 687218 254288 687454
rect 253968 687134 254288 687218
rect 253968 686898 254010 687134
rect 254246 686898 254288 687134
rect 253968 686866 254288 686898
rect 284688 687454 285008 687486
rect 284688 687218 284730 687454
rect 284966 687218 285008 687454
rect 284688 687134 285008 687218
rect 284688 686898 284730 687134
rect 284966 686898 285008 687134
rect 284688 686866 285008 686898
rect 315408 687454 315728 687486
rect 315408 687218 315450 687454
rect 315686 687218 315728 687454
rect 315408 687134 315728 687218
rect 315408 686898 315450 687134
rect 315686 686898 315728 687134
rect 315408 686866 315728 686898
rect 346128 687454 346448 687486
rect 346128 687218 346170 687454
rect 346406 687218 346448 687454
rect 346128 687134 346448 687218
rect 346128 686898 346170 687134
rect 346406 686898 346448 687134
rect 346128 686866 346448 686898
rect 376848 687454 377168 687486
rect 376848 687218 376890 687454
rect 377126 687218 377168 687454
rect 376848 687134 377168 687218
rect 376848 686898 376890 687134
rect 377126 686898 377168 687134
rect 376848 686866 377168 686898
rect 407568 687454 407888 687486
rect 407568 687218 407610 687454
rect 407846 687218 407888 687454
rect 407568 687134 407888 687218
rect 407568 686898 407610 687134
rect 407846 686898 407888 687134
rect 407568 686866 407888 686898
rect 438288 687454 438608 687486
rect 438288 687218 438330 687454
rect 438566 687218 438608 687454
rect 438288 687134 438608 687218
rect 438288 686898 438330 687134
rect 438566 686898 438608 687134
rect 438288 686866 438608 686898
rect 469008 687454 469328 687486
rect 469008 687218 469050 687454
rect 469286 687218 469328 687454
rect 469008 687134 469328 687218
rect 469008 686898 469050 687134
rect 469286 686898 469328 687134
rect 469008 686866 469328 686898
rect 499728 687454 500048 687486
rect 499728 687218 499770 687454
rect 500006 687218 500048 687454
rect 499728 687134 500048 687218
rect 499728 686898 499770 687134
rect 500006 686898 500048 687134
rect 499728 686866 500048 686898
rect 530448 687454 530768 687486
rect 530448 687218 530490 687454
rect 530726 687218 530768 687454
rect 530448 687134 530768 687218
rect 530448 686898 530490 687134
rect 530726 686898 530768 687134
rect 530448 686866 530768 686898
rect 561168 687454 561488 687486
rect 561168 687218 561210 687454
rect 561446 687218 561488 687454
rect 561168 687134 561488 687218
rect 561168 686898 561210 687134
rect 561446 686898 561488 687134
rect 561168 686866 561488 686898
rect 567234 676894 567854 709082
rect 567234 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 567854 676894
rect 567234 676574 567854 676658
rect 567234 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 567854 676574
rect 23568 669454 23888 669486
rect 23568 669218 23610 669454
rect 23846 669218 23888 669454
rect 23568 669134 23888 669218
rect 23568 668898 23610 669134
rect 23846 668898 23888 669134
rect 23568 668866 23888 668898
rect 54288 669454 54608 669486
rect 54288 669218 54330 669454
rect 54566 669218 54608 669454
rect 54288 669134 54608 669218
rect 54288 668898 54330 669134
rect 54566 668898 54608 669134
rect 54288 668866 54608 668898
rect 85008 669454 85328 669486
rect 85008 669218 85050 669454
rect 85286 669218 85328 669454
rect 85008 669134 85328 669218
rect 85008 668898 85050 669134
rect 85286 668898 85328 669134
rect 85008 668866 85328 668898
rect 115728 669454 116048 669486
rect 115728 669218 115770 669454
rect 116006 669218 116048 669454
rect 115728 669134 116048 669218
rect 115728 668898 115770 669134
rect 116006 668898 116048 669134
rect 115728 668866 116048 668898
rect 146448 669454 146768 669486
rect 146448 669218 146490 669454
rect 146726 669218 146768 669454
rect 146448 669134 146768 669218
rect 146448 668898 146490 669134
rect 146726 668898 146768 669134
rect 146448 668866 146768 668898
rect 177168 669454 177488 669486
rect 177168 669218 177210 669454
rect 177446 669218 177488 669454
rect 177168 669134 177488 669218
rect 177168 668898 177210 669134
rect 177446 668898 177488 669134
rect 177168 668866 177488 668898
rect 207888 669454 208208 669486
rect 207888 669218 207930 669454
rect 208166 669218 208208 669454
rect 207888 669134 208208 669218
rect 207888 668898 207930 669134
rect 208166 668898 208208 669134
rect 207888 668866 208208 668898
rect 238608 669454 238928 669486
rect 238608 669218 238650 669454
rect 238886 669218 238928 669454
rect 238608 669134 238928 669218
rect 238608 668898 238650 669134
rect 238886 668898 238928 669134
rect 238608 668866 238928 668898
rect 269328 669454 269648 669486
rect 269328 669218 269370 669454
rect 269606 669218 269648 669454
rect 269328 669134 269648 669218
rect 269328 668898 269370 669134
rect 269606 668898 269648 669134
rect 269328 668866 269648 668898
rect 300048 669454 300368 669486
rect 300048 669218 300090 669454
rect 300326 669218 300368 669454
rect 300048 669134 300368 669218
rect 300048 668898 300090 669134
rect 300326 668898 300368 669134
rect 300048 668866 300368 668898
rect 330768 669454 331088 669486
rect 330768 669218 330810 669454
rect 331046 669218 331088 669454
rect 330768 669134 331088 669218
rect 330768 668898 330810 669134
rect 331046 668898 331088 669134
rect 330768 668866 331088 668898
rect 361488 669454 361808 669486
rect 361488 669218 361530 669454
rect 361766 669218 361808 669454
rect 361488 669134 361808 669218
rect 361488 668898 361530 669134
rect 361766 668898 361808 669134
rect 361488 668866 361808 668898
rect 392208 669454 392528 669486
rect 392208 669218 392250 669454
rect 392486 669218 392528 669454
rect 392208 669134 392528 669218
rect 392208 668898 392250 669134
rect 392486 668898 392528 669134
rect 392208 668866 392528 668898
rect 422928 669454 423248 669486
rect 422928 669218 422970 669454
rect 423206 669218 423248 669454
rect 422928 669134 423248 669218
rect 422928 668898 422970 669134
rect 423206 668898 423248 669134
rect 422928 668866 423248 668898
rect 453648 669454 453968 669486
rect 453648 669218 453690 669454
rect 453926 669218 453968 669454
rect 453648 669134 453968 669218
rect 453648 668898 453690 669134
rect 453926 668898 453968 669134
rect 453648 668866 453968 668898
rect 484368 669454 484688 669486
rect 484368 669218 484410 669454
rect 484646 669218 484688 669454
rect 484368 669134 484688 669218
rect 484368 668898 484410 669134
rect 484646 668898 484688 669134
rect 484368 668866 484688 668898
rect 515088 669454 515408 669486
rect 515088 669218 515130 669454
rect 515366 669218 515408 669454
rect 515088 669134 515408 669218
rect 515088 668898 515130 669134
rect 515366 668898 515408 669134
rect 515088 668866 515408 668898
rect 545808 669454 546128 669486
rect 545808 669218 545850 669454
rect 546086 669218 546128 669454
rect 545808 669134 546128 669218
rect 545808 668898 545850 669134
rect 546086 668898 546128 669134
rect 545808 668866 546128 668898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect 8208 651454 8528 651486
rect 8208 651218 8250 651454
rect 8486 651218 8528 651454
rect 8208 651134 8528 651218
rect 8208 650898 8250 651134
rect 8486 650898 8528 651134
rect 8208 650866 8528 650898
rect 38928 651454 39248 651486
rect 38928 651218 38970 651454
rect 39206 651218 39248 651454
rect 38928 651134 39248 651218
rect 38928 650898 38970 651134
rect 39206 650898 39248 651134
rect 38928 650866 39248 650898
rect 69648 651454 69968 651486
rect 69648 651218 69690 651454
rect 69926 651218 69968 651454
rect 69648 651134 69968 651218
rect 69648 650898 69690 651134
rect 69926 650898 69968 651134
rect 69648 650866 69968 650898
rect 100368 651454 100688 651486
rect 100368 651218 100410 651454
rect 100646 651218 100688 651454
rect 100368 651134 100688 651218
rect 100368 650898 100410 651134
rect 100646 650898 100688 651134
rect 100368 650866 100688 650898
rect 131088 651454 131408 651486
rect 131088 651218 131130 651454
rect 131366 651218 131408 651454
rect 131088 651134 131408 651218
rect 131088 650898 131130 651134
rect 131366 650898 131408 651134
rect 131088 650866 131408 650898
rect 161808 651454 162128 651486
rect 161808 651218 161850 651454
rect 162086 651218 162128 651454
rect 161808 651134 162128 651218
rect 161808 650898 161850 651134
rect 162086 650898 162128 651134
rect 161808 650866 162128 650898
rect 192528 651454 192848 651486
rect 192528 651218 192570 651454
rect 192806 651218 192848 651454
rect 192528 651134 192848 651218
rect 192528 650898 192570 651134
rect 192806 650898 192848 651134
rect 192528 650866 192848 650898
rect 223248 651454 223568 651486
rect 223248 651218 223290 651454
rect 223526 651218 223568 651454
rect 223248 651134 223568 651218
rect 223248 650898 223290 651134
rect 223526 650898 223568 651134
rect 223248 650866 223568 650898
rect 253968 651454 254288 651486
rect 253968 651218 254010 651454
rect 254246 651218 254288 651454
rect 253968 651134 254288 651218
rect 253968 650898 254010 651134
rect 254246 650898 254288 651134
rect 253968 650866 254288 650898
rect 284688 651454 285008 651486
rect 284688 651218 284730 651454
rect 284966 651218 285008 651454
rect 284688 651134 285008 651218
rect 284688 650898 284730 651134
rect 284966 650898 285008 651134
rect 284688 650866 285008 650898
rect 315408 651454 315728 651486
rect 315408 651218 315450 651454
rect 315686 651218 315728 651454
rect 315408 651134 315728 651218
rect 315408 650898 315450 651134
rect 315686 650898 315728 651134
rect 315408 650866 315728 650898
rect 346128 651454 346448 651486
rect 346128 651218 346170 651454
rect 346406 651218 346448 651454
rect 346128 651134 346448 651218
rect 346128 650898 346170 651134
rect 346406 650898 346448 651134
rect 346128 650866 346448 650898
rect 376848 651454 377168 651486
rect 376848 651218 376890 651454
rect 377126 651218 377168 651454
rect 376848 651134 377168 651218
rect 376848 650898 376890 651134
rect 377126 650898 377168 651134
rect 376848 650866 377168 650898
rect 407568 651454 407888 651486
rect 407568 651218 407610 651454
rect 407846 651218 407888 651454
rect 407568 651134 407888 651218
rect 407568 650898 407610 651134
rect 407846 650898 407888 651134
rect 407568 650866 407888 650898
rect 438288 651454 438608 651486
rect 438288 651218 438330 651454
rect 438566 651218 438608 651454
rect 438288 651134 438608 651218
rect 438288 650898 438330 651134
rect 438566 650898 438608 651134
rect 438288 650866 438608 650898
rect 469008 651454 469328 651486
rect 469008 651218 469050 651454
rect 469286 651218 469328 651454
rect 469008 651134 469328 651218
rect 469008 650898 469050 651134
rect 469286 650898 469328 651134
rect 469008 650866 469328 650898
rect 499728 651454 500048 651486
rect 499728 651218 499770 651454
rect 500006 651218 500048 651454
rect 499728 651134 500048 651218
rect 499728 650898 499770 651134
rect 500006 650898 500048 651134
rect 499728 650866 500048 650898
rect 530448 651454 530768 651486
rect 530448 651218 530490 651454
rect 530726 651218 530768 651454
rect 530448 651134 530768 651218
rect 530448 650898 530490 651134
rect 530726 650898 530768 651134
rect 530448 650866 530768 650898
rect 561168 651454 561488 651486
rect 561168 651218 561210 651454
rect 561446 651218 561488 651454
rect 561168 651134 561488 651218
rect 561168 650898 561210 651134
rect 561446 650898 561488 651134
rect 561168 650866 561488 650898
rect 567234 640894 567854 676338
rect 567234 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 567854 640894
rect 567234 640574 567854 640658
rect 567234 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 567854 640574
rect 23568 633454 23888 633486
rect 23568 633218 23610 633454
rect 23846 633218 23888 633454
rect 23568 633134 23888 633218
rect 23568 632898 23610 633134
rect 23846 632898 23888 633134
rect 23568 632866 23888 632898
rect 54288 633454 54608 633486
rect 54288 633218 54330 633454
rect 54566 633218 54608 633454
rect 54288 633134 54608 633218
rect 54288 632898 54330 633134
rect 54566 632898 54608 633134
rect 54288 632866 54608 632898
rect 85008 633454 85328 633486
rect 85008 633218 85050 633454
rect 85286 633218 85328 633454
rect 85008 633134 85328 633218
rect 85008 632898 85050 633134
rect 85286 632898 85328 633134
rect 85008 632866 85328 632898
rect 115728 633454 116048 633486
rect 115728 633218 115770 633454
rect 116006 633218 116048 633454
rect 115728 633134 116048 633218
rect 115728 632898 115770 633134
rect 116006 632898 116048 633134
rect 115728 632866 116048 632898
rect 146448 633454 146768 633486
rect 146448 633218 146490 633454
rect 146726 633218 146768 633454
rect 146448 633134 146768 633218
rect 146448 632898 146490 633134
rect 146726 632898 146768 633134
rect 146448 632866 146768 632898
rect 177168 633454 177488 633486
rect 177168 633218 177210 633454
rect 177446 633218 177488 633454
rect 177168 633134 177488 633218
rect 177168 632898 177210 633134
rect 177446 632898 177488 633134
rect 177168 632866 177488 632898
rect 207888 633454 208208 633486
rect 207888 633218 207930 633454
rect 208166 633218 208208 633454
rect 207888 633134 208208 633218
rect 207888 632898 207930 633134
rect 208166 632898 208208 633134
rect 207888 632866 208208 632898
rect 238608 633454 238928 633486
rect 238608 633218 238650 633454
rect 238886 633218 238928 633454
rect 238608 633134 238928 633218
rect 238608 632898 238650 633134
rect 238886 632898 238928 633134
rect 238608 632866 238928 632898
rect 269328 633454 269648 633486
rect 269328 633218 269370 633454
rect 269606 633218 269648 633454
rect 269328 633134 269648 633218
rect 269328 632898 269370 633134
rect 269606 632898 269648 633134
rect 269328 632866 269648 632898
rect 300048 633454 300368 633486
rect 300048 633218 300090 633454
rect 300326 633218 300368 633454
rect 300048 633134 300368 633218
rect 300048 632898 300090 633134
rect 300326 632898 300368 633134
rect 300048 632866 300368 632898
rect 330768 633454 331088 633486
rect 330768 633218 330810 633454
rect 331046 633218 331088 633454
rect 330768 633134 331088 633218
rect 330768 632898 330810 633134
rect 331046 632898 331088 633134
rect 330768 632866 331088 632898
rect 361488 633454 361808 633486
rect 361488 633218 361530 633454
rect 361766 633218 361808 633454
rect 361488 633134 361808 633218
rect 361488 632898 361530 633134
rect 361766 632898 361808 633134
rect 361488 632866 361808 632898
rect 392208 633454 392528 633486
rect 392208 633218 392250 633454
rect 392486 633218 392528 633454
rect 392208 633134 392528 633218
rect 392208 632898 392250 633134
rect 392486 632898 392528 633134
rect 392208 632866 392528 632898
rect 422928 633454 423248 633486
rect 422928 633218 422970 633454
rect 423206 633218 423248 633454
rect 422928 633134 423248 633218
rect 422928 632898 422970 633134
rect 423206 632898 423248 633134
rect 422928 632866 423248 632898
rect 453648 633454 453968 633486
rect 453648 633218 453690 633454
rect 453926 633218 453968 633454
rect 453648 633134 453968 633218
rect 453648 632898 453690 633134
rect 453926 632898 453968 633134
rect 453648 632866 453968 632898
rect 484368 633454 484688 633486
rect 484368 633218 484410 633454
rect 484646 633218 484688 633454
rect 484368 633134 484688 633218
rect 484368 632898 484410 633134
rect 484646 632898 484688 633134
rect 484368 632866 484688 632898
rect 515088 633454 515408 633486
rect 515088 633218 515130 633454
rect 515366 633218 515408 633454
rect 515088 633134 515408 633218
rect 515088 632898 515130 633134
rect 515366 632898 515408 633134
rect 515088 632866 515408 632898
rect 545808 633454 546128 633486
rect 545808 633218 545850 633454
rect 546086 633218 546128 633454
rect 545808 633134 546128 633218
rect 545808 632898 545850 633134
rect 546086 632898 546128 633134
rect 545808 632866 546128 632898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect 8208 615454 8528 615486
rect 8208 615218 8250 615454
rect 8486 615218 8528 615454
rect 8208 615134 8528 615218
rect 8208 614898 8250 615134
rect 8486 614898 8528 615134
rect 8208 614866 8528 614898
rect 38928 615454 39248 615486
rect 38928 615218 38970 615454
rect 39206 615218 39248 615454
rect 38928 615134 39248 615218
rect 38928 614898 38970 615134
rect 39206 614898 39248 615134
rect 38928 614866 39248 614898
rect 69648 615454 69968 615486
rect 69648 615218 69690 615454
rect 69926 615218 69968 615454
rect 69648 615134 69968 615218
rect 69648 614898 69690 615134
rect 69926 614898 69968 615134
rect 69648 614866 69968 614898
rect 100368 615454 100688 615486
rect 100368 615218 100410 615454
rect 100646 615218 100688 615454
rect 100368 615134 100688 615218
rect 100368 614898 100410 615134
rect 100646 614898 100688 615134
rect 100368 614866 100688 614898
rect 131088 615454 131408 615486
rect 131088 615218 131130 615454
rect 131366 615218 131408 615454
rect 131088 615134 131408 615218
rect 131088 614898 131130 615134
rect 131366 614898 131408 615134
rect 131088 614866 131408 614898
rect 161808 615454 162128 615486
rect 161808 615218 161850 615454
rect 162086 615218 162128 615454
rect 161808 615134 162128 615218
rect 161808 614898 161850 615134
rect 162086 614898 162128 615134
rect 161808 614866 162128 614898
rect 192528 615454 192848 615486
rect 192528 615218 192570 615454
rect 192806 615218 192848 615454
rect 192528 615134 192848 615218
rect 192528 614898 192570 615134
rect 192806 614898 192848 615134
rect 192528 614866 192848 614898
rect 223248 615454 223568 615486
rect 223248 615218 223290 615454
rect 223526 615218 223568 615454
rect 223248 615134 223568 615218
rect 223248 614898 223290 615134
rect 223526 614898 223568 615134
rect 223248 614866 223568 614898
rect 253968 615454 254288 615486
rect 253968 615218 254010 615454
rect 254246 615218 254288 615454
rect 253968 615134 254288 615218
rect 253968 614898 254010 615134
rect 254246 614898 254288 615134
rect 253968 614866 254288 614898
rect 284688 615454 285008 615486
rect 284688 615218 284730 615454
rect 284966 615218 285008 615454
rect 284688 615134 285008 615218
rect 284688 614898 284730 615134
rect 284966 614898 285008 615134
rect 284688 614866 285008 614898
rect 315408 615454 315728 615486
rect 315408 615218 315450 615454
rect 315686 615218 315728 615454
rect 315408 615134 315728 615218
rect 315408 614898 315450 615134
rect 315686 614898 315728 615134
rect 315408 614866 315728 614898
rect 346128 615454 346448 615486
rect 346128 615218 346170 615454
rect 346406 615218 346448 615454
rect 346128 615134 346448 615218
rect 346128 614898 346170 615134
rect 346406 614898 346448 615134
rect 346128 614866 346448 614898
rect 376848 615454 377168 615486
rect 376848 615218 376890 615454
rect 377126 615218 377168 615454
rect 376848 615134 377168 615218
rect 376848 614898 376890 615134
rect 377126 614898 377168 615134
rect 376848 614866 377168 614898
rect 407568 615454 407888 615486
rect 407568 615218 407610 615454
rect 407846 615218 407888 615454
rect 407568 615134 407888 615218
rect 407568 614898 407610 615134
rect 407846 614898 407888 615134
rect 407568 614866 407888 614898
rect 438288 615454 438608 615486
rect 438288 615218 438330 615454
rect 438566 615218 438608 615454
rect 438288 615134 438608 615218
rect 438288 614898 438330 615134
rect 438566 614898 438608 615134
rect 438288 614866 438608 614898
rect 469008 615454 469328 615486
rect 469008 615218 469050 615454
rect 469286 615218 469328 615454
rect 469008 615134 469328 615218
rect 469008 614898 469050 615134
rect 469286 614898 469328 615134
rect 469008 614866 469328 614898
rect 499728 615454 500048 615486
rect 499728 615218 499770 615454
rect 500006 615218 500048 615454
rect 499728 615134 500048 615218
rect 499728 614898 499770 615134
rect 500006 614898 500048 615134
rect 499728 614866 500048 614898
rect 530448 615454 530768 615486
rect 530448 615218 530490 615454
rect 530726 615218 530768 615454
rect 530448 615134 530768 615218
rect 530448 614898 530490 615134
rect 530726 614898 530768 615134
rect 530448 614866 530768 614898
rect 561168 615454 561488 615486
rect 561168 615218 561210 615454
rect 561446 615218 561488 615454
rect 561168 615134 561488 615218
rect 561168 614898 561210 615134
rect 561446 614898 561488 615134
rect 561168 614866 561488 614898
rect 567234 604894 567854 640338
rect 567234 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 567854 604894
rect 567234 604574 567854 604658
rect 567234 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 567854 604574
rect 23568 597454 23888 597486
rect 23568 597218 23610 597454
rect 23846 597218 23888 597454
rect 23568 597134 23888 597218
rect 23568 596898 23610 597134
rect 23846 596898 23888 597134
rect 23568 596866 23888 596898
rect 54288 597454 54608 597486
rect 54288 597218 54330 597454
rect 54566 597218 54608 597454
rect 54288 597134 54608 597218
rect 54288 596898 54330 597134
rect 54566 596898 54608 597134
rect 54288 596866 54608 596898
rect 85008 597454 85328 597486
rect 85008 597218 85050 597454
rect 85286 597218 85328 597454
rect 85008 597134 85328 597218
rect 85008 596898 85050 597134
rect 85286 596898 85328 597134
rect 85008 596866 85328 596898
rect 115728 597454 116048 597486
rect 115728 597218 115770 597454
rect 116006 597218 116048 597454
rect 115728 597134 116048 597218
rect 115728 596898 115770 597134
rect 116006 596898 116048 597134
rect 115728 596866 116048 596898
rect 146448 597454 146768 597486
rect 146448 597218 146490 597454
rect 146726 597218 146768 597454
rect 146448 597134 146768 597218
rect 146448 596898 146490 597134
rect 146726 596898 146768 597134
rect 146448 596866 146768 596898
rect 177168 597454 177488 597486
rect 177168 597218 177210 597454
rect 177446 597218 177488 597454
rect 177168 597134 177488 597218
rect 177168 596898 177210 597134
rect 177446 596898 177488 597134
rect 177168 596866 177488 596898
rect 207888 597454 208208 597486
rect 207888 597218 207930 597454
rect 208166 597218 208208 597454
rect 207888 597134 208208 597218
rect 207888 596898 207930 597134
rect 208166 596898 208208 597134
rect 207888 596866 208208 596898
rect 238608 597454 238928 597486
rect 238608 597218 238650 597454
rect 238886 597218 238928 597454
rect 238608 597134 238928 597218
rect 238608 596898 238650 597134
rect 238886 596898 238928 597134
rect 238608 596866 238928 596898
rect 269328 597454 269648 597486
rect 269328 597218 269370 597454
rect 269606 597218 269648 597454
rect 269328 597134 269648 597218
rect 269328 596898 269370 597134
rect 269606 596898 269648 597134
rect 269328 596866 269648 596898
rect 300048 597454 300368 597486
rect 300048 597218 300090 597454
rect 300326 597218 300368 597454
rect 300048 597134 300368 597218
rect 300048 596898 300090 597134
rect 300326 596898 300368 597134
rect 300048 596866 300368 596898
rect 330768 597454 331088 597486
rect 330768 597218 330810 597454
rect 331046 597218 331088 597454
rect 330768 597134 331088 597218
rect 330768 596898 330810 597134
rect 331046 596898 331088 597134
rect 330768 596866 331088 596898
rect 361488 597454 361808 597486
rect 361488 597218 361530 597454
rect 361766 597218 361808 597454
rect 361488 597134 361808 597218
rect 361488 596898 361530 597134
rect 361766 596898 361808 597134
rect 361488 596866 361808 596898
rect 392208 597454 392528 597486
rect 392208 597218 392250 597454
rect 392486 597218 392528 597454
rect 392208 597134 392528 597218
rect 392208 596898 392250 597134
rect 392486 596898 392528 597134
rect 392208 596866 392528 596898
rect 422928 597454 423248 597486
rect 422928 597218 422970 597454
rect 423206 597218 423248 597454
rect 422928 597134 423248 597218
rect 422928 596898 422970 597134
rect 423206 596898 423248 597134
rect 422928 596866 423248 596898
rect 453648 597454 453968 597486
rect 453648 597218 453690 597454
rect 453926 597218 453968 597454
rect 453648 597134 453968 597218
rect 453648 596898 453690 597134
rect 453926 596898 453968 597134
rect 453648 596866 453968 596898
rect 484368 597454 484688 597486
rect 484368 597218 484410 597454
rect 484646 597218 484688 597454
rect 484368 597134 484688 597218
rect 484368 596898 484410 597134
rect 484646 596898 484688 597134
rect 484368 596866 484688 596898
rect 515088 597454 515408 597486
rect 515088 597218 515130 597454
rect 515366 597218 515408 597454
rect 515088 597134 515408 597218
rect 515088 596898 515130 597134
rect 515366 596898 515408 597134
rect 515088 596866 515408 596898
rect 545808 597454 546128 597486
rect 545808 597218 545850 597454
rect 546086 597218 546128 597454
rect 545808 597134 546128 597218
rect 545808 596898 545850 597134
rect 546086 596898 546128 597134
rect 545808 596866 546128 596898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect 8208 579454 8528 579486
rect 8208 579218 8250 579454
rect 8486 579218 8528 579454
rect 8208 579134 8528 579218
rect 8208 578898 8250 579134
rect 8486 578898 8528 579134
rect 8208 578866 8528 578898
rect 38928 579454 39248 579486
rect 38928 579218 38970 579454
rect 39206 579218 39248 579454
rect 38928 579134 39248 579218
rect 38928 578898 38970 579134
rect 39206 578898 39248 579134
rect 38928 578866 39248 578898
rect 69648 579454 69968 579486
rect 69648 579218 69690 579454
rect 69926 579218 69968 579454
rect 69648 579134 69968 579218
rect 69648 578898 69690 579134
rect 69926 578898 69968 579134
rect 69648 578866 69968 578898
rect 100368 579454 100688 579486
rect 100368 579218 100410 579454
rect 100646 579218 100688 579454
rect 100368 579134 100688 579218
rect 100368 578898 100410 579134
rect 100646 578898 100688 579134
rect 100368 578866 100688 578898
rect 131088 579454 131408 579486
rect 131088 579218 131130 579454
rect 131366 579218 131408 579454
rect 131088 579134 131408 579218
rect 131088 578898 131130 579134
rect 131366 578898 131408 579134
rect 131088 578866 131408 578898
rect 161808 579454 162128 579486
rect 161808 579218 161850 579454
rect 162086 579218 162128 579454
rect 161808 579134 162128 579218
rect 161808 578898 161850 579134
rect 162086 578898 162128 579134
rect 161808 578866 162128 578898
rect 192528 579454 192848 579486
rect 192528 579218 192570 579454
rect 192806 579218 192848 579454
rect 192528 579134 192848 579218
rect 192528 578898 192570 579134
rect 192806 578898 192848 579134
rect 192528 578866 192848 578898
rect 223248 579454 223568 579486
rect 223248 579218 223290 579454
rect 223526 579218 223568 579454
rect 223248 579134 223568 579218
rect 223248 578898 223290 579134
rect 223526 578898 223568 579134
rect 223248 578866 223568 578898
rect 253968 579454 254288 579486
rect 253968 579218 254010 579454
rect 254246 579218 254288 579454
rect 253968 579134 254288 579218
rect 253968 578898 254010 579134
rect 254246 578898 254288 579134
rect 253968 578866 254288 578898
rect 284688 579454 285008 579486
rect 284688 579218 284730 579454
rect 284966 579218 285008 579454
rect 284688 579134 285008 579218
rect 284688 578898 284730 579134
rect 284966 578898 285008 579134
rect 284688 578866 285008 578898
rect 315408 579454 315728 579486
rect 315408 579218 315450 579454
rect 315686 579218 315728 579454
rect 315408 579134 315728 579218
rect 315408 578898 315450 579134
rect 315686 578898 315728 579134
rect 315408 578866 315728 578898
rect 346128 579454 346448 579486
rect 346128 579218 346170 579454
rect 346406 579218 346448 579454
rect 346128 579134 346448 579218
rect 346128 578898 346170 579134
rect 346406 578898 346448 579134
rect 346128 578866 346448 578898
rect 376848 579454 377168 579486
rect 376848 579218 376890 579454
rect 377126 579218 377168 579454
rect 376848 579134 377168 579218
rect 376848 578898 376890 579134
rect 377126 578898 377168 579134
rect 376848 578866 377168 578898
rect 407568 579454 407888 579486
rect 407568 579218 407610 579454
rect 407846 579218 407888 579454
rect 407568 579134 407888 579218
rect 407568 578898 407610 579134
rect 407846 578898 407888 579134
rect 407568 578866 407888 578898
rect 438288 579454 438608 579486
rect 438288 579218 438330 579454
rect 438566 579218 438608 579454
rect 438288 579134 438608 579218
rect 438288 578898 438330 579134
rect 438566 578898 438608 579134
rect 438288 578866 438608 578898
rect 469008 579454 469328 579486
rect 469008 579218 469050 579454
rect 469286 579218 469328 579454
rect 469008 579134 469328 579218
rect 469008 578898 469050 579134
rect 469286 578898 469328 579134
rect 469008 578866 469328 578898
rect 499728 579454 500048 579486
rect 499728 579218 499770 579454
rect 500006 579218 500048 579454
rect 499728 579134 500048 579218
rect 499728 578898 499770 579134
rect 500006 578898 500048 579134
rect 499728 578866 500048 578898
rect 530448 579454 530768 579486
rect 530448 579218 530490 579454
rect 530726 579218 530768 579454
rect 530448 579134 530768 579218
rect 530448 578898 530490 579134
rect 530726 578898 530768 579134
rect 530448 578866 530768 578898
rect 561168 579454 561488 579486
rect 561168 579218 561210 579454
rect 561446 579218 561488 579454
rect 561168 579134 561488 579218
rect 561168 578898 561210 579134
rect 561446 578898 561488 579134
rect 561168 578866 561488 578898
rect 567234 568894 567854 604338
rect 567234 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 567854 568894
rect 567234 568574 567854 568658
rect 567234 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 567854 568574
rect 23568 561454 23888 561486
rect 23568 561218 23610 561454
rect 23846 561218 23888 561454
rect 23568 561134 23888 561218
rect 23568 560898 23610 561134
rect 23846 560898 23888 561134
rect 23568 560866 23888 560898
rect 54288 561454 54608 561486
rect 54288 561218 54330 561454
rect 54566 561218 54608 561454
rect 54288 561134 54608 561218
rect 54288 560898 54330 561134
rect 54566 560898 54608 561134
rect 54288 560866 54608 560898
rect 85008 561454 85328 561486
rect 85008 561218 85050 561454
rect 85286 561218 85328 561454
rect 85008 561134 85328 561218
rect 85008 560898 85050 561134
rect 85286 560898 85328 561134
rect 85008 560866 85328 560898
rect 115728 561454 116048 561486
rect 115728 561218 115770 561454
rect 116006 561218 116048 561454
rect 115728 561134 116048 561218
rect 115728 560898 115770 561134
rect 116006 560898 116048 561134
rect 115728 560866 116048 560898
rect 146448 561454 146768 561486
rect 146448 561218 146490 561454
rect 146726 561218 146768 561454
rect 146448 561134 146768 561218
rect 146448 560898 146490 561134
rect 146726 560898 146768 561134
rect 146448 560866 146768 560898
rect 177168 561454 177488 561486
rect 177168 561218 177210 561454
rect 177446 561218 177488 561454
rect 177168 561134 177488 561218
rect 177168 560898 177210 561134
rect 177446 560898 177488 561134
rect 177168 560866 177488 560898
rect 207888 561454 208208 561486
rect 207888 561218 207930 561454
rect 208166 561218 208208 561454
rect 207888 561134 208208 561218
rect 207888 560898 207930 561134
rect 208166 560898 208208 561134
rect 207888 560866 208208 560898
rect 238608 561454 238928 561486
rect 238608 561218 238650 561454
rect 238886 561218 238928 561454
rect 238608 561134 238928 561218
rect 238608 560898 238650 561134
rect 238886 560898 238928 561134
rect 238608 560866 238928 560898
rect 269328 561454 269648 561486
rect 269328 561218 269370 561454
rect 269606 561218 269648 561454
rect 269328 561134 269648 561218
rect 269328 560898 269370 561134
rect 269606 560898 269648 561134
rect 269328 560866 269648 560898
rect 300048 561454 300368 561486
rect 300048 561218 300090 561454
rect 300326 561218 300368 561454
rect 300048 561134 300368 561218
rect 300048 560898 300090 561134
rect 300326 560898 300368 561134
rect 300048 560866 300368 560898
rect 330768 561454 331088 561486
rect 330768 561218 330810 561454
rect 331046 561218 331088 561454
rect 330768 561134 331088 561218
rect 330768 560898 330810 561134
rect 331046 560898 331088 561134
rect 330768 560866 331088 560898
rect 361488 561454 361808 561486
rect 361488 561218 361530 561454
rect 361766 561218 361808 561454
rect 361488 561134 361808 561218
rect 361488 560898 361530 561134
rect 361766 560898 361808 561134
rect 361488 560866 361808 560898
rect 392208 561454 392528 561486
rect 392208 561218 392250 561454
rect 392486 561218 392528 561454
rect 392208 561134 392528 561218
rect 392208 560898 392250 561134
rect 392486 560898 392528 561134
rect 392208 560866 392528 560898
rect 422928 561454 423248 561486
rect 422928 561218 422970 561454
rect 423206 561218 423248 561454
rect 422928 561134 423248 561218
rect 422928 560898 422970 561134
rect 423206 560898 423248 561134
rect 422928 560866 423248 560898
rect 453648 561454 453968 561486
rect 453648 561218 453690 561454
rect 453926 561218 453968 561454
rect 453648 561134 453968 561218
rect 453648 560898 453690 561134
rect 453926 560898 453968 561134
rect 453648 560866 453968 560898
rect 484368 561454 484688 561486
rect 484368 561218 484410 561454
rect 484646 561218 484688 561454
rect 484368 561134 484688 561218
rect 484368 560898 484410 561134
rect 484646 560898 484688 561134
rect 484368 560866 484688 560898
rect 515088 561454 515408 561486
rect 515088 561218 515130 561454
rect 515366 561218 515408 561454
rect 515088 561134 515408 561218
rect 515088 560898 515130 561134
rect 515366 560898 515408 561134
rect 515088 560866 515408 560898
rect 545808 561454 546128 561486
rect 545808 561218 545850 561454
rect 546086 561218 546128 561454
rect 545808 561134 546128 561218
rect 545808 560898 545850 561134
rect 546086 560898 546128 561134
rect 545808 560866 546128 560898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect 8208 543454 8528 543486
rect 8208 543218 8250 543454
rect 8486 543218 8528 543454
rect 8208 543134 8528 543218
rect 8208 542898 8250 543134
rect 8486 542898 8528 543134
rect 8208 542866 8528 542898
rect 38928 543454 39248 543486
rect 38928 543218 38970 543454
rect 39206 543218 39248 543454
rect 38928 543134 39248 543218
rect 38928 542898 38970 543134
rect 39206 542898 39248 543134
rect 38928 542866 39248 542898
rect 69648 543454 69968 543486
rect 69648 543218 69690 543454
rect 69926 543218 69968 543454
rect 69648 543134 69968 543218
rect 69648 542898 69690 543134
rect 69926 542898 69968 543134
rect 69648 542866 69968 542898
rect 100368 543454 100688 543486
rect 100368 543218 100410 543454
rect 100646 543218 100688 543454
rect 100368 543134 100688 543218
rect 100368 542898 100410 543134
rect 100646 542898 100688 543134
rect 100368 542866 100688 542898
rect 131088 543454 131408 543486
rect 131088 543218 131130 543454
rect 131366 543218 131408 543454
rect 131088 543134 131408 543218
rect 131088 542898 131130 543134
rect 131366 542898 131408 543134
rect 131088 542866 131408 542898
rect 161808 543454 162128 543486
rect 161808 543218 161850 543454
rect 162086 543218 162128 543454
rect 161808 543134 162128 543218
rect 161808 542898 161850 543134
rect 162086 542898 162128 543134
rect 161808 542866 162128 542898
rect 192528 543454 192848 543486
rect 192528 543218 192570 543454
rect 192806 543218 192848 543454
rect 192528 543134 192848 543218
rect 192528 542898 192570 543134
rect 192806 542898 192848 543134
rect 192528 542866 192848 542898
rect 223248 543454 223568 543486
rect 223248 543218 223290 543454
rect 223526 543218 223568 543454
rect 223248 543134 223568 543218
rect 223248 542898 223290 543134
rect 223526 542898 223568 543134
rect 223248 542866 223568 542898
rect 253968 543454 254288 543486
rect 253968 543218 254010 543454
rect 254246 543218 254288 543454
rect 253968 543134 254288 543218
rect 253968 542898 254010 543134
rect 254246 542898 254288 543134
rect 253968 542866 254288 542898
rect 284688 543454 285008 543486
rect 284688 543218 284730 543454
rect 284966 543218 285008 543454
rect 284688 543134 285008 543218
rect 284688 542898 284730 543134
rect 284966 542898 285008 543134
rect 284688 542866 285008 542898
rect 315408 543454 315728 543486
rect 315408 543218 315450 543454
rect 315686 543218 315728 543454
rect 315408 543134 315728 543218
rect 315408 542898 315450 543134
rect 315686 542898 315728 543134
rect 315408 542866 315728 542898
rect 346128 543454 346448 543486
rect 346128 543218 346170 543454
rect 346406 543218 346448 543454
rect 346128 543134 346448 543218
rect 346128 542898 346170 543134
rect 346406 542898 346448 543134
rect 346128 542866 346448 542898
rect 376848 543454 377168 543486
rect 376848 543218 376890 543454
rect 377126 543218 377168 543454
rect 376848 543134 377168 543218
rect 376848 542898 376890 543134
rect 377126 542898 377168 543134
rect 376848 542866 377168 542898
rect 407568 543454 407888 543486
rect 407568 543218 407610 543454
rect 407846 543218 407888 543454
rect 407568 543134 407888 543218
rect 407568 542898 407610 543134
rect 407846 542898 407888 543134
rect 407568 542866 407888 542898
rect 438288 543454 438608 543486
rect 438288 543218 438330 543454
rect 438566 543218 438608 543454
rect 438288 543134 438608 543218
rect 438288 542898 438330 543134
rect 438566 542898 438608 543134
rect 438288 542866 438608 542898
rect 469008 543454 469328 543486
rect 469008 543218 469050 543454
rect 469286 543218 469328 543454
rect 469008 543134 469328 543218
rect 469008 542898 469050 543134
rect 469286 542898 469328 543134
rect 469008 542866 469328 542898
rect 499728 543454 500048 543486
rect 499728 543218 499770 543454
rect 500006 543218 500048 543454
rect 499728 543134 500048 543218
rect 499728 542898 499770 543134
rect 500006 542898 500048 543134
rect 499728 542866 500048 542898
rect 530448 543454 530768 543486
rect 530448 543218 530490 543454
rect 530726 543218 530768 543454
rect 530448 543134 530768 543218
rect 530448 542898 530490 543134
rect 530726 542898 530768 543134
rect 530448 542866 530768 542898
rect 561168 543454 561488 543486
rect 561168 543218 561210 543454
rect 561446 543218 561488 543454
rect 561168 543134 561488 543218
rect 561168 542898 561210 543134
rect 561446 542898 561488 543134
rect 561168 542866 561488 542898
rect 567234 532894 567854 568338
rect 567234 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 567854 532894
rect 567234 532574 567854 532658
rect 567234 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 567854 532574
rect 23568 525454 23888 525486
rect 23568 525218 23610 525454
rect 23846 525218 23888 525454
rect 23568 525134 23888 525218
rect 23568 524898 23610 525134
rect 23846 524898 23888 525134
rect 23568 524866 23888 524898
rect 54288 525454 54608 525486
rect 54288 525218 54330 525454
rect 54566 525218 54608 525454
rect 54288 525134 54608 525218
rect 54288 524898 54330 525134
rect 54566 524898 54608 525134
rect 54288 524866 54608 524898
rect 85008 525454 85328 525486
rect 85008 525218 85050 525454
rect 85286 525218 85328 525454
rect 85008 525134 85328 525218
rect 85008 524898 85050 525134
rect 85286 524898 85328 525134
rect 85008 524866 85328 524898
rect 115728 525454 116048 525486
rect 115728 525218 115770 525454
rect 116006 525218 116048 525454
rect 115728 525134 116048 525218
rect 115728 524898 115770 525134
rect 116006 524898 116048 525134
rect 115728 524866 116048 524898
rect 146448 525454 146768 525486
rect 146448 525218 146490 525454
rect 146726 525218 146768 525454
rect 146448 525134 146768 525218
rect 146448 524898 146490 525134
rect 146726 524898 146768 525134
rect 146448 524866 146768 524898
rect 177168 525454 177488 525486
rect 177168 525218 177210 525454
rect 177446 525218 177488 525454
rect 177168 525134 177488 525218
rect 177168 524898 177210 525134
rect 177446 524898 177488 525134
rect 177168 524866 177488 524898
rect 207888 525454 208208 525486
rect 207888 525218 207930 525454
rect 208166 525218 208208 525454
rect 207888 525134 208208 525218
rect 207888 524898 207930 525134
rect 208166 524898 208208 525134
rect 207888 524866 208208 524898
rect 238608 525454 238928 525486
rect 238608 525218 238650 525454
rect 238886 525218 238928 525454
rect 238608 525134 238928 525218
rect 238608 524898 238650 525134
rect 238886 524898 238928 525134
rect 238608 524866 238928 524898
rect 269328 525454 269648 525486
rect 269328 525218 269370 525454
rect 269606 525218 269648 525454
rect 269328 525134 269648 525218
rect 269328 524898 269370 525134
rect 269606 524898 269648 525134
rect 269328 524866 269648 524898
rect 300048 525454 300368 525486
rect 300048 525218 300090 525454
rect 300326 525218 300368 525454
rect 300048 525134 300368 525218
rect 300048 524898 300090 525134
rect 300326 524898 300368 525134
rect 300048 524866 300368 524898
rect 330768 525454 331088 525486
rect 330768 525218 330810 525454
rect 331046 525218 331088 525454
rect 330768 525134 331088 525218
rect 330768 524898 330810 525134
rect 331046 524898 331088 525134
rect 330768 524866 331088 524898
rect 361488 525454 361808 525486
rect 361488 525218 361530 525454
rect 361766 525218 361808 525454
rect 361488 525134 361808 525218
rect 361488 524898 361530 525134
rect 361766 524898 361808 525134
rect 361488 524866 361808 524898
rect 392208 525454 392528 525486
rect 392208 525218 392250 525454
rect 392486 525218 392528 525454
rect 392208 525134 392528 525218
rect 392208 524898 392250 525134
rect 392486 524898 392528 525134
rect 392208 524866 392528 524898
rect 422928 525454 423248 525486
rect 422928 525218 422970 525454
rect 423206 525218 423248 525454
rect 422928 525134 423248 525218
rect 422928 524898 422970 525134
rect 423206 524898 423248 525134
rect 422928 524866 423248 524898
rect 453648 525454 453968 525486
rect 453648 525218 453690 525454
rect 453926 525218 453968 525454
rect 453648 525134 453968 525218
rect 453648 524898 453690 525134
rect 453926 524898 453968 525134
rect 453648 524866 453968 524898
rect 484368 525454 484688 525486
rect 484368 525218 484410 525454
rect 484646 525218 484688 525454
rect 484368 525134 484688 525218
rect 484368 524898 484410 525134
rect 484646 524898 484688 525134
rect 484368 524866 484688 524898
rect 515088 525454 515408 525486
rect 515088 525218 515130 525454
rect 515366 525218 515408 525454
rect 515088 525134 515408 525218
rect 515088 524898 515130 525134
rect 515366 524898 515408 525134
rect 515088 524866 515408 524898
rect 545808 525454 546128 525486
rect 545808 525218 545850 525454
rect 546086 525218 546128 525454
rect 545808 525134 546128 525218
rect 545808 524898 545850 525134
rect 546086 524898 546128 525134
rect 545808 524866 546128 524898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect 8208 507454 8528 507486
rect 8208 507218 8250 507454
rect 8486 507218 8528 507454
rect 8208 507134 8528 507218
rect 8208 506898 8250 507134
rect 8486 506898 8528 507134
rect 8208 506866 8528 506898
rect 38928 507454 39248 507486
rect 38928 507218 38970 507454
rect 39206 507218 39248 507454
rect 38928 507134 39248 507218
rect 38928 506898 38970 507134
rect 39206 506898 39248 507134
rect 38928 506866 39248 506898
rect 69648 507454 69968 507486
rect 69648 507218 69690 507454
rect 69926 507218 69968 507454
rect 69648 507134 69968 507218
rect 69648 506898 69690 507134
rect 69926 506898 69968 507134
rect 69648 506866 69968 506898
rect 100368 507454 100688 507486
rect 100368 507218 100410 507454
rect 100646 507218 100688 507454
rect 100368 507134 100688 507218
rect 100368 506898 100410 507134
rect 100646 506898 100688 507134
rect 100368 506866 100688 506898
rect 131088 507454 131408 507486
rect 131088 507218 131130 507454
rect 131366 507218 131408 507454
rect 131088 507134 131408 507218
rect 131088 506898 131130 507134
rect 131366 506898 131408 507134
rect 131088 506866 131408 506898
rect 161808 507454 162128 507486
rect 161808 507218 161850 507454
rect 162086 507218 162128 507454
rect 161808 507134 162128 507218
rect 161808 506898 161850 507134
rect 162086 506898 162128 507134
rect 161808 506866 162128 506898
rect 192528 507454 192848 507486
rect 192528 507218 192570 507454
rect 192806 507218 192848 507454
rect 192528 507134 192848 507218
rect 192528 506898 192570 507134
rect 192806 506898 192848 507134
rect 192528 506866 192848 506898
rect 223248 507454 223568 507486
rect 223248 507218 223290 507454
rect 223526 507218 223568 507454
rect 223248 507134 223568 507218
rect 223248 506898 223290 507134
rect 223526 506898 223568 507134
rect 223248 506866 223568 506898
rect 253968 507454 254288 507486
rect 253968 507218 254010 507454
rect 254246 507218 254288 507454
rect 253968 507134 254288 507218
rect 253968 506898 254010 507134
rect 254246 506898 254288 507134
rect 253968 506866 254288 506898
rect 284688 507454 285008 507486
rect 284688 507218 284730 507454
rect 284966 507218 285008 507454
rect 284688 507134 285008 507218
rect 284688 506898 284730 507134
rect 284966 506898 285008 507134
rect 284688 506866 285008 506898
rect 315408 507454 315728 507486
rect 315408 507218 315450 507454
rect 315686 507218 315728 507454
rect 315408 507134 315728 507218
rect 315408 506898 315450 507134
rect 315686 506898 315728 507134
rect 315408 506866 315728 506898
rect 346128 507454 346448 507486
rect 346128 507218 346170 507454
rect 346406 507218 346448 507454
rect 346128 507134 346448 507218
rect 346128 506898 346170 507134
rect 346406 506898 346448 507134
rect 346128 506866 346448 506898
rect 376848 507454 377168 507486
rect 376848 507218 376890 507454
rect 377126 507218 377168 507454
rect 376848 507134 377168 507218
rect 376848 506898 376890 507134
rect 377126 506898 377168 507134
rect 376848 506866 377168 506898
rect 407568 507454 407888 507486
rect 407568 507218 407610 507454
rect 407846 507218 407888 507454
rect 407568 507134 407888 507218
rect 407568 506898 407610 507134
rect 407846 506898 407888 507134
rect 407568 506866 407888 506898
rect 438288 507454 438608 507486
rect 438288 507218 438330 507454
rect 438566 507218 438608 507454
rect 438288 507134 438608 507218
rect 438288 506898 438330 507134
rect 438566 506898 438608 507134
rect 438288 506866 438608 506898
rect 469008 507454 469328 507486
rect 469008 507218 469050 507454
rect 469286 507218 469328 507454
rect 469008 507134 469328 507218
rect 469008 506898 469050 507134
rect 469286 506898 469328 507134
rect 469008 506866 469328 506898
rect 499728 507454 500048 507486
rect 499728 507218 499770 507454
rect 500006 507218 500048 507454
rect 499728 507134 500048 507218
rect 499728 506898 499770 507134
rect 500006 506898 500048 507134
rect 499728 506866 500048 506898
rect 530448 507454 530768 507486
rect 530448 507218 530490 507454
rect 530726 507218 530768 507454
rect 530448 507134 530768 507218
rect 530448 506898 530490 507134
rect 530726 506898 530768 507134
rect 530448 506866 530768 506898
rect 561168 507454 561488 507486
rect 561168 507218 561210 507454
rect 561446 507218 561488 507454
rect 561168 507134 561488 507218
rect 561168 506898 561210 507134
rect 561446 506898 561488 507134
rect 561168 506866 561488 506898
rect 567234 496894 567854 532338
rect 567234 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 567854 496894
rect 567234 496574 567854 496658
rect 567234 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 567854 496574
rect 23568 489454 23888 489486
rect 23568 489218 23610 489454
rect 23846 489218 23888 489454
rect 23568 489134 23888 489218
rect 23568 488898 23610 489134
rect 23846 488898 23888 489134
rect 23568 488866 23888 488898
rect 54288 489454 54608 489486
rect 54288 489218 54330 489454
rect 54566 489218 54608 489454
rect 54288 489134 54608 489218
rect 54288 488898 54330 489134
rect 54566 488898 54608 489134
rect 54288 488866 54608 488898
rect 85008 489454 85328 489486
rect 85008 489218 85050 489454
rect 85286 489218 85328 489454
rect 85008 489134 85328 489218
rect 85008 488898 85050 489134
rect 85286 488898 85328 489134
rect 85008 488866 85328 488898
rect 115728 489454 116048 489486
rect 115728 489218 115770 489454
rect 116006 489218 116048 489454
rect 115728 489134 116048 489218
rect 115728 488898 115770 489134
rect 116006 488898 116048 489134
rect 115728 488866 116048 488898
rect 146448 489454 146768 489486
rect 146448 489218 146490 489454
rect 146726 489218 146768 489454
rect 146448 489134 146768 489218
rect 146448 488898 146490 489134
rect 146726 488898 146768 489134
rect 146448 488866 146768 488898
rect 177168 489454 177488 489486
rect 177168 489218 177210 489454
rect 177446 489218 177488 489454
rect 177168 489134 177488 489218
rect 177168 488898 177210 489134
rect 177446 488898 177488 489134
rect 177168 488866 177488 488898
rect 207888 489454 208208 489486
rect 207888 489218 207930 489454
rect 208166 489218 208208 489454
rect 207888 489134 208208 489218
rect 207888 488898 207930 489134
rect 208166 488898 208208 489134
rect 207888 488866 208208 488898
rect 238608 489454 238928 489486
rect 238608 489218 238650 489454
rect 238886 489218 238928 489454
rect 238608 489134 238928 489218
rect 238608 488898 238650 489134
rect 238886 488898 238928 489134
rect 238608 488866 238928 488898
rect 269328 489454 269648 489486
rect 269328 489218 269370 489454
rect 269606 489218 269648 489454
rect 269328 489134 269648 489218
rect 269328 488898 269370 489134
rect 269606 488898 269648 489134
rect 269328 488866 269648 488898
rect 300048 489454 300368 489486
rect 300048 489218 300090 489454
rect 300326 489218 300368 489454
rect 300048 489134 300368 489218
rect 300048 488898 300090 489134
rect 300326 488898 300368 489134
rect 300048 488866 300368 488898
rect 330768 489454 331088 489486
rect 330768 489218 330810 489454
rect 331046 489218 331088 489454
rect 330768 489134 331088 489218
rect 330768 488898 330810 489134
rect 331046 488898 331088 489134
rect 330768 488866 331088 488898
rect 361488 489454 361808 489486
rect 361488 489218 361530 489454
rect 361766 489218 361808 489454
rect 361488 489134 361808 489218
rect 361488 488898 361530 489134
rect 361766 488898 361808 489134
rect 361488 488866 361808 488898
rect 392208 489454 392528 489486
rect 392208 489218 392250 489454
rect 392486 489218 392528 489454
rect 392208 489134 392528 489218
rect 392208 488898 392250 489134
rect 392486 488898 392528 489134
rect 392208 488866 392528 488898
rect 422928 489454 423248 489486
rect 422928 489218 422970 489454
rect 423206 489218 423248 489454
rect 422928 489134 423248 489218
rect 422928 488898 422970 489134
rect 423206 488898 423248 489134
rect 422928 488866 423248 488898
rect 453648 489454 453968 489486
rect 453648 489218 453690 489454
rect 453926 489218 453968 489454
rect 453648 489134 453968 489218
rect 453648 488898 453690 489134
rect 453926 488898 453968 489134
rect 453648 488866 453968 488898
rect 484368 489454 484688 489486
rect 484368 489218 484410 489454
rect 484646 489218 484688 489454
rect 484368 489134 484688 489218
rect 484368 488898 484410 489134
rect 484646 488898 484688 489134
rect 484368 488866 484688 488898
rect 515088 489454 515408 489486
rect 515088 489218 515130 489454
rect 515366 489218 515408 489454
rect 515088 489134 515408 489218
rect 515088 488898 515130 489134
rect 515366 488898 515408 489134
rect 515088 488866 515408 488898
rect 545808 489454 546128 489486
rect 545808 489218 545850 489454
rect 546086 489218 546128 489454
rect 545808 489134 546128 489218
rect 545808 488898 545850 489134
rect 546086 488898 546128 489134
rect 545808 488866 546128 488898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect 8208 471454 8528 471486
rect 8208 471218 8250 471454
rect 8486 471218 8528 471454
rect 8208 471134 8528 471218
rect 8208 470898 8250 471134
rect 8486 470898 8528 471134
rect 8208 470866 8528 470898
rect 38928 471454 39248 471486
rect 38928 471218 38970 471454
rect 39206 471218 39248 471454
rect 38928 471134 39248 471218
rect 38928 470898 38970 471134
rect 39206 470898 39248 471134
rect 38928 470866 39248 470898
rect 69648 471454 69968 471486
rect 69648 471218 69690 471454
rect 69926 471218 69968 471454
rect 69648 471134 69968 471218
rect 69648 470898 69690 471134
rect 69926 470898 69968 471134
rect 69648 470866 69968 470898
rect 100368 471454 100688 471486
rect 100368 471218 100410 471454
rect 100646 471218 100688 471454
rect 100368 471134 100688 471218
rect 100368 470898 100410 471134
rect 100646 470898 100688 471134
rect 100368 470866 100688 470898
rect 131088 471454 131408 471486
rect 131088 471218 131130 471454
rect 131366 471218 131408 471454
rect 131088 471134 131408 471218
rect 131088 470898 131130 471134
rect 131366 470898 131408 471134
rect 131088 470866 131408 470898
rect 161808 471454 162128 471486
rect 161808 471218 161850 471454
rect 162086 471218 162128 471454
rect 161808 471134 162128 471218
rect 161808 470898 161850 471134
rect 162086 470898 162128 471134
rect 161808 470866 162128 470898
rect 192528 471454 192848 471486
rect 192528 471218 192570 471454
rect 192806 471218 192848 471454
rect 192528 471134 192848 471218
rect 192528 470898 192570 471134
rect 192806 470898 192848 471134
rect 192528 470866 192848 470898
rect 223248 471454 223568 471486
rect 223248 471218 223290 471454
rect 223526 471218 223568 471454
rect 223248 471134 223568 471218
rect 223248 470898 223290 471134
rect 223526 470898 223568 471134
rect 223248 470866 223568 470898
rect 253968 471454 254288 471486
rect 253968 471218 254010 471454
rect 254246 471218 254288 471454
rect 253968 471134 254288 471218
rect 253968 470898 254010 471134
rect 254246 470898 254288 471134
rect 253968 470866 254288 470898
rect 284688 471454 285008 471486
rect 284688 471218 284730 471454
rect 284966 471218 285008 471454
rect 284688 471134 285008 471218
rect 284688 470898 284730 471134
rect 284966 470898 285008 471134
rect 284688 470866 285008 470898
rect 315408 471454 315728 471486
rect 315408 471218 315450 471454
rect 315686 471218 315728 471454
rect 315408 471134 315728 471218
rect 315408 470898 315450 471134
rect 315686 470898 315728 471134
rect 315408 470866 315728 470898
rect 346128 471454 346448 471486
rect 346128 471218 346170 471454
rect 346406 471218 346448 471454
rect 346128 471134 346448 471218
rect 346128 470898 346170 471134
rect 346406 470898 346448 471134
rect 346128 470866 346448 470898
rect 376848 471454 377168 471486
rect 376848 471218 376890 471454
rect 377126 471218 377168 471454
rect 376848 471134 377168 471218
rect 376848 470898 376890 471134
rect 377126 470898 377168 471134
rect 376848 470866 377168 470898
rect 407568 471454 407888 471486
rect 407568 471218 407610 471454
rect 407846 471218 407888 471454
rect 407568 471134 407888 471218
rect 407568 470898 407610 471134
rect 407846 470898 407888 471134
rect 407568 470866 407888 470898
rect 438288 471454 438608 471486
rect 438288 471218 438330 471454
rect 438566 471218 438608 471454
rect 438288 471134 438608 471218
rect 438288 470898 438330 471134
rect 438566 470898 438608 471134
rect 438288 470866 438608 470898
rect 469008 471454 469328 471486
rect 469008 471218 469050 471454
rect 469286 471218 469328 471454
rect 469008 471134 469328 471218
rect 469008 470898 469050 471134
rect 469286 470898 469328 471134
rect 469008 470866 469328 470898
rect 499728 471454 500048 471486
rect 499728 471218 499770 471454
rect 500006 471218 500048 471454
rect 499728 471134 500048 471218
rect 499728 470898 499770 471134
rect 500006 470898 500048 471134
rect 499728 470866 500048 470898
rect 530448 471454 530768 471486
rect 530448 471218 530490 471454
rect 530726 471218 530768 471454
rect 530448 471134 530768 471218
rect 530448 470898 530490 471134
rect 530726 470898 530768 471134
rect 530448 470866 530768 470898
rect 561168 471454 561488 471486
rect 561168 471218 561210 471454
rect 561446 471218 561488 471454
rect 561168 471134 561488 471218
rect 561168 470898 561210 471134
rect 561446 470898 561488 471134
rect 561168 470866 561488 470898
rect 567234 460894 567854 496338
rect 567234 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 567854 460894
rect 567234 460574 567854 460658
rect 567234 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 567854 460574
rect 23568 453454 23888 453486
rect 23568 453218 23610 453454
rect 23846 453218 23888 453454
rect 23568 453134 23888 453218
rect 23568 452898 23610 453134
rect 23846 452898 23888 453134
rect 23568 452866 23888 452898
rect 54288 453454 54608 453486
rect 54288 453218 54330 453454
rect 54566 453218 54608 453454
rect 54288 453134 54608 453218
rect 54288 452898 54330 453134
rect 54566 452898 54608 453134
rect 54288 452866 54608 452898
rect 85008 453454 85328 453486
rect 85008 453218 85050 453454
rect 85286 453218 85328 453454
rect 85008 453134 85328 453218
rect 85008 452898 85050 453134
rect 85286 452898 85328 453134
rect 85008 452866 85328 452898
rect 115728 453454 116048 453486
rect 115728 453218 115770 453454
rect 116006 453218 116048 453454
rect 115728 453134 116048 453218
rect 115728 452898 115770 453134
rect 116006 452898 116048 453134
rect 115728 452866 116048 452898
rect 146448 453454 146768 453486
rect 146448 453218 146490 453454
rect 146726 453218 146768 453454
rect 146448 453134 146768 453218
rect 146448 452898 146490 453134
rect 146726 452898 146768 453134
rect 146448 452866 146768 452898
rect 177168 453454 177488 453486
rect 177168 453218 177210 453454
rect 177446 453218 177488 453454
rect 177168 453134 177488 453218
rect 177168 452898 177210 453134
rect 177446 452898 177488 453134
rect 177168 452866 177488 452898
rect 207888 453454 208208 453486
rect 207888 453218 207930 453454
rect 208166 453218 208208 453454
rect 207888 453134 208208 453218
rect 207888 452898 207930 453134
rect 208166 452898 208208 453134
rect 207888 452866 208208 452898
rect 238608 453454 238928 453486
rect 238608 453218 238650 453454
rect 238886 453218 238928 453454
rect 238608 453134 238928 453218
rect 238608 452898 238650 453134
rect 238886 452898 238928 453134
rect 238608 452866 238928 452898
rect 269328 453454 269648 453486
rect 269328 453218 269370 453454
rect 269606 453218 269648 453454
rect 269328 453134 269648 453218
rect 269328 452898 269370 453134
rect 269606 452898 269648 453134
rect 269328 452866 269648 452898
rect 300048 453454 300368 453486
rect 300048 453218 300090 453454
rect 300326 453218 300368 453454
rect 300048 453134 300368 453218
rect 300048 452898 300090 453134
rect 300326 452898 300368 453134
rect 300048 452866 300368 452898
rect 330768 453454 331088 453486
rect 330768 453218 330810 453454
rect 331046 453218 331088 453454
rect 330768 453134 331088 453218
rect 330768 452898 330810 453134
rect 331046 452898 331088 453134
rect 330768 452866 331088 452898
rect 361488 453454 361808 453486
rect 361488 453218 361530 453454
rect 361766 453218 361808 453454
rect 361488 453134 361808 453218
rect 361488 452898 361530 453134
rect 361766 452898 361808 453134
rect 361488 452866 361808 452898
rect 392208 453454 392528 453486
rect 392208 453218 392250 453454
rect 392486 453218 392528 453454
rect 392208 453134 392528 453218
rect 392208 452898 392250 453134
rect 392486 452898 392528 453134
rect 392208 452866 392528 452898
rect 422928 453454 423248 453486
rect 422928 453218 422970 453454
rect 423206 453218 423248 453454
rect 422928 453134 423248 453218
rect 422928 452898 422970 453134
rect 423206 452898 423248 453134
rect 422928 452866 423248 452898
rect 453648 453454 453968 453486
rect 453648 453218 453690 453454
rect 453926 453218 453968 453454
rect 453648 453134 453968 453218
rect 453648 452898 453690 453134
rect 453926 452898 453968 453134
rect 453648 452866 453968 452898
rect 484368 453454 484688 453486
rect 484368 453218 484410 453454
rect 484646 453218 484688 453454
rect 484368 453134 484688 453218
rect 484368 452898 484410 453134
rect 484646 452898 484688 453134
rect 484368 452866 484688 452898
rect 515088 453454 515408 453486
rect 515088 453218 515130 453454
rect 515366 453218 515408 453454
rect 515088 453134 515408 453218
rect 515088 452898 515130 453134
rect 515366 452898 515408 453134
rect 515088 452866 515408 452898
rect 545808 453454 546128 453486
rect 545808 453218 545850 453454
rect 546086 453218 546128 453454
rect 545808 453134 546128 453218
rect 545808 452898 545850 453134
rect 546086 452898 546128 453134
rect 545808 452866 546128 452898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect 8208 435454 8528 435486
rect 8208 435218 8250 435454
rect 8486 435218 8528 435454
rect 8208 435134 8528 435218
rect 8208 434898 8250 435134
rect 8486 434898 8528 435134
rect 8208 434866 8528 434898
rect 38928 435454 39248 435486
rect 38928 435218 38970 435454
rect 39206 435218 39248 435454
rect 38928 435134 39248 435218
rect 38928 434898 38970 435134
rect 39206 434898 39248 435134
rect 38928 434866 39248 434898
rect 69648 435454 69968 435486
rect 69648 435218 69690 435454
rect 69926 435218 69968 435454
rect 69648 435134 69968 435218
rect 69648 434898 69690 435134
rect 69926 434898 69968 435134
rect 69648 434866 69968 434898
rect 100368 435454 100688 435486
rect 100368 435218 100410 435454
rect 100646 435218 100688 435454
rect 100368 435134 100688 435218
rect 100368 434898 100410 435134
rect 100646 434898 100688 435134
rect 100368 434866 100688 434898
rect 131088 435454 131408 435486
rect 131088 435218 131130 435454
rect 131366 435218 131408 435454
rect 131088 435134 131408 435218
rect 131088 434898 131130 435134
rect 131366 434898 131408 435134
rect 131088 434866 131408 434898
rect 161808 435454 162128 435486
rect 161808 435218 161850 435454
rect 162086 435218 162128 435454
rect 161808 435134 162128 435218
rect 161808 434898 161850 435134
rect 162086 434898 162128 435134
rect 161808 434866 162128 434898
rect 192528 435454 192848 435486
rect 192528 435218 192570 435454
rect 192806 435218 192848 435454
rect 192528 435134 192848 435218
rect 192528 434898 192570 435134
rect 192806 434898 192848 435134
rect 192528 434866 192848 434898
rect 223248 435454 223568 435486
rect 223248 435218 223290 435454
rect 223526 435218 223568 435454
rect 223248 435134 223568 435218
rect 223248 434898 223290 435134
rect 223526 434898 223568 435134
rect 223248 434866 223568 434898
rect 253968 435454 254288 435486
rect 253968 435218 254010 435454
rect 254246 435218 254288 435454
rect 253968 435134 254288 435218
rect 253968 434898 254010 435134
rect 254246 434898 254288 435134
rect 253968 434866 254288 434898
rect 284688 435454 285008 435486
rect 284688 435218 284730 435454
rect 284966 435218 285008 435454
rect 284688 435134 285008 435218
rect 284688 434898 284730 435134
rect 284966 434898 285008 435134
rect 284688 434866 285008 434898
rect 315408 435454 315728 435486
rect 315408 435218 315450 435454
rect 315686 435218 315728 435454
rect 315408 435134 315728 435218
rect 315408 434898 315450 435134
rect 315686 434898 315728 435134
rect 315408 434866 315728 434898
rect 346128 435454 346448 435486
rect 346128 435218 346170 435454
rect 346406 435218 346448 435454
rect 346128 435134 346448 435218
rect 346128 434898 346170 435134
rect 346406 434898 346448 435134
rect 346128 434866 346448 434898
rect 376848 435454 377168 435486
rect 376848 435218 376890 435454
rect 377126 435218 377168 435454
rect 376848 435134 377168 435218
rect 376848 434898 376890 435134
rect 377126 434898 377168 435134
rect 376848 434866 377168 434898
rect 407568 435454 407888 435486
rect 407568 435218 407610 435454
rect 407846 435218 407888 435454
rect 407568 435134 407888 435218
rect 407568 434898 407610 435134
rect 407846 434898 407888 435134
rect 407568 434866 407888 434898
rect 438288 435454 438608 435486
rect 438288 435218 438330 435454
rect 438566 435218 438608 435454
rect 438288 435134 438608 435218
rect 438288 434898 438330 435134
rect 438566 434898 438608 435134
rect 438288 434866 438608 434898
rect 469008 435454 469328 435486
rect 469008 435218 469050 435454
rect 469286 435218 469328 435454
rect 469008 435134 469328 435218
rect 469008 434898 469050 435134
rect 469286 434898 469328 435134
rect 469008 434866 469328 434898
rect 499728 435454 500048 435486
rect 499728 435218 499770 435454
rect 500006 435218 500048 435454
rect 499728 435134 500048 435218
rect 499728 434898 499770 435134
rect 500006 434898 500048 435134
rect 499728 434866 500048 434898
rect 530448 435454 530768 435486
rect 530448 435218 530490 435454
rect 530726 435218 530768 435454
rect 530448 435134 530768 435218
rect 530448 434898 530490 435134
rect 530726 434898 530768 435134
rect 530448 434866 530768 434898
rect 561168 435454 561488 435486
rect 561168 435218 561210 435454
rect 561446 435218 561488 435454
rect 561168 435134 561488 435218
rect 561168 434898 561210 435134
rect 561446 434898 561488 435134
rect 561168 434866 561488 434898
rect 567234 424894 567854 460338
rect 567234 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 567854 424894
rect 567234 424574 567854 424658
rect 567234 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 567854 424574
rect 23568 417454 23888 417486
rect 23568 417218 23610 417454
rect 23846 417218 23888 417454
rect 23568 417134 23888 417218
rect 23568 416898 23610 417134
rect 23846 416898 23888 417134
rect 23568 416866 23888 416898
rect 54288 417454 54608 417486
rect 54288 417218 54330 417454
rect 54566 417218 54608 417454
rect 54288 417134 54608 417218
rect 54288 416898 54330 417134
rect 54566 416898 54608 417134
rect 54288 416866 54608 416898
rect 85008 417454 85328 417486
rect 85008 417218 85050 417454
rect 85286 417218 85328 417454
rect 85008 417134 85328 417218
rect 85008 416898 85050 417134
rect 85286 416898 85328 417134
rect 85008 416866 85328 416898
rect 115728 417454 116048 417486
rect 115728 417218 115770 417454
rect 116006 417218 116048 417454
rect 115728 417134 116048 417218
rect 115728 416898 115770 417134
rect 116006 416898 116048 417134
rect 115728 416866 116048 416898
rect 146448 417454 146768 417486
rect 146448 417218 146490 417454
rect 146726 417218 146768 417454
rect 146448 417134 146768 417218
rect 146448 416898 146490 417134
rect 146726 416898 146768 417134
rect 146448 416866 146768 416898
rect 177168 417454 177488 417486
rect 177168 417218 177210 417454
rect 177446 417218 177488 417454
rect 177168 417134 177488 417218
rect 177168 416898 177210 417134
rect 177446 416898 177488 417134
rect 177168 416866 177488 416898
rect 207888 417454 208208 417486
rect 207888 417218 207930 417454
rect 208166 417218 208208 417454
rect 207888 417134 208208 417218
rect 207888 416898 207930 417134
rect 208166 416898 208208 417134
rect 207888 416866 208208 416898
rect 238608 417454 238928 417486
rect 238608 417218 238650 417454
rect 238886 417218 238928 417454
rect 238608 417134 238928 417218
rect 238608 416898 238650 417134
rect 238886 416898 238928 417134
rect 238608 416866 238928 416898
rect 269328 417454 269648 417486
rect 269328 417218 269370 417454
rect 269606 417218 269648 417454
rect 269328 417134 269648 417218
rect 269328 416898 269370 417134
rect 269606 416898 269648 417134
rect 269328 416866 269648 416898
rect 300048 417454 300368 417486
rect 300048 417218 300090 417454
rect 300326 417218 300368 417454
rect 300048 417134 300368 417218
rect 300048 416898 300090 417134
rect 300326 416898 300368 417134
rect 300048 416866 300368 416898
rect 330768 417454 331088 417486
rect 330768 417218 330810 417454
rect 331046 417218 331088 417454
rect 330768 417134 331088 417218
rect 330768 416898 330810 417134
rect 331046 416898 331088 417134
rect 330768 416866 331088 416898
rect 361488 417454 361808 417486
rect 361488 417218 361530 417454
rect 361766 417218 361808 417454
rect 361488 417134 361808 417218
rect 361488 416898 361530 417134
rect 361766 416898 361808 417134
rect 361488 416866 361808 416898
rect 392208 417454 392528 417486
rect 392208 417218 392250 417454
rect 392486 417218 392528 417454
rect 392208 417134 392528 417218
rect 392208 416898 392250 417134
rect 392486 416898 392528 417134
rect 392208 416866 392528 416898
rect 422928 417454 423248 417486
rect 422928 417218 422970 417454
rect 423206 417218 423248 417454
rect 422928 417134 423248 417218
rect 422928 416898 422970 417134
rect 423206 416898 423248 417134
rect 422928 416866 423248 416898
rect 453648 417454 453968 417486
rect 453648 417218 453690 417454
rect 453926 417218 453968 417454
rect 453648 417134 453968 417218
rect 453648 416898 453690 417134
rect 453926 416898 453968 417134
rect 453648 416866 453968 416898
rect 484368 417454 484688 417486
rect 484368 417218 484410 417454
rect 484646 417218 484688 417454
rect 484368 417134 484688 417218
rect 484368 416898 484410 417134
rect 484646 416898 484688 417134
rect 484368 416866 484688 416898
rect 515088 417454 515408 417486
rect 515088 417218 515130 417454
rect 515366 417218 515408 417454
rect 515088 417134 515408 417218
rect 515088 416898 515130 417134
rect 515366 416898 515408 417134
rect 515088 416866 515408 416898
rect 545808 417454 546128 417486
rect 545808 417218 545850 417454
rect 546086 417218 546128 417454
rect 545808 417134 546128 417218
rect 545808 416898 545850 417134
rect 546086 416898 546128 417134
rect 545808 416866 546128 416898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect 8208 399454 8528 399486
rect 8208 399218 8250 399454
rect 8486 399218 8528 399454
rect 8208 399134 8528 399218
rect 8208 398898 8250 399134
rect 8486 398898 8528 399134
rect 8208 398866 8528 398898
rect 38928 399454 39248 399486
rect 38928 399218 38970 399454
rect 39206 399218 39248 399454
rect 38928 399134 39248 399218
rect 38928 398898 38970 399134
rect 39206 398898 39248 399134
rect 38928 398866 39248 398898
rect 69648 399454 69968 399486
rect 69648 399218 69690 399454
rect 69926 399218 69968 399454
rect 69648 399134 69968 399218
rect 69648 398898 69690 399134
rect 69926 398898 69968 399134
rect 69648 398866 69968 398898
rect 100368 399454 100688 399486
rect 100368 399218 100410 399454
rect 100646 399218 100688 399454
rect 100368 399134 100688 399218
rect 100368 398898 100410 399134
rect 100646 398898 100688 399134
rect 100368 398866 100688 398898
rect 131088 399454 131408 399486
rect 131088 399218 131130 399454
rect 131366 399218 131408 399454
rect 131088 399134 131408 399218
rect 131088 398898 131130 399134
rect 131366 398898 131408 399134
rect 131088 398866 131408 398898
rect 161808 399454 162128 399486
rect 161808 399218 161850 399454
rect 162086 399218 162128 399454
rect 161808 399134 162128 399218
rect 161808 398898 161850 399134
rect 162086 398898 162128 399134
rect 161808 398866 162128 398898
rect 192528 399454 192848 399486
rect 192528 399218 192570 399454
rect 192806 399218 192848 399454
rect 192528 399134 192848 399218
rect 192528 398898 192570 399134
rect 192806 398898 192848 399134
rect 192528 398866 192848 398898
rect 223248 399454 223568 399486
rect 223248 399218 223290 399454
rect 223526 399218 223568 399454
rect 223248 399134 223568 399218
rect 223248 398898 223290 399134
rect 223526 398898 223568 399134
rect 223248 398866 223568 398898
rect 253968 399454 254288 399486
rect 253968 399218 254010 399454
rect 254246 399218 254288 399454
rect 253968 399134 254288 399218
rect 253968 398898 254010 399134
rect 254246 398898 254288 399134
rect 253968 398866 254288 398898
rect 284688 399454 285008 399486
rect 284688 399218 284730 399454
rect 284966 399218 285008 399454
rect 284688 399134 285008 399218
rect 284688 398898 284730 399134
rect 284966 398898 285008 399134
rect 284688 398866 285008 398898
rect 315408 399454 315728 399486
rect 315408 399218 315450 399454
rect 315686 399218 315728 399454
rect 315408 399134 315728 399218
rect 315408 398898 315450 399134
rect 315686 398898 315728 399134
rect 315408 398866 315728 398898
rect 346128 399454 346448 399486
rect 346128 399218 346170 399454
rect 346406 399218 346448 399454
rect 346128 399134 346448 399218
rect 346128 398898 346170 399134
rect 346406 398898 346448 399134
rect 346128 398866 346448 398898
rect 376848 399454 377168 399486
rect 376848 399218 376890 399454
rect 377126 399218 377168 399454
rect 376848 399134 377168 399218
rect 376848 398898 376890 399134
rect 377126 398898 377168 399134
rect 376848 398866 377168 398898
rect 407568 399454 407888 399486
rect 407568 399218 407610 399454
rect 407846 399218 407888 399454
rect 407568 399134 407888 399218
rect 407568 398898 407610 399134
rect 407846 398898 407888 399134
rect 407568 398866 407888 398898
rect 438288 399454 438608 399486
rect 438288 399218 438330 399454
rect 438566 399218 438608 399454
rect 438288 399134 438608 399218
rect 438288 398898 438330 399134
rect 438566 398898 438608 399134
rect 438288 398866 438608 398898
rect 469008 399454 469328 399486
rect 469008 399218 469050 399454
rect 469286 399218 469328 399454
rect 469008 399134 469328 399218
rect 469008 398898 469050 399134
rect 469286 398898 469328 399134
rect 469008 398866 469328 398898
rect 499728 399454 500048 399486
rect 499728 399218 499770 399454
rect 500006 399218 500048 399454
rect 499728 399134 500048 399218
rect 499728 398898 499770 399134
rect 500006 398898 500048 399134
rect 499728 398866 500048 398898
rect 530448 399454 530768 399486
rect 530448 399218 530490 399454
rect 530726 399218 530768 399454
rect 530448 399134 530768 399218
rect 530448 398898 530490 399134
rect 530726 398898 530768 399134
rect 530448 398866 530768 398898
rect 561168 399454 561488 399486
rect 561168 399218 561210 399454
rect 561446 399218 561488 399454
rect 561168 399134 561488 399218
rect 561168 398898 561210 399134
rect 561446 398898 561488 399134
rect 561168 398866 561488 398898
rect 567234 388894 567854 424338
rect 567234 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 567854 388894
rect 567234 388574 567854 388658
rect 567234 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 567854 388574
rect 23568 381454 23888 381486
rect 23568 381218 23610 381454
rect 23846 381218 23888 381454
rect 23568 381134 23888 381218
rect 23568 380898 23610 381134
rect 23846 380898 23888 381134
rect 23568 380866 23888 380898
rect 54288 381454 54608 381486
rect 54288 381218 54330 381454
rect 54566 381218 54608 381454
rect 54288 381134 54608 381218
rect 54288 380898 54330 381134
rect 54566 380898 54608 381134
rect 54288 380866 54608 380898
rect 85008 381454 85328 381486
rect 85008 381218 85050 381454
rect 85286 381218 85328 381454
rect 85008 381134 85328 381218
rect 85008 380898 85050 381134
rect 85286 380898 85328 381134
rect 85008 380866 85328 380898
rect 115728 381454 116048 381486
rect 115728 381218 115770 381454
rect 116006 381218 116048 381454
rect 115728 381134 116048 381218
rect 115728 380898 115770 381134
rect 116006 380898 116048 381134
rect 115728 380866 116048 380898
rect 146448 381454 146768 381486
rect 146448 381218 146490 381454
rect 146726 381218 146768 381454
rect 146448 381134 146768 381218
rect 146448 380898 146490 381134
rect 146726 380898 146768 381134
rect 146448 380866 146768 380898
rect 177168 381454 177488 381486
rect 177168 381218 177210 381454
rect 177446 381218 177488 381454
rect 177168 381134 177488 381218
rect 177168 380898 177210 381134
rect 177446 380898 177488 381134
rect 177168 380866 177488 380898
rect 207888 381454 208208 381486
rect 207888 381218 207930 381454
rect 208166 381218 208208 381454
rect 207888 381134 208208 381218
rect 207888 380898 207930 381134
rect 208166 380898 208208 381134
rect 207888 380866 208208 380898
rect 238608 381454 238928 381486
rect 238608 381218 238650 381454
rect 238886 381218 238928 381454
rect 238608 381134 238928 381218
rect 238608 380898 238650 381134
rect 238886 380898 238928 381134
rect 238608 380866 238928 380898
rect 269328 381454 269648 381486
rect 269328 381218 269370 381454
rect 269606 381218 269648 381454
rect 269328 381134 269648 381218
rect 269328 380898 269370 381134
rect 269606 380898 269648 381134
rect 269328 380866 269648 380898
rect 300048 381454 300368 381486
rect 300048 381218 300090 381454
rect 300326 381218 300368 381454
rect 300048 381134 300368 381218
rect 300048 380898 300090 381134
rect 300326 380898 300368 381134
rect 300048 380866 300368 380898
rect 330768 381454 331088 381486
rect 330768 381218 330810 381454
rect 331046 381218 331088 381454
rect 330768 381134 331088 381218
rect 330768 380898 330810 381134
rect 331046 380898 331088 381134
rect 330768 380866 331088 380898
rect 361488 381454 361808 381486
rect 361488 381218 361530 381454
rect 361766 381218 361808 381454
rect 361488 381134 361808 381218
rect 361488 380898 361530 381134
rect 361766 380898 361808 381134
rect 361488 380866 361808 380898
rect 392208 381454 392528 381486
rect 392208 381218 392250 381454
rect 392486 381218 392528 381454
rect 392208 381134 392528 381218
rect 392208 380898 392250 381134
rect 392486 380898 392528 381134
rect 392208 380866 392528 380898
rect 422928 381454 423248 381486
rect 422928 381218 422970 381454
rect 423206 381218 423248 381454
rect 422928 381134 423248 381218
rect 422928 380898 422970 381134
rect 423206 380898 423248 381134
rect 422928 380866 423248 380898
rect 453648 381454 453968 381486
rect 453648 381218 453690 381454
rect 453926 381218 453968 381454
rect 453648 381134 453968 381218
rect 453648 380898 453690 381134
rect 453926 380898 453968 381134
rect 453648 380866 453968 380898
rect 484368 381454 484688 381486
rect 484368 381218 484410 381454
rect 484646 381218 484688 381454
rect 484368 381134 484688 381218
rect 484368 380898 484410 381134
rect 484646 380898 484688 381134
rect 484368 380866 484688 380898
rect 515088 381454 515408 381486
rect 515088 381218 515130 381454
rect 515366 381218 515408 381454
rect 515088 381134 515408 381218
rect 515088 380898 515130 381134
rect 515366 380898 515408 381134
rect 515088 380866 515408 380898
rect 545808 381454 546128 381486
rect 545808 381218 545850 381454
rect 546086 381218 546128 381454
rect 545808 381134 546128 381218
rect 545808 380898 545850 381134
rect 546086 380898 546128 381134
rect 545808 380866 546128 380898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect 8208 363454 8528 363486
rect 8208 363218 8250 363454
rect 8486 363218 8528 363454
rect 8208 363134 8528 363218
rect 8208 362898 8250 363134
rect 8486 362898 8528 363134
rect 8208 362866 8528 362898
rect 38928 363454 39248 363486
rect 38928 363218 38970 363454
rect 39206 363218 39248 363454
rect 38928 363134 39248 363218
rect 38928 362898 38970 363134
rect 39206 362898 39248 363134
rect 38928 362866 39248 362898
rect 69648 363454 69968 363486
rect 69648 363218 69690 363454
rect 69926 363218 69968 363454
rect 69648 363134 69968 363218
rect 69648 362898 69690 363134
rect 69926 362898 69968 363134
rect 69648 362866 69968 362898
rect 100368 363454 100688 363486
rect 100368 363218 100410 363454
rect 100646 363218 100688 363454
rect 100368 363134 100688 363218
rect 100368 362898 100410 363134
rect 100646 362898 100688 363134
rect 100368 362866 100688 362898
rect 131088 363454 131408 363486
rect 131088 363218 131130 363454
rect 131366 363218 131408 363454
rect 131088 363134 131408 363218
rect 131088 362898 131130 363134
rect 131366 362898 131408 363134
rect 131088 362866 131408 362898
rect 161808 363454 162128 363486
rect 161808 363218 161850 363454
rect 162086 363218 162128 363454
rect 161808 363134 162128 363218
rect 161808 362898 161850 363134
rect 162086 362898 162128 363134
rect 161808 362866 162128 362898
rect 192528 363454 192848 363486
rect 192528 363218 192570 363454
rect 192806 363218 192848 363454
rect 192528 363134 192848 363218
rect 192528 362898 192570 363134
rect 192806 362898 192848 363134
rect 192528 362866 192848 362898
rect 223248 363454 223568 363486
rect 223248 363218 223290 363454
rect 223526 363218 223568 363454
rect 223248 363134 223568 363218
rect 223248 362898 223290 363134
rect 223526 362898 223568 363134
rect 223248 362866 223568 362898
rect 253968 363454 254288 363486
rect 253968 363218 254010 363454
rect 254246 363218 254288 363454
rect 253968 363134 254288 363218
rect 253968 362898 254010 363134
rect 254246 362898 254288 363134
rect 253968 362866 254288 362898
rect 284688 363454 285008 363486
rect 284688 363218 284730 363454
rect 284966 363218 285008 363454
rect 284688 363134 285008 363218
rect 284688 362898 284730 363134
rect 284966 362898 285008 363134
rect 284688 362866 285008 362898
rect 315408 363454 315728 363486
rect 315408 363218 315450 363454
rect 315686 363218 315728 363454
rect 315408 363134 315728 363218
rect 315408 362898 315450 363134
rect 315686 362898 315728 363134
rect 315408 362866 315728 362898
rect 346128 363454 346448 363486
rect 346128 363218 346170 363454
rect 346406 363218 346448 363454
rect 346128 363134 346448 363218
rect 346128 362898 346170 363134
rect 346406 362898 346448 363134
rect 346128 362866 346448 362898
rect 376848 363454 377168 363486
rect 376848 363218 376890 363454
rect 377126 363218 377168 363454
rect 376848 363134 377168 363218
rect 376848 362898 376890 363134
rect 377126 362898 377168 363134
rect 376848 362866 377168 362898
rect 407568 363454 407888 363486
rect 407568 363218 407610 363454
rect 407846 363218 407888 363454
rect 407568 363134 407888 363218
rect 407568 362898 407610 363134
rect 407846 362898 407888 363134
rect 407568 362866 407888 362898
rect 438288 363454 438608 363486
rect 438288 363218 438330 363454
rect 438566 363218 438608 363454
rect 438288 363134 438608 363218
rect 438288 362898 438330 363134
rect 438566 362898 438608 363134
rect 438288 362866 438608 362898
rect 469008 363454 469328 363486
rect 469008 363218 469050 363454
rect 469286 363218 469328 363454
rect 469008 363134 469328 363218
rect 469008 362898 469050 363134
rect 469286 362898 469328 363134
rect 469008 362866 469328 362898
rect 499728 363454 500048 363486
rect 499728 363218 499770 363454
rect 500006 363218 500048 363454
rect 499728 363134 500048 363218
rect 499728 362898 499770 363134
rect 500006 362898 500048 363134
rect 499728 362866 500048 362898
rect 530448 363454 530768 363486
rect 530448 363218 530490 363454
rect 530726 363218 530768 363454
rect 530448 363134 530768 363218
rect 530448 362898 530490 363134
rect 530726 362898 530768 363134
rect 530448 362866 530768 362898
rect 561168 363454 561488 363486
rect 561168 363218 561210 363454
rect 561446 363218 561488 363454
rect 561168 363134 561488 363218
rect 561168 362898 561210 363134
rect 561446 362898 561488 363134
rect 561168 362866 561488 362898
rect 567234 352894 567854 388338
rect 567234 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 567854 352894
rect 567234 352574 567854 352658
rect 567234 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 567854 352574
rect 23568 345454 23888 345486
rect 23568 345218 23610 345454
rect 23846 345218 23888 345454
rect 23568 345134 23888 345218
rect 23568 344898 23610 345134
rect 23846 344898 23888 345134
rect 23568 344866 23888 344898
rect 54288 345454 54608 345486
rect 54288 345218 54330 345454
rect 54566 345218 54608 345454
rect 54288 345134 54608 345218
rect 54288 344898 54330 345134
rect 54566 344898 54608 345134
rect 54288 344866 54608 344898
rect 85008 345454 85328 345486
rect 85008 345218 85050 345454
rect 85286 345218 85328 345454
rect 85008 345134 85328 345218
rect 85008 344898 85050 345134
rect 85286 344898 85328 345134
rect 85008 344866 85328 344898
rect 115728 345454 116048 345486
rect 115728 345218 115770 345454
rect 116006 345218 116048 345454
rect 115728 345134 116048 345218
rect 115728 344898 115770 345134
rect 116006 344898 116048 345134
rect 115728 344866 116048 344898
rect 146448 345454 146768 345486
rect 146448 345218 146490 345454
rect 146726 345218 146768 345454
rect 146448 345134 146768 345218
rect 146448 344898 146490 345134
rect 146726 344898 146768 345134
rect 146448 344866 146768 344898
rect 177168 345454 177488 345486
rect 177168 345218 177210 345454
rect 177446 345218 177488 345454
rect 177168 345134 177488 345218
rect 177168 344898 177210 345134
rect 177446 344898 177488 345134
rect 177168 344866 177488 344898
rect 207888 345454 208208 345486
rect 207888 345218 207930 345454
rect 208166 345218 208208 345454
rect 207888 345134 208208 345218
rect 207888 344898 207930 345134
rect 208166 344898 208208 345134
rect 207888 344866 208208 344898
rect 238608 345454 238928 345486
rect 238608 345218 238650 345454
rect 238886 345218 238928 345454
rect 238608 345134 238928 345218
rect 238608 344898 238650 345134
rect 238886 344898 238928 345134
rect 238608 344866 238928 344898
rect 269328 345454 269648 345486
rect 269328 345218 269370 345454
rect 269606 345218 269648 345454
rect 269328 345134 269648 345218
rect 269328 344898 269370 345134
rect 269606 344898 269648 345134
rect 269328 344866 269648 344898
rect 300048 345454 300368 345486
rect 300048 345218 300090 345454
rect 300326 345218 300368 345454
rect 300048 345134 300368 345218
rect 300048 344898 300090 345134
rect 300326 344898 300368 345134
rect 300048 344866 300368 344898
rect 330768 345454 331088 345486
rect 330768 345218 330810 345454
rect 331046 345218 331088 345454
rect 330768 345134 331088 345218
rect 330768 344898 330810 345134
rect 331046 344898 331088 345134
rect 330768 344866 331088 344898
rect 361488 345454 361808 345486
rect 361488 345218 361530 345454
rect 361766 345218 361808 345454
rect 361488 345134 361808 345218
rect 361488 344898 361530 345134
rect 361766 344898 361808 345134
rect 361488 344866 361808 344898
rect 392208 345454 392528 345486
rect 392208 345218 392250 345454
rect 392486 345218 392528 345454
rect 392208 345134 392528 345218
rect 392208 344898 392250 345134
rect 392486 344898 392528 345134
rect 392208 344866 392528 344898
rect 422928 345454 423248 345486
rect 422928 345218 422970 345454
rect 423206 345218 423248 345454
rect 422928 345134 423248 345218
rect 422928 344898 422970 345134
rect 423206 344898 423248 345134
rect 422928 344866 423248 344898
rect 453648 345454 453968 345486
rect 453648 345218 453690 345454
rect 453926 345218 453968 345454
rect 453648 345134 453968 345218
rect 453648 344898 453690 345134
rect 453926 344898 453968 345134
rect 453648 344866 453968 344898
rect 484368 345454 484688 345486
rect 484368 345218 484410 345454
rect 484646 345218 484688 345454
rect 484368 345134 484688 345218
rect 484368 344898 484410 345134
rect 484646 344898 484688 345134
rect 484368 344866 484688 344898
rect 515088 345454 515408 345486
rect 515088 345218 515130 345454
rect 515366 345218 515408 345454
rect 515088 345134 515408 345218
rect 515088 344898 515130 345134
rect 515366 344898 515408 345134
rect 515088 344866 515408 344898
rect 545808 345454 546128 345486
rect 545808 345218 545850 345454
rect 546086 345218 546128 345454
rect 545808 345134 546128 345218
rect 545808 344898 545850 345134
rect 546086 344898 546128 345134
rect 545808 344866 546128 344898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect 8208 327454 8528 327486
rect 8208 327218 8250 327454
rect 8486 327218 8528 327454
rect 8208 327134 8528 327218
rect 8208 326898 8250 327134
rect 8486 326898 8528 327134
rect 8208 326866 8528 326898
rect 38928 327454 39248 327486
rect 38928 327218 38970 327454
rect 39206 327218 39248 327454
rect 38928 327134 39248 327218
rect 38928 326898 38970 327134
rect 39206 326898 39248 327134
rect 38928 326866 39248 326898
rect 69648 327454 69968 327486
rect 69648 327218 69690 327454
rect 69926 327218 69968 327454
rect 69648 327134 69968 327218
rect 69648 326898 69690 327134
rect 69926 326898 69968 327134
rect 69648 326866 69968 326898
rect 100368 327454 100688 327486
rect 100368 327218 100410 327454
rect 100646 327218 100688 327454
rect 100368 327134 100688 327218
rect 100368 326898 100410 327134
rect 100646 326898 100688 327134
rect 100368 326866 100688 326898
rect 131088 327454 131408 327486
rect 131088 327218 131130 327454
rect 131366 327218 131408 327454
rect 131088 327134 131408 327218
rect 131088 326898 131130 327134
rect 131366 326898 131408 327134
rect 131088 326866 131408 326898
rect 161808 327454 162128 327486
rect 161808 327218 161850 327454
rect 162086 327218 162128 327454
rect 161808 327134 162128 327218
rect 161808 326898 161850 327134
rect 162086 326898 162128 327134
rect 161808 326866 162128 326898
rect 192528 327454 192848 327486
rect 192528 327218 192570 327454
rect 192806 327218 192848 327454
rect 192528 327134 192848 327218
rect 192528 326898 192570 327134
rect 192806 326898 192848 327134
rect 192528 326866 192848 326898
rect 223248 327454 223568 327486
rect 223248 327218 223290 327454
rect 223526 327218 223568 327454
rect 223248 327134 223568 327218
rect 223248 326898 223290 327134
rect 223526 326898 223568 327134
rect 223248 326866 223568 326898
rect 253968 327454 254288 327486
rect 253968 327218 254010 327454
rect 254246 327218 254288 327454
rect 253968 327134 254288 327218
rect 253968 326898 254010 327134
rect 254246 326898 254288 327134
rect 253968 326866 254288 326898
rect 284688 327454 285008 327486
rect 284688 327218 284730 327454
rect 284966 327218 285008 327454
rect 284688 327134 285008 327218
rect 284688 326898 284730 327134
rect 284966 326898 285008 327134
rect 284688 326866 285008 326898
rect 315408 327454 315728 327486
rect 315408 327218 315450 327454
rect 315686 327218 315728 327454
rect 315408 327134 315728 327218
rect 315408 326898 315450 327134
rect 315686 326898 315728 327134
rect 315408 326866 315728 326898
rect 346128 327454 346448 327486
rect 346128 327218 346170 327454
rect 346406 327218 346448 327454
rect 346128 327134 346448 327218
rect 346128 326898 346170 327134
rect 346406 326898 346448 327134
rect 346128 326866 346448 326898
rect 376848 327454 377168 327486
rect 376848 327218 376890 327454
rect 377126 327218 377168 327454
rect 376848 327134 377168 327218
rect 376848 326898 376890 327134
rect 377126 326898 377168 327134
rect 376848 326866 377168 326898
rect 407568 327454 407888 327486
rect 407568 327218 407610 327454
rect 407846 327218 407888 327454
rect 407568 327134 407888 327218
rect 407568 326898 407610 327134
rect 407846 326898 407888 327134
rect 407568 326866 407888 326898
rect 438288 327454 438608 327486
rect 438288 327218 438330 327454
rect 438566 327218 438608 327454
rect 438288 327134 438608 327218
rect 438288 326898 438330 327134
rect 438566 326898 438608 327134
rect 438288 326866 438608 326898
rect 469008 327454 469328 327486
rect 469008 327218 469050 327454
rect 469286 327218 469328 327454
rect 469008 327134 469328 327218
rect 469008 326898 469050 327134
rect 469286 326898 469328 327134
rect 469008 326866 469328 326898
rect 499728 327454 500048 327486
rect 499728 327218 499770 327454
rect 500006 327218 500048 327454
rect 499728 327134 500048 327218
rect 499728 326898 499770 327134
rect 500006 326898 500048 327134
rect 499728 326866 500048 326898
rect 530448 327454 530768 327486
rect 530448 327218 530490 327454
rect 530726 327218 530768 327454
rect 530448 327134 530768 327218
rect 530448 326898 530490 327134
rect 530726 326898 530768 327134
rect 530448 326866 530768 326898
rect 561168 327454 561488 327486
rect 561168 327218 561210 327454
rect 561446 327218 561488 327454
rect 561168 327134 561488 327218
rect 561168 326898 561210 327134
rect 561446 326898 561488 327134
rect 561168 326866 561488 326898
rect 567234 316894 567854 352338
rect 567234 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 567854 316894
rect 567234 316574 567854 316658
rect 567234 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 567854 316574
rect 23568 309454 23888 309486
rect 23568 309218 23610 309454
rect 23846 309218 23888 309454
rect 23568 309134 23888 309218
rect 23568 308898 23610 309134
rect 23846 308898 23888 309134
rect 23568 308866 23888 308898
rect 54288 309454 54608 309486
rect 54288 309218 54330 309454
rect 54566 309218 54608 309454
rect 54288 309134 54608 309218
rect 54288 308898 54330 309134
rect 54566 308898 54608 309134
rect 54288 308866 54608 308898
rect 85008 309454 85328 309486
rect 85008 309218 85050 309454
rect 85286 309218 85328 309454
rect 85008 309134 85328 309218
rect 85008 308898 85050 309134
rect 85286 308898 85328 309134
rect 85008 308866 85328 308898
rect 115728 309454 116048 309486
rect 115728 309218 115770 309454
rect 116006 309218 116048 309454
rect 115728 309134 116048 309218
rect 115728 308898 115770 309134
rect 116006 308898 116048 309134
rect 115728 308866 116048 308898
rect 146448 309454 146768 309486
rect 146448 309218 146490 309454
rect 146726 309218 146768 309454
rect 146448 309134 146768 309218
rect 146448 308898 146490 309134
rect 146726 308898 146768 309134
rect 146448 308866 146768 308898
rect 177168 309454 177488 309486
rect 177168 309218 177210 309454
rect 177446 309218 177488 309454
rect 177168 309134 177488 309218
rect 177168 308898 177210 309134
rect 177446 308898 177488 309134
rect 177168 308866 177488 308898
rect 207888 309454 208208 309486
rect 207888 309218 207930 309454
rect 208166 309218 208208 309454
rect 207888 309134 208208 309218
rect 207888 308898 207930 309134
rect 208166 308898 208208 309134
rect 207888 308866 208208 308898
rect 238608 309454 238928 309486
rect 238608 309218 238650 309454
rect 238886 309218 238928 309454
rect 238608 309134 238928 309218
rect 238608 308898 238650 309134
rect 238886 308898 238928 309134
rect 238608 308866 238928 308898
rect 269328 309454 269648 309486
rect 269328 309218 269370 309454
rect 269606 309218 269648 309454
rect 269328 309134 269648 309218
rect 269328 308898 269370 309134
rect 269606 308898 269648 309134
rect 269328 308866 269648 308898
rect 300048 309454 300368 309486
rect 300048 309218 300090 309454
rect 300326 309218 300368 309454
rect 300048 309134 300368 309218
rect 300048 308898 300090 309134
rect 300326 308898 300368 309134
rect 300048 308866 300368 308898
rect 330768 309454 331088 309486
rect 330768 309218 330810 309454
rect 331046 309218 331088 309454
rect 330768 309134 331088 309218
rect 330768 308898 330810 309134
rect 331046 308898 331088 309134
rect 330768 308866 331088 308898
rect 361488 309454 361808 309486
rect 361488 309218 361530 309454
rect 361766 309218 361808 309454
rect 361488 309134 361808 309218
rect 361488 308898 361530 309134
rect 361766 308898 361808 309134
rect 361488 308866 361808 308898
rect 392208 309454 392528 309486
rect 392208 309218 392250 309454
rect 392486 309218 392528 309454
rect 392208 309134 392528 309218
rect 392208 308898 392250 309134
rect 392486 308898 392528 309134
rect 392208 308866 392528 308898
rect 422928 309454 423248 309486
rect 422928 309218 422970 309454
rect 423206 309218 423248 309454
rect 422928 309134 423248 309218
rect 422928 308898 422970 309134
rect 423206 308898 423248 309134
rect 422928 308866 423248 308898
rect 453648 309454 453968 309486
rect 453648 309218 453690 309454
rect 453926 309218 453968 309454
rect 453648 309134 453968 309218
rect 453648 308898 453690 309134
rect 453926 308898 453968 309134
rect 453648 308866 453968 308898
rect 484368 309454 484688 309486
rect 484368 309218 484410 309454
rect 484646 309218 484688 309454
rect 484368 309134 484688 309218
rect 484368 308898 484410 309134
rect 484646 308898 484688 309134
rect 484368 308866 484688 308898
rect 515088 309454 515408 309486
rect 515088 309218 515130 309454
rect 515366 309218 515408 309454
rect 515088 309134 515408 309218
rect 515088 308898 515130 309134
rect 515366 308898 515408 309134
rect 515088 308866 515408 308898
rect 545808 309454 546128 309486
rect 545808 309218 545850 309454
rect 546086 309218 546128 309454
rect 545808 309134 546128 309218
rect 545808 308898 545850 309134
rect 546086 308898 546128 309134
rect 545808 308866 546128 308898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect 8208 291454 8528 291486
rect 8208 291218 8250 291454
rect 8486 291218 8528 291454
rect 8208 291134 8528 291218
rect 8208 290898 8250 291134
rect 8486 290898 8528 291134
rect 8208 290866 8528 290898
rect 38928 291454 39248 291486
rect 38928 291218 38970 291454
rect 39206 291218 39248 291454
rect 38928 291134 39248 291218
rect 38928 290898 38970 291134
rect 39206 290898 39248 291134
rect 38928 290866 39248 290898
rect 69648 291454 69968 291486
rect 69648 291218 69690 291454
rect 69926 291218 69968 291454
rect 69648 291134 69968 291218
rect 69648 290898 69690 291134
rect 69926 290898 69968 291134
rect 69648 290866 69968 290898
rect 100368 291454 100688 291486
rect 100368 291218 100410 291454
rect 100646 291218 100688 291454
rect 100368 291134 100688 291218
rect 100368 290898 100410 291134
rect 100646 290898 100688 291134
rect 100368 290866 100688 290898
rect 131088 291454 131408 291486
rect 131088 291218 131130 291454
rect 131366 291218 131408 291454
rect 131088 291134 131408 291218
rect 131088 290898 131130 291134
rect 131366 290898 131408 291134
rect 131088 290866 131408 290898
rect 161808 291454 162128 291486
rect 161808 291218 161850 291454
rect 162086 291218 162128 291454
rect 161808 291134 162128 291218
rect 161808 290898 161850 291134
rect 162086 290898 162128 291134
rect 161808 290866 162128 290898
rect 192528 291454 192848 291486
rect 192528 291218 192570 291454
rect 192806 291218 192848 291454
rect 192528 291134 192848 291218
rect 192528 290898 192570 291134
rect 192806 290898 192848 291134
rect 192528 290866 192848 290898
rect 223248 291454 223568 291486
rect 223248 291218 223290 291454
rect 223526 291218 223568 291454
rect 223248 291134 223568 291218
rect 223248 290898 223290 291134
rect 223526 290898 223568 291134
rect 223248 290866 223568 290898
rect 253968 291454 254288 291486
rect 253968 291218 254010 291454
rect 254246 291218 254288 291454
rect 253968 291134 254288 291218
rect 253968 290898 254010 291134
rect 254246 290898 254288 291134
rect 253968 290866 254288 290898
rect 284688 291454 285008 291486
rect 284688 291218 284730 291454
rect 284966 291218 285008 291454
rect 284688 291134 285008 291218
rect 284688 290898 284730 291134
rect 284966 290898 285008 291134
rect 284688 290866 285008 290898
rect 315408 291454 315728 291486
rect 315408 291218 315450 291454
rect 315686 291218 315728 291454
rect 315408 291134 315728 291218
rect 315408 290898 315450 291134
rect 315686 290898 315728 291134
rect 315408 290866 315728 290898
rect 346128 291454 346448 291486
rect 346128 291218 346170 291454
rect 346406 291218 346448 291454
rect 346128 291134 346448 291218
rect 346128 290898 346170 291134
rect 346406 290898 346448 291134
rect 346128 290866 346448 290898
rect 376848 291454 377168 291486
rect 376848 291218 376890 291454
rect 377126 291218 377168 291454
rect 376848 291134 377168 291218
rect 376848 290898 376890 291134
rect 377126 290898 377168 291134
rect 376848 290866 377168 290898
rect 407568 291454 407888 291486
rect 407568 291218 407610 291454
rect 407846 291218 407888 291454
rect 407568 291134 407888 291218
rect 407568 290898 407610 291134
rect 407846 290898 407888 291134
rect 407568 290866 407888 290898
rect 438288 291454 438608 291486
rect 438288 291218 438330 291454
rect 438566 291218 438608 291454
rect 438288 291134 438608 291218
rect 438288 290898 438330 291134
rect 438566 290898 438608 291134
rect 438288 290866 438608 290898
rect 469008 291454 469328 291486
rect 469008 291218 469050 291454
rect 469286 291218 469328 291454
rect 469008 291134 469328 291218
rect 469008 290898 469050 291134
rect 469286 290898 469328 291134
rect 469008 290866 469328 290898
rect 499728 291454 500048 291486
rect 499728 291218 499770 291454
rect 500006 291218 500048 291454
rect 499728 291134 500048 291218
rect 499728 290898 499770 291134
rect 500006 290898 500048 291134
rect 499728 290866 500048 290898
rect 530448 291454 530768 291486
rect 530448 291218 530490 291454
rect 530726 291218 530768 291454
rect 530448 291134 530768 291218
rect 530448 290898 530490 291134
rect 530726 290898 530768 291134
rect 530448 290866 530768 290898
rect 561168 291454 561488 291486
rect 561168 291218 561210 291454
rect 561446 291218 561488 291454
rect 561168 291134 561488 291218
rect 561168 290898 561210 291134
rect 561446 290898 561488 291134
rect 561168 290866 561488 290898
rect 567234 280894 567854 316338
rect 567234 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 567854 280894
rect 567234 280574 567854 280658
rect 567234 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 567854 280574
rect 23568 273454 23888 273486
rect 23568 273218 23610 273454
rect 23846 273218 23888 273454
rect 23568 273134 23888 273218
rect 23568 272898 23610 273134
rect 23846 272898 23888 273134
rect 23568 272866 23888 272898
rect 54288 273454 54608 273486
rect 54288 273218 54330 273454
rect 54566 273218 54608 273454
rect 54288 273134 54608 273218
rect 54288 272898 54330 273134
rect 54566 272898 54608 273134
rect 54288 272866 54608 272898
rect 85008 273454 85328 273486
rect 85008 273218 85050 273454
rect 85286 273218 85328 273454
rect 85008 273134 85328 273218
rect 85008 272898 85050 273134
rect 85286 272898 85328 273134
rect 85008 272866 85328 272898
rect 115728 273454 116048 273486
rect 115728 273218 115770 273454
rect 116006 273218 116048 273454
rect 115728 273134 116048 273218
rect 115728 272898 115770 273134
rect 116006 272898 116048 273134
rect 115728 272866 116048 272898
rect 146448 273454 146768 273486
rect 146448 273218 146490 273454
rect 146726 273218 146768 273454
rect 146448 273134 146768 273218
rect 146448 272898 146490 273134
rect 146726 272898 146768 273134
rect 146448 272866 146768 272898
rect 177168 273454 177488 273486
rect 177168 273218 177210 273454
rect 177446 273218 177488 273454
rect 177168 273134 177488 273218
rect 177168 272898 177210 273134
rect 177446 272898 177488 273134
rect 177168 272866 177488 272898
rect 207888 273454 208208 273486
rect 207888 273218 207930 273454
rect 208166 273218 208208 273454
rect 207888 273134 208208 273218
rect 207888 272898 207930 273134
rect 208166 272898 208208 273134
rect 207888 272866 208208 272898
rect 238608 273454 238928 273486
rect 238608 273218 238650 273454
rect 238886 273218 238928 273454
rect 238608 273134 238928 273218
rect 238608 272898 238650 273134
rect 238886 272898 238928 273134
rect 238608 272866 238928 272898
rect 269328 273454 269648 273486
rect 269328 273218 269370 273454
rect 269606 273218 269648 273454
rect 269328 273134 269648 273218
rect 269328 272898 269370 273134
rect 269606 272898 269648 273134
rect 269328 272866 269648 272898
rect 300048 273454 300368 273486
rect 300048 273218 300090 273454
rect 300326 273218 300368 273454
rect 300048 273134 300368 273218
rect 300048 272898 300090 273134
rect 300326 272898 300368 273134
rect 300048 272866 300368 272898
rect 330768 273454 331088 273486
rect 330768 273218 330810 273454
rect 331046 273218 331088 273454
rect 330768 273134 331088 273218
rect 330768 272898 330810 273134
rect 331046 272898 331088 273134
rect 330768 272866 331088 272898
rect 361488 273454 361808 273486
rect 361488 273218 361530 273454
rect 361766 273218 361808 273454
rect 361488 273134 361808 273218
rect 361488 272898 361530 273134
rect 361766 272898 361808 273134
rect 361488 272866 361808 272898
rect 392208 273454 392528 273486
rect 392208 273218 392250 273454
rect 392486 273218 392528 273454
rect 392208 273134 392528 273218
rect 392208 272898 392250 273134
rect 392486 272898 392528 273134
rect 392208 272866 392528 272898
rect 422928 273454 423248 273486
rect 422928 273218 422970 273454
rect 423206 273218 423248 273454
rect 422928 273134 423248 273218
rect 422928 272898 422970 273134
rect 423206 272898 423248 273134
rect 422928 272866 423248 272898
rect 453648 273454 453968 273486
rect 453648 273218 453690 273454
rect 453926 273218 453968 273454
rect 453648 273134 453968 273218
rect 453648 272898 453690 273134
rect 453926 272898 453968 273134
rect 453648 272866 453968 272898
rect 484368 273454 484688 273486
rect 484368 273218 484410 273454
rect 484646 273218 484688 273454
rect 484368 273134 484688 273218
rect 484368 272898 484410 273134
rect 484646 272898 484688 273134
rect 484368 272866 484688 272898
rect 515088 273454 515408 273486
rect 515088 273218 515130 273454
rect 515366 273218 515408 273454
rect 515088 273134 515408 273218
rect 515088 272898 515130 273134
rect 515366 272898 515408 273134
rect 515088 272866 515408 272898
rect 545808 273454 546128 273486
rect 545808 273218 545850 273454
rect 546086 273218 546128 273454
rect 545808 273134 546128 273218
rect 545808 272898 545850 273134
rect 546086 272898 546128 273134
rect 545808 272866 546128 272898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect 8208 255454 8528 255486
rect 8208 255218 8250 255454
rect 8486 255218 8528 255454
rect 8208 255134 8528 255218
rect 8208 254898 8250 255134
rect 8486 254898 8528 255134
rect 8208 254866 8528 254898
rect 38928 255454 39248 255486
rect 38928 255218 38970 255454
rect 39206 255218 39248 255454
rect 38928 255134 39248 255218
rect 38928 254898 38970 255134
rect 39206 254898 39248 255134
rect 38928 254866 39248 254898
rect 69648 255454 69968 255486
rect 69648 255218 69690 255454
rect 69926 255218 69968 255454
rect 69648 255134 69968 255218
rect 69648 254898 69690 255134
rect 69926 254898 69968 255134
rect 69648 254866 69968 254898
rect 100368 255454 100688 255486
rect 100368 255218 100410 255454
rect 100646 255218 100688 255454
rect 100368 255134 100688 255218
rect 100368 254898 100410 255134
rect 100646 254898 100688 255134
rect 100368 254866 100688 254898
rect 131088 255454 131408 255486
rect 131088 255218 131130 255454
rect 131366 255218 131408 255454
rect 131088 255134 131408 255218
rect 131088 254898 131130 255134
rect 131366 254898 131408 255134
rect 131088 254866 131408 254898
rect 161808 255454 162128 255486
rect 161808 255218 161850 255454
rect 162086 255218 162128 255454
rect 161808 255134 162128 255218
rect 161808 254898 161850 255134
rect 162086 254898 162128 255134
rect 161808 254866 162128 254898
rect 192528 255454 192848 255486
rect 192528 255218 192570 255454
rect 192806 255218 192848 255454
rect 192528 255134 192848 255218
rect 192528 254898 192570 255134
rect 192806 254898 192848 255134
rect 192528 254866 192848 254898
rect 223248 255454 223568 255486
rect 223248 255218 223290 255454
rect 223526 255218 223568 255454
rect 223248 255134 223568 255218
rect 223248 254898 223290 255134
rect 223526 254898 223568 255134
rect 223248 254866 223568 254898
rect 253968 255454 254288 255486
rect 253968 255218 254010 255454
rect 254246 255218 254288 255454
rect 253968 255134 254288 255218
rect 253968 254898 254010 255134
rect 254246 254898 254288 255134
rect 253968 254866 254288 254898
rect 284688 255454 285008 255486
rect 284688 255218 284730 255454
rect 284966 255218 285008 255454
rect 284688 255134 285008 255218
rect 284688 254898 284730 255134
rect 284966 254898 285008 255134
rect 284688 254866 285008 254898
rect 315408 255454 315728 255486
rect 315408 255218 315450 255454
rect 315686 255218 315728 255454
rect 315408 255134 315728 255218
rect 315408 254898 315450 255134
rect 315686 254898 315728 255134
rect 315408 254866 315728 254898
rect 346128 255454 346448 255486
rect 346128 255218 346170 255454
rect 346406 255218 346448 255454
rect 346128 255134 346448 255218
rect 346128 254898 346170 255134
rect 346406 254898 346448 255134
rect 346128 254866 346448 254898
rect 376848 255454 377168 255486
rect 376848 255218 376890 255454
rect 377126 255218 377168 255454
rect 376848 255134 377168 255218
rect 376848 254898 376890 255134
rect 377126 254898 377168 255134
rect 376848 254866 377168 254898
rect 407568 255454 407888 255486
rect 407568 255218 407610 255454
rect 407846 255218 407888 255454
rect 407568 255134 407888 255218
rect 407568 254898 407610 255134
rect 407846 254898 407888 255134
rect 407568 254866 407888 254898
rect 438288 255454 438608 255486
rect 438288 255218 438330 255454
rect 438566 255218 438608 255454
rect 438288 255134 438608 255218
rect 438288 254898 438330 255134
rect 438566 254898 438608 255134
rect 438288 254866 438608 254898
rect 469008 255454 469328 255486
rect 469008 255218 469050 255454
rect 469286 255218 469328 255454
rect 469008 255134 469328 255218
rect 469008 254898 469050 255134
rect 469286 254898 469328 255134
rect 469008 254866 469328 254898
rect 499728 255454 500048 255486
rect 499728 255218 499770 255454
rect 500006 255218 500048 255454
rect 499728 255134 500048 255218
rect 499728 254898 499770 255134
rect 500006 254898 500048 255134
rect 499728 254866 500048 254898
rect 530448 255454 530768 255486
rect 530448 255218 530490 255454
rect 530726 255218 530768 255454
rect 530448 255134 530768 255218
rect 530448 254898 530490 255134
rect 530726 254898 530768 255134
rect 530448 254866 530768 254898
rect 561168 255454 561488 255486
rect 561168 255218 561210 255454
rect 561446 255218 561488 255454
rect 561168 255134 561488 255218
rect 561168 254898 561210 255134
rect 561446 254898 561488 255134
rect 561168 254866 561488 254898
rect 567234 244894 567854 280338
rect 567234 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 567854 244894
rect 567234 244574 567854 244658
rect 567234 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 567854 244574
rect 23568 237454 23888 237486
rect 23568 237218 23610 237454
rect 23846 237218 23888 237454
rect 23568 237134 23888 237218
rect 23568 236898 23610 237134
rect 23846 236898 23888 237134
rect 23568 236866 23888 236898
rect 54288 237454 54608 237486
rect 54288 237218 54330 237454
rect 54566 237218 54608 237454
rect 54288 237134 54608 237218
rect 54288 236898 54330 237134
rect 54566 236898 54608 237134
rect 54288 236866 54608 236898
rect 85008 237454 85328 237486
rect 85008 237218 85050 237454
rect 85286 237218 85328 237454
rect 85008 237134 85328 237218
rect 85008 236898 85050 237134
rect 85286 236898 85328 237134
rect 85008 236866 85328 236898
rect 115728 237454 116048 237486
rect 115728 237218 115770 237454
rect 116006 237218 116048 237454
rect 115728 237134 116048 237218
rect 115728 236898 115770 237134
rect 116006 236898 116048 237134
rect 115728 236866 116048 236898
rect 146448 237454 146768 237486
rect 146448 237218 146490 237454
rect 146726 237218 146768 237454
rect 146448 237134 146768 237218
rect 146448 236898 146490 237134
rect 146726 236898 146768 237134
rect 146448 236866 146768 236898
rect 177168 237454 177488 237486
rect 177168 237218 177210 237454
rect 177446 237218 177488 237454
rect 177168 237134 177488 237218
rect 177168 236898 177210 237134
rect 177446 236898 177488 237134
rect 177168 236866 177488 236898
rect 207888 237454 208208 237486
rect 207888 237218 207930 237454
rect 208166 237218 208208 237454
rect 207888 237134 208208 237218
rect 207888 236898 207930 237134
rect 208166 236898 208208 237134
rect 207888 236866 208208 236898
rect 238608 237454 238928 237486
rect 238608 237218 238650 237454
rect 238886 237218 238928 237454
rect 238608 237134 238928 237218
rect 238608 236898 238650 237134
rect 238886 236898 238928 237134
rect 238608 236866 238928 236898
rect 269328 237454 269648 237486
rect 269328 237218 269370 237454
rect 269606 237218 269648 237454
rect 269328 237134 269648 237218
rect 269328 236898 269370 237134
rect 269606 236898 269648 237134
rect 269328 236866 269648 236898
rect 300048 237454 300368 237486
rect 300048 237218 300090 237454
rect 300326 237218 300368 237454
rect 300048 237134 300368 237218
rect 300048 236898 300090 237134
rect 300326 236898 300368 237134
rect 300048 236866 300368 236898
rect 330768 237454 331088 237486
rect 330768 237218 330810 237454
rect 331046 237218 331088 237454
rect 330768 237134 331088 237218
rect 330768 236898 330810 237134
rect 331046 236898 331088 237134
rect 330768 236866 331088 236898
rect 361488 237454 361808 237486
rect 361488 237218 361530 237454
rect 361766 237218 361808 237454
rect 361488 237134 361808 237218
rect 361488 236898 361530 237134
rect 361766 236898 361808 237134
rect 361488 236866 361808 236898
rect 392208 237454 392528 237486
rect 392208 237218 392250 237454
rect 392486 237218 392528 237454
rect 392208 237134 392528 237218
rect 392208 236898 392250 237134
rect 392486 236898 392528 237134
rect 392208 236866 392528 236898
rect 422928 237454 423248 237486
rect 422928 237218 422970 237454
rect 423206 237218 423248 237454
rect 422928 237134 423248 237218
rect 422928 236898 422970 237134
rect 423206 236898 423248 237134
rect 422928 236866 423248 236898
rect 453648 237454 453968 237486
rect 453648 237218 453690 237454
rect 453926 237218 453968 237454
rect 453648 237134 453968 237218
rect 453648 236898 453690 237134
rect 453926 236898 453968 237134
rect 453648 236866 453968 236898
rect 484368 237454 484688 237486
rect 484368 237218 484410 237454
rect 484646 237218 484688 237454
rect 484368 237134 484688 237218
rect 484368 236898 484410 237134
rect 484646 236898 484688 237134
rect 484368 236866 484688 236898
rect 515088 237454 515408 237486
rect 515088 237218 515130 237454
rect 515366 237218 515408 237454
rect 515088 237134 515408 237218
rect 515088 236898 515130 237134
rect 515366 236898 515408 237134
rect 515088 236866 515408 236898
rect 545808 237454 546128 237486
rect 545808 237218 545850 237454
rect 546086 237218 546128 237454
rect 545808 237134 546128 237218
rect 545808 236898 545850 237134
rect 546086 236898 546128 237134
rect 545808 236866 546128 236898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect 8208 219454 8528 219486
rect 8208 219218 8250 219454
rect 8486 219218 8528 219454
rect 8208 219134 8528 219218
rect 8208 218898 8250 219134
rect 8486 218898 8528 219134
rect 8208 218866 8528 218898
rect 38928 219454 39248 219486
rect 38928 219218 38970 219454
rect 39206 219218 39248 219454
rect 38928 219134 39248 219218
rect 38928 218898 38970 219134
rect 39206 218898 39248 219134
rect 38928 218866 39248 218898
rect 69648 219454 69968 219486
rect 69648 219218 69690 219454
rect 69926 219218 69968 219454
rect 69648 219134 69968 219218
rect 69648 218898 69690 219134
rect 69926 218898 69968 219134
rect 69648 218866 69968 218898
rect 100368 219454 100688 219486
rect 100368 219218 100410 219454
rect 100646 219218 100688 219454
rect 100368 219134 100688 219218
rect 100368 218898 100410 219134
rect 100646 218898 100688 219134
rect 100368 218866 100688 218898
rect 131088 219454 131408 219486
rect 131088 219218 131130 219454
rect 131366 219218 131408 219454
rect 131088 219134 131408 219218
rect 131088 218898 131130 219134
rect 131366 218898 131408 219134
rect 131088 218866 131408 218898
rect 161808 219454 162128 219486
rect 161808 219218 161850 219454
rect 162086 219218 162128 219454
rect 161808 219134 162128 219218
rect 161808 218898 161850 219134
rect 162086 218898 162128 219134
rect 161808 218866 162128 218898
rect 192528 219454 192848 219486
rect 192528 219218 192570 219454
rect 192806 219218 192848 219454
rect 192528 219134 192848 219218
rect 192528 218898 192570 219134
rect 192806 218898 192848 219134
rect 192528 218866 192848 218898
rect 223248 219454 223568 219486
rect 223248 219218 223290 219454
rect 223526 219218 223568 219454
rect 223248 219134 223568 219218
rect 223248 218898 223290 219134
rect 223526 218898 223568 219134
rect 223248 218866 223568 218898
rect 253968 219454 254288 219486
rect 253968 219218 254010 219454
rect 254246 219218 254288 219454
rect 253968 219134 254288 219218
rect 253968 218898 254010 219134
rect 254246 218898 254288 219134
rect 253968 218866 254288 218898
rect 284688 219454 285008 219486
rect 284688 219218 284730 219454
rect 284966 219218 285008 219454
rect 284688 219134 285008 219218
rect 284688 218898 284730 219134
rect 284966 218898 285008 219134
rect 284688 218866 285008 218898
rect 315408 219454 315728 219486
rect 315408 219218 315450 219454
rect 315686 219218 315728 219454
rect 315408 219134 315728 219218
rect 315408 218898 315450 219134
rect 315686 218898 315728 219134
rect 315408 218866 315728 218898
rect 346128 219454 346448 219486
rect 346128 219218 346170 219454
rect 346406 219218 346448 219454
rect 346128 219134 346448 219218
rect 346128 218898 346170 219134
rect 346406 218898 346448 219134
rect 346128 218866 346448 218898
rect 376848 219454 377168 219486
rect 376848 219218 376890 219454
rect 377126 219218 377168 219454
rect 376848 219134 377168 219218
rect 376848 218898 376890 219134
rect 377126 218898 377168 219134
rect 376848 218866 377168 218898
rect 407568 219454 407888 219486
rect 407568 219218 407610 219454
rect 407846 219218 407888 219454
rect 407568 219134 407888 219218
rect 407568 218898 407610 219134
rect 407846 218898 407888 219134
rect 407568 218866 407888 218898
rect 438288 219454 438608 219486
rect 438288 219218 438330 219454
rect 438566 219218 438608 219454
rect 438288 219134 438608 219218
rect 438288 218898 438330 219134
rect 438566 218898 438608 219134
rect 438288 218866 438608 218898
rect 469008 219454 469328 219486
rect 469008 219218 469050 219454
rect 469286 219218 469328 219454
rect 469008 219134 469328 219218
rect 469008 218898 469050 219134
rect 469286 218898 469328 219134
rect 469008 218866 469328 218898
rect 499728 219454 500048 219486
rect 499728 219218 499770 219454
rect 500006 219218 500048 219454
rect 499728 219134 500048 219218
rect 499728 218898 499770 219134
rect 500006 218898 500048 219134
rect 499728 218866 500048 218898
rect 530448 219454 530768 219486
rect 530448 219218 530490 219454
rect 530726 219218 530768 219454
rect 530448 219134 530768 219218
rect 530448 218898 530490 219134
rect 530726 218898 530768 219134
rect 530448 218866 530768 218898
rect 561168 219454 561488 219486
rect 561168 219218 561210 219454
rect 561446 219218 561488 219454
rect 561168 219134 561488 219218
rect 561168 218898 561210 219134
rect 561446 218898 561488 219134
rect 561168 218866 561488 218898
rect 567234 208894 567854 244338
rect 567234 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 567854 208894
rect 567234 208574 567854 208658
rect 567234 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 567854 208574
rect 23568 201454 23888 201486
rect 23568 201218 23610 201454
rect 23846 201218 23888 201454
rect 23568 201134 23888 201218
rect 23568 200898 23610 201134
rect 23846 200898 23888 201134
rect 23568 200866 23888 200898
rect 54288 201454 54608 201486
rect 54288 201218 54330 201454
rect 54566 201218 54608 201454
rect 54288 201134 54608 201218
rect 54288 200898 54330 201134
rect 54566 200898 54608 201134
rect 54288 200866 54608 200898
rect 85008 201454 85328 201486
rect 85008 201218 85050 201454
rect 85286 201218 85328 201454
rect 85008 201134 85328 201218
rect 85008 200898 85050 201134
rect 85286 200898 85328 201134
rect 85008 200866 85328 200898
rect 115728 201454 116048 201486
rect 115728 201218 115770 201454
rect 116006 201218 116048 201454
rect 115728 201134 116048 201218
rect 115728 200898 115770 201134
rect 116006 200898 116048 201134
rect 115728 200866 116048 200898
rect 146448 201454 146768 201486
rect 146448 201218 146490 201454
rect 146726 201218 146768 201454
rect 146448 201134 146768 201218
rect 146448 200898 146490 201134
rect 146726 200898 146768 201134
rect 146448 200866 146768 200898
rect 177168 201454 177488 201486
rect 177168 201218 177210 201454
rect 177446 201218 177488 201454
rect 177168 201134 177488 201218
rect 177168 200898 177210 201134
rect 177446 200898 177488 201134
rect 177168 200866 177488 200898
rect 207888 201454 208208 201486
rect 207888 201218 207930 201454
rect 208166 201218 208208 201454
rect 207888 201134 208208 201218
rect 207888 200898 207930 201134
rect 208166 200898 208208 201134
rect 207888 200866 208208 200898
rect 238608 201454 238928 201486
rect 238608 201218 238650 201454
rect 238886 201218 238928 201454
rect 238608 201134 238928 201218
rect 238608 200898 238650 201134
rect 238886 200898 238928 201134
rect 238608 200866 238928 200898
rect 269328 201454 269648 201486
rect 269328 201218 269370 201454
rect 269606 201218 269648 201454
rect 269328 201134 269648 201218
rect 269328 200898 269370 201134
rect 269606 200898 269648 201134
rect 269328 200866 269648 200898
rect 300048 201454 300368 201486
rect 300048 201218 300090 201454
rect 300326 201218 300368 201454
rect 300048 201134 300368 201218
rect 300048 200898 300090 201134
rect 300326 200898 300368 201134
rect 300048 200866 300368 200898
rect 330768 201454 331088 201486
rect 330768 201218 330810 201454
rect 331046 201218 331088 201454
rect 330768 201134 331088 201218
rect 330768 200898 330810 201134
rect 331046 200898 331088 201134
rect 330768 200866 331088 200898
rect 361488 201454 361808 201486
rect 361488 201218 361530 201454
rect 361766 201218 361808 201454
rect 361488 201134 361808 201218
rect 361488 200898 361530 201134
rect 361766 200898 361808 201134
rect 361488 200866 361808 200898
rect 392208 201454 392528 201486
rect 392208 201218 392250 201454
rect 392486 201218 392528 201454
rect 392208 201134 392528 201218
rect 392208 200898 392250 201134
rect 392486 200898 392528 201134
rect 392208 200866 392528 200898
rect 422928 201454 423248 201486
rect 422928 201218 422970 201454
rect 423206 201218 423248 201454
rect 422928 201134 423248 201218
rect 422928 200898 422970 201134
rect 423206 200898 423248 201134
rect 422928 200866 423248 200898
rect 453648 201454 453968 201486
rect 453648 201218 453690 201454
rect 453926 201218 453968 201454
rect 453648 201134 453968 201218
rect 453648 200898 453690 201134
rect 453926 200898 453968 201134
rect 453648 200866 453968 200898
rect 484368 201454 484688 201486
rect 484368 201218 484410 201454
rect 484646 201218 484688 201454
rect 484368 201134 484688 201218
rect 484368 200898 484410 201134
rect 484646 200898 484688 201134
rect 484368 200866 484688 200898
rect 515088 201454 515408 201486
rect 515088 201218 515130 201454
rect 515366 201218 515408 201454
rect 515088 201134 515408 201218
rect 515088 200898 515130 201134
rect 515366 200898 515408 201134
rect 515088 200866 515408 200898
rect 545808 201454 546128 201486
rect 545808 201218 545850 201454
rect 546086 201218 546128 201454
rect 545808 201134 546128 201218
rect 545808 200898 545850 201134
rect 546086 200898 546128 201134
rect 545808 200866 546128 200898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect 8208 183454 8528 183486
rect 8208 183218 8250 183454
rect 8486 183218 8528 183454
rect 8208 183134 8528 183218
rect 8208 182898 8250 183134
rect 8486 182898 8528 183134
rect 8208 182866 8528 182898
rect 38928 183454 39248 183486
rect 38928 183218 38970 183454
rect 39206 183218 39248 183454
rect 38928 183134 39248 183218
rect 38928 182898 38970 183134
rect 39206 182898 39248 183134
rect 38928 182866 39248 182898
rect 69648 183454 69968 183486
rect 69648 183218 69690 183454
rect 69926 183218 69968 183454
rect 69648 183134 69968 183218
rect 69648 182898 69690 183134
rect 69926 182898 69968 183134
rect 69648 182866 69968 182898
rect 100368 183454 100688 183486
rect 100368 183218 100410 183454
rect 100646 183218 100688 183454
rect 100368 183134 100688 183218
rect 100368 182898 100410 183134
rect 100646 182898 100688 183134
rect 100368 182866 100688 182898
rect 131088 183454 131408 183486
rect 131088 183218 131130 183454
rect 131366 183218 131408 183454
rect 131088 183134 131408 183218
rect 131088 182898 131130 183134
rect 131366 182898 131408 183134
rect 131088 182866 131408 182898
rect 161808 183454 162128 183486
rect 161808 183218 161850 183454
rect 162086 183218 162128 183454
rect 161808 183134 162128 183218
rect 161808 182898 161850 183134
rect 162086 182898 162128 183134
rect 161808 182866 162128 182898
rect 192528 183454 192848 183486
rect 192528 183218 192570 183454
rect 192806 183218 192848 183454
rect 192528 183134 192848 183218
rect 192528 182898 192570 183134
rect 192806 182898 192848 183134
rect 192528 182866 192848 182898
rect 223248 183454 223568 183486
rect 223248 183218 223290 183454
rect 223526 183218 223568 183454
rect 223248 183134 223568 183218
rect 223248 182898 223290 183134
rect 223526 182898 223568 183134
rect 223248 182866 223568 182898
rect 253968 183454 254288 183486
rect 253968 183218 254010 183454
rect 254246 183218 254288 183454
rect 253968 183134 254288 183218
rect 253968 182898 254010 183134
rect 254246 182898 254288 183134
rect 253968 182866 254288 182898
rect 284688 183454 285008 183486
rect 284688 183218 284730 183454
rect 284966 183218 285008 183454
rect 284688 183134 285008 183218
rect 284688 182898 284730 183134
rect 284966 182898 285008 183134
rect 284688 182866 285008 182898
rect 315408 183454 315728 183486
rect 315408 183218 315450 183454
rect 315686 183218 315728 183454
rect 315408 183134 315728 183218
rect 315408 182898 315450 183134
rect 315686 182898 315728 183134
rect 315408 182866 315728 182898
rect 346128 183454 346448 183486
rect 346128 183218 346170 183454
rect 346406 183218 346448 183454
rect 346128 183134 346448 183218
rect 346128 182898 346170 183134
rect 346406 182898 346448 183134
rect 346128 182866 346448 182898
rect 376848 183454 377168 183486
rect 376848 183218 376890 183454
rect 377126 183218 377168 183454
rect 376848 183134 377168 183218
rect 376848 182898 376890 183134
rect 377126 182898 377168 183134
rect 376848 182866 377168 182898
rect 407568 183454 407888 183486
rect 407568 183218 407610 183454
rect 407846 183218 407888 183454
rect 407568 183134 407888 183218
rect 407568 182898 407610 183134
rect 407846 182898 407888 183134
rect 407568 182866 407888 182898
rect 438288 183454 438608 183486
rect 438288 183218 438330 183454
rect 438566 183218 438608 183454
rect 438288 183134 438608 183218
rect 438288 182898 438330 183134
rect 438566 182898 438608 183134
rect 438288 182866 438608 182898
rect 469008 183454 469328 183486
rect 469008 183218 469050 183454
rect 469286 183218 469328 183454
rect 469008 183134 469328 183218
rect 469008 182898 469050 183134
rect 469286 182898 469328 183134
rect 469008 182866 469328 182898
rect 499728 183454 500048 183486
rect 499728 183218 499770 183454
rect 500006 183218 500048 183454
rect 499728 183134 500048 183218
rect 499728 182898 499770 183134
rect 500006 182898 500048 183134
rect 499728 182866 500048 182898
rect 530448 183454 530768 183486
rect 530448 183218 530490 183454
rect 530726 183218 530768 183454
rect 530448 183134 530768 183218
rect 530448 182898 530490 183134
rect 530726 182898 530768 183134
rect 530448 182866 530768 182898
rect 561168 183454 561488 183486
rect 561168 183218 561210 183454
rect 561446 183218 561488 183454
rect 561168 183134 561488 183218
rect 561168 182898 561210 183134
rect 561446 182898 561488 183134
rect 561168 182866 561488 182898
rect 567234 172894 567854 208338
rect 567234 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 567854 172894
rect 567234 172574 567854 172658
rect 567234 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 567854 172574
rect 23568 165454 23888 165486
rect 23568 165218 23610 165454
rect 23846 165218 23888 165454
rect 23568 165134 23888 165218
rect 23568 164898 23610 165134
rect 23846 164898 23888 165134
rect 23568 164866 23888 164898
rect 54288 165454 54608 165486
rect 54288 165218 54330 165454
rect 54566 165218 54608 165454
rect 54288 165134 54608 165218
rect 54288 164898 54330 165134
rect 54566 164898 54608 165134
rect 54288 164866 54608 164898
rect 85008 165454 85328 165486
rect 85008 165218 85050 165454
rect 85286 165218 85328 165454
rect 85008 165134 85328 165218
rect 85008 164898 85050 165134
rect 85286 164898 85328 165134
rect 85008 164866 85328 164898
rect 115728 165454 116048 165486
rect 115728 165218 115770 165454
rect 116006 165218 116048 165454
rect 115728 165134 116048 165218
rect 115728 164898 115770 165134
rect 116006 164898 116048 165134
rect 115728 164866 116048 164898
rect 146448 165454 146768 165486
rect 146448 165218 146490 165454
rect 146726 165218 146768 165454
rect 146448 165134 146768 165218
rect 146448 164898 146490 165134
rect 146726 164898 146768 165134
rect 146448 164866 146768 164898
rect 177168 165454 177488 165486
rect 177168 165218 177210 165454
rect 177446 165218 177488 165454
rect 177168 165134 177488 165218
rect 177168 164898 177210 165134
rect 177446 164898 177488 165134
rect 177168 164866 177488 164898
rect 207888 165454 208208 165486
rect 207888 165218 207930 165454
rect 208166 165218 208208 165454
rect 207888 165134 208208 165218
rect 207888 164898 207930 165134
rect 208166 164898 208208 165134
rect 207888 164866 208208 164898
rect 238608 165454 238928 165486
rect 238608 165218 238650 165454
rect 238886 165218 238928 165454
rect 238608 165134 238928 165218
rect 238608 164898 238650 165134
rect 238886 164898 238928 165134
rect 238608 164866 238928 164898
rect 269328 165454 269648 165486
rect 269328 165218 269370 165454
rect 269606 165218 269648 165454
rect 269328 165134 269648 165218
rect 269328 164898 269370 165134
rect 269606 164898 269648 165134
rect 269328 164866 269648 164898
rect 300048 165454 300368 165486
rect 300048 165218 300090 165454
rect 300326 165218 300368 165454
rect 300048 165134 300368 165218
rect 300048 164898 300090 165134
rect 300326 164898 300368 165134
rect 300048 164866 300368 164898
rect 330768 165454 331088 165486
rect 330768 165218 330810 165454
rect 331046 165218 331088 165454
rect 330768 165134 331088 165218
rect 330768 164898 330810 165134
rect 331046 164898 331088 165134
rect 330768 164866 331088 164898
rect 361488 165454 361808 165486
rect 361488 165218 361530 165454
rect 361766 165218 361808 165454
rect 361488 165134 361808 165218
rect 361488 164898 361530 165134
rect 361766 164898 361808 165134
rect 361488 164866 361808 164898
rect 392208 165454 392528 165486
rect 392208 165218 392250 165454
rect 392486 165218 392528 165454
rect 392208 165134 392528 165218
rect 392208 164898 392250 165134
rect 392486 164898 392528 165134
rect 392208 164866 392528 164898
rect 422928 165454 423248 165486
rect 422928 165218 422970 165454
rect 423206 165218 423248 165454
rect 422928 165134 423248 165218
rect 422928 164898 422970 165134
rect 423206 164898 423248 165134
rect 422928 164866 423248 164898
rect 453648 165454 453968 165486
rect 453648 165218 453690 165454
rect 453926 165218 453968 165454
rect 453648 165134 453968 165218
rect 453648 164898 453690 165134
rect 453926 164898 453968 165134
rect 453648 164866 453968 164898
rect 484368 165454 484688 165486
rect 484368 165218 484410 165454
rect 484646 165218 484688 165454
rect 484368 165134 484688 165218
rect 484368 164898 484410 165134
rect 484646 164898 484688 165134
rect 484368 164866 484688 164898
rect 515088 165454 515408 165486
rect 515088 165218 515130 165454
rect 515366 165218 515408 165454
rect 515088 165134 515408 165218
rect 515088 164898 515130 165134
rect 515366 164898 515408 165134
rect 515088 164866 515408 164898
rect 545808 165454 546128 165486
rect 545808 165218 545850 165454
rect 546086 165218 546128 165454
rect 545808 165134 546128 165218
rect 545808 164898 545850 165134
rect 546086 164898 546128 165134
rect 545808 164866 546128 164898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect 8208 147454 8528 147486
rect 8208 147218 8250 147454
rect 8486 147218 8528 147454
rect 8208 147134 8528 147218
rect 8208 146898 8250 147134
rect 8486 146898 8528 147134
rect 8208 146866 8528 146898
rect 38928 147454 39248 147486
rect 38928 147218 38970 147454
rect 39206 147218 39248 147454
rect 38928 147134 39248 147218
rect 38928 146898 38970 147134
rect 39206 146898 39248 147134
rect 38928 146866 39248 146898
rect 69648 147454 69968 147486
rect 69648 147218 69690 147454
rect 69926 147218 69968 147454
rect 69648 147134 69968 147218
rect 69648 146898 69690 147134
rect 69926 146898 69968 147134
rect 69648 146866 69968 146898
rect 100368 147454 100688 147486
rect 100368 147218 100410 147454
rect 100646 147218 100688 147454
rect 100368 147134 100688 147218
rect 100368 146898 100410 147134
rect 100646 146898 100688 147134
rect 100368 146866 100688 146898
rect 131088 147454 131408 147486
rect 131088 147218 131130 147454
rect 131366 147218 131408 147454
rect 131088 147134 131408 147218
rect 131088 146898 131130 147134
rect 131366 146898 131408 147134
rect 131088 146866 131408 146898
rect 161808 147454 162128 147486
rect 161808 147218 161850 147454
rect 162086 147218 162128 147454
rect 161808 147134 162128 147218
rect 161808 146898 161850 147134
rect 162086 146898 162128 147134
rect 161808 146866 162128 146898
rect 192528 147454 192848 147486
rect 192528 147218 192570 147454
rect 192806 147218 192848 147454
rect 192528 147134 192848 147218
rect 192528 146898 192570 147134
rect 192806 146898 192848 147134
rect 192528 146866 192848 146898
rect 223248 147454 223568 147486
rect 223248 147218 223290 147454
rect 223526 147218 223568 147454
rect 223248 147134 223568 147218
rect 223248 146898 223290 147134
rect 223526 146898 223568 147134
rect 223248 146866 223568 146898
rect 253968 147454 254288 147486
rect 253968 147218 254010 147454
rect 254246 147218 254288 147454
rect 253968 147134 254288 147218
rect 253968 146898 254010 147134
rect 254246 146898 254288 147134
rect 253968 146866 254288 146898
rect 284688 147454 285008 147486
rect 284688 147218 284730 147454
rect 284966 147218 285008 147454
rect 284688 147134 285008 147218
rect 284688 146898 284730 147134
rect 284966 146898 285008 147134
rect 284688 146866 285008 146898
rect 315408 147454 315728 147486
rect 315408 147218 315450 147454
rect 315686 147218 315728 147454
rect 315408 147134 315728 147218
rect 315408 146898 315450 147134
rect 315686 146898 315728 147134
rect 315408 146866 315728 146898
rect 346128 147454 346448 147486
rect 346128 147218 346170 147454
rect 346406 147218 346448 147454
rect 346128 147134 346448 147218
rect 346128 146898 346170 147134
rect 346406 146898 346448 147134
rect 346128 146866 346448 146898
rect 376848 147454 377168 147486
rect 376848 147218 376890 147454
rect 377126 147218 377168 147454
rect 376848 147134 377168 147218
rect 376848 146898 376890 147134
rect 377126 146898 377168 147134
rect 376848 146866 377168 146898
rect 407568 147454 407888 147486
rect 407568 147218 407610 147454
rect 407846 147218 407888 147454
rect 407568 147134 407888 147218
rect 407568 146898 407610 147134
rect 407846 146898 407888 147134
rect 407568 146866 407888 146898
rect 438288 147454 438608 147486
rect 438288 147218 438330 147454
rect 438566 147218 438608 147454
rect 438288 147134 438608 147218
rect 438288 146898 438330 147134
rect 438566 146898 438608 147134
rect 438288 146866 438608 146898
rect 469008 147454 469328 147486
rect 469008 147218 469050 147454
rect 469286 147218 469328 147454
rect 469008 147134 469328 147218
rect 469008 146898 469050 147134
rect 469286 146898 469328 147134
rect 469008 146866 469328 146898
rect 499728 147454 500048 147486
rect 499728 147218 499770 147454
rect 500006 147218 500048 147454
rect 499728 147134 500048 147218
rect 499728 146898 499770 147134
rect 500006 146898 500048 147134
rect 499728 146866 500048 146898
rect 530448 147454 530768 147486
rect 530448 147218 530490 147454
rect 530726 147218 530768 147454
rect 530448 147134 530768 147218
rect 530448 146898 530490 147134
rect 530726 146898 530768 147134
rect 530448 146866 530768 146898
rect 561168 147454 561488 147486
rect 561168 147218 561210 147454
rect 561446 147218 561488 147454
rect 561168 147134 561488 147218
rect 561168 146898 561210 147134
rect 561446 146898 561488 147134
rect 561168 146866 561488 146898
rect 567234 136894 567854 172338
rect 567234 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 567854 136894
rect 567234 136574 567854 136658
rect 567234 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 567854 136574
rect 23568 129454 23888 129486
rect 23568 129218 23610 129454
rect 23846 129218 23888 129454
rect 23568 129134 23888 129218
rect 23568 128898 23610 129134
rect 23846 128898 23888 129134
rect 23568 128866 23888 128898
rect 54288 129454 54608 129486
rect 54288 129218 54330 129454
rect 54566 129218 54608 129454
rect 54288 129134 54608 129218
rect 54288 128898 54330 129134
rect 54566 128898 54608 129134
rect 54288 128866 54608 128898
rect 85008 129454 85328 129486
rect 85008 129218 85050 129454
rect 85286 129218 85328 129454
rect 85008 129134 85328 129218
rect 85008 128898 85050 129134
rect 85286 128898 85328 129134
rect 85008 128866 85328 128898
rect 115728 129454 116048 129486
rect 115728 129218 115770 129454
rect 116006 129218 116048 129454
rect 115728 129134 116048 129218
rect 115728 128898 115770 129134
rect 116006 128898 116048 129134
rect 115728 128866 116048 128898
rect 146448 129454 146768 129486
rect 146448 129218 146490 129454
rect 146726 129218 146768 129454
rect 146448 129134 146768 129218
rect 146448 128898 146490 129134
rect 146726 128898 146768 129134
rect 146448 128866 146768 128898
rect 177168 129454 177488 129486
rect 177168 129218 177210 129454
rect 177446 129218 177488 129454
rect 177168 129134 177488 129218
rect 177168 128898 177210 129134
rect 177446 128898 177488 129134
rect 177168 128866 177488 128898
rect 207888 129454 208208 129486
rect 207888 129218 207930 129454
rect 208166 129218 208208 129454
rect 207888 129134 208208 129218
rect 207888 128898 207930 129134
rect 208166 128898 208208 129134
rect 207888 128866 208208 128898
rect 238608 129454 238928 129486
rect 238608 129218 238650 129454
rect 238886 129218 238928 129454
rect 238608 129134 238928 129218
rect 238608 128898 238650 129134
rect 238886 128898 238928 129134
rect 238608 128866 238928 128898
rect 269328 129454 269648 129486
rect 269328 129218 269370 129454
rect 269606 129218 269648 129454
rect 269328 129134 269648 129218
rect 269328 128898 269370 129134
rect 269606 128898 269648 129134
rect 269328 128866 269648 128898
rect 300048 129454 300368 129486
rect 300048 129218 300090 129454
rect 300326 129218 300368 129454
rect 300048 129134 300368 129218
rect 300048 128898 300090 129134
rect 300326 128898 300368 129134
rect 300048 128866 300368 128898
rect 330768 129454 331088 129486
rect 330768 129218 330810 129454
rect 331046 129218 331088 129454
rect 330768 129134 331088 129218
rect 330768 128898 330810 129134
rect 331046 128898 331088 129134
rect 330768 128866 331088 128898
rect 361488 129454 361808 129486
rect 361488 129218 361530 129454
rect 361766 129218 361808 129454
rect 361488 129134 361808 129218
rect 361488 128898 361530 129134
rect 361766 128898 361808 129134
rect 361488 128866 361808 128898
rect 392208 129454 392528 129486
rect 392208 129218 392250 129454
rect 392486 129218 392528 129454
rect 392208 129134 392528 129218
rect 392208 128898 392250 129134
rect 392486 128898 392528 129134
rect 392208 128866 392528 128898
rect 422928 129454 423248 129486
rect 422928 129218 422970 129454
rect 423206 129218 423248 129454
rect 422928 129134 423248 129218
rect 422928 128898 422970 129134
rect 423206 128898 423248 129134
rect 422928 128866 423248 128898
rect 453648 129454 453968 129486
rect 453648 129218 453690 129454
rect 453926 129218 453968 129454
rect 453648 129134 453968 129218
rect 453648 128898 453690 129134
rect 453926 128898 453968 129134
rect 453648 128866 453968 128898
rect 484368 129454 484688 129486
rect 484368 129218 484410 129454
rect 484646 129218 484688 129454
rect 484368 129134 484688 129218
rect 484368 128898 484410 129134
rect 484646 128898 484688 129134
rect 484368 128866 484688 128898
rect 515088 129454 515408 129486
rect 515088 129218 515130 129454
rect 515366 129218 515408 129454
rect 515088 129134 515408 129218
rect 515088 128898 515130 129134
rect 515366 128898 515408 129134
rect 515088 128866 515408 128898
rect 545808 129454 546128 129486
rect 545808 129218 545850 129454
rect 546086 129218 546128 129454
rect 545808 129134 546128 129218
rect 545808 128898 545850 129134
rect 546086 128898 546128 129134
rect 545808 128866 546128 128898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect 8208 111454 8528 111486
rect 8208 111218 8250 111454
rect 8486 111218 8528 111454
rect 8208 111134 8528 111218
rect 8208 110898 8250 111134
rect 8486 110898 8528 111134
rect 8208 110866 8528 110898
rect 38928 111454 39248 111486
rect 38928 111218 38970 111454
rect 39206 111218 39248 111454
rect 38928 111134 39248 111218
rect 38928 110898 38970 111134
rect 39206 110898 39248 111134
rect 38928 110866 39248 110898
rect 69648 111454 69968 111486
rect 69648 111218 69690 111454
rect 69926 111218 69968 111454
rect 69648 111134 69968 111218
rect 69648 110898 69690 111134
rect 69926 110898 69968 111134
rect 69648 110866 69968 110898
rect 100368 111454 100688 111486
rect 100368 111218 100410 111454
rect 100646 111218 100688 111454
rect 100368 111134 100688 111218
rect 100368 110898 100410 111134
rect 100646 110898 100688 111134
rect 100368 110866 100688 110898
rect 131088 111454 131408 111486
rect 131088 111218 131130 111454
rect 131366 111218 131408 111454
rect 131088 111134 131408 111218
rect 131088 110898 131130 111134
rect 131366 110898 131408 111134
rect 131088 110866 131408 110898
rect 161808 111454 162128 111486
rect 161808 111218 161850 111454
rect 162086 111218 162128 111454
rect 161808 111134 162128 111218
rect 161808 110898 161850 111134
rect 162086 110898 162128 111134
rect 161808 110866 162128 110898
rect 192528 111454 192848 111486
rect 192528 111218 192570 111454
rect 192806 111218 192848 111454
rect 192528 111134 192848 111218
rect 192528 110898 192570 111134
rect 192806 110898 192848 111134
rect 192528 110866 192848 110898
rect 223248 111454 223568 111486
rect 223248 111218 223290 111454
rect 223526 111218 223568 111454
rect 223248 111134 223568 111218
rect 223248 110898 223290 111134
rect 223526 110898 223568 111134
rect 223248 110866 223568 110898
rect 253968 111454 254288 111486
rect 253968 111218 254010 111454
rect 254246 111218 254288 111454
rect 253968 111134 254288 111218
rect 253968 110898 254010 111134
rect 254246 110898 254288 111134
rect 253968 110866 254288 110898
rect 284688 111454 285008 111486
rect 284688 111218 284730 111454
rect 284966 111218 285008 111454
rect 284688 111134 285008 111218
rect 284688 110898 284730 111134
rect 284966 110898 285008 111134
rect 284688 110866 285008 110898
rect 315408 111454 315728 111486
rect 315408 111218 315450 111454
rect 315686 111218 315728 111454
rect 315408 111134 315728 111218
rect 315408 110898 315450 111134
rect 315686 110898 315728 111134
rect 315408 110866 315728 110898
rect 346128 111454 346448 111486
rect 346128 111218 346170 111454
rect 346406 111218 346448 111454
rect 346128 111134 346448 111218
rect 346128 110898 346170 111134
rect 346406 110898 346448 111134
rect 346128 110866 346448 110898
rect 376848 111454 377168 111486
rect 376848 111218 376890 111454
rect 377126 111218 377168 111454
rect 376848 111134 377168 111218
rect 376848 110898 376890 111134
rect 377126 110898 377168 111134
rect 376848 110866 377168 110898
rect 407568 111454 407888 111486
rect 407568 111218 407610 111454
rect 407846 111218 407888 111454
rect 407568 111134 407888 111218
rect 407568 110898 407610 111134
rect 407846 110898 407888 111134
rect 407568 110866 407888 110898
rect 438288 111454 438608 111486
rect 438288 111218 438330 111454
rect 438566 111218 438608 111454
rect 438288 111134 438608 111218
rect 438288 110898 438330 111134
rect 438566 110898 438608 111134
rect 438288 110866 438608 110898
rect 469008 111454 469328 111486
rect 469008 111218 469050 111454
rect 469286 111218 469328 111454
rect 469008 111134 469328 111218
rect 469008 110898 469050 111134
rect 469286 110898 469328 111134
rect 469008 110866 469328 110898
rect 499728 111454 500048 111486
rect 499728 111218 499770 111454
rect 500006 111218 500048 111454
rect 499728 111134 500048 111218
rect 499728 110898 499770 111134
rect 500006 110898 500048 111134
rect 499728 110866 500048 110898
rect 530448 111454 530768 111486
rect 530448 111218 530490 111454
rect 530726 111218 530768 111454
rect 530448 111134 530768 111218
rect 530448 110898 530490 111134
rect 530726 110898 530768 111134
rect 530448 110866 530768 110898
rect 561168 111454 561488 111486
rect 561168 111218 561210 111454
rect 561446 111218 561488 111454
rect 561168 111134 561488 111218
rect 561168 110898 561210 111134
rect 561446 110898 561488 111134
rect 561168 110866 561488 110898
rect 567234 100894 567854 136338
rect 567234 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 567854 100894
rect 567234 100574 567854 100658
rect 567234 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 567854 100574
rect 23568 93454 23888 93486
rect 23568 93218 23610 93454
rect 23846 93218 23888 93454
rect 23568 93134 23888 93218
rect 23568 92898 23610 93134
rect 23846 92898 23888 93134
rect 23568 92866 23888 92898
rect 54288 93454 54608 93486
rect 54288 93218 54330 93454
rect 54566 93218 54608 93454
rect 54288 93134 54608 93218
rect 54288 92898 54330 93134
rect 54566 92898 54608 93134
rect 54288 92866 54608 92898
rect 85008 93454 85328 93486
rect 85008 93218 85050 93454
rect 85286 93218 85328 93454
rect 85008 93134 85328 93218
rect 85008 92898 85050 93134
rect 85286 92898 85328 93134
rect 85008 92866 85328 92898
rect 115728 93454 116048 93486
rect 115728 93218 115770 93454
rect 116006 93218 116048 93454
rect 115728 93134 116048 93218
rect 115728 92898 115770 93134
rect 116006 92898 116048 93134
rect 115728 92866 116048 92898
rect 146448 93454 146768 93486
rect 146448 93218 146490 93454
rect 146726 93218 146768 93454
rect 146448 93134 146768 93218
rect 146448 92898 146490 93134
rect 146726 92898 146768 93134
rect 146448 92866 146768 92898
rect 177168 93454 177488 93486
rect 177168 93218 177210 93454
rect 177446 93218 177488 93454
rect 177168 93134 177488 93218
rect 177168 92898 177210 93134
rect 177446 92898 177488 93134
rect 177168 92866 177488 92898
rect 207888 93454 208208 93486
rect 207888 93218 207930 93454
rect 208166 93218 208208 93454
rect 207888 93134 208208 93218
rect 207888 92898 207930 93134
rect 208166 92898 208208 93134
rect 207888 92866 208208 92898
rect 238608 93454 238928 93486
rect 238608 93218 238650 93454
rect 238886 93218 238928 93454
rect 238608 93134 238928 93218
rect 238608 92898 238650 93134
rect 238886 92898 238928 93134
rect 238608 92866 238928 92898
rect 269328 93454 269648 93486
rect 269328 93218 269370 93454
rect 269606 93218 269648 93454
rect 269328 93134 269648 93218
rect 269328 92898 269370 93134
rect 269606 92898 269648 93134
rect 269328 92866 269648 92898
rect 300048 93454 300368 93486
rect 300048 93218 300090 93454
rect 300326 93218 300368 93454
rect 300048 93134 300368 93218
rect 300048 92898 300090 93134
rect 300326 92898 300368 93134
rect 300048 92866 300368 92898
rect 330768 93454 331088 93486
rect 330768 93218 330810 93454
rect 331046 93218 331088 93454
rect 330768 93134 331088 93218
rect 330768 92898 330810 93134
rect 331046 92898 331088 93134
rect 330768 92866 331088 92898
rect 361488 93454 361808 93486
rect 361488 93218 361530 93454
rect 361766 93218 361808 93454
rect 361488 93134 361808 93218
rect 361488 92898 361530 93134
rect 361766 92898 361808 93134
rect 361488 92866 361808 92898
rect 392208 93454 392528 93486
rect 392208 93218 392250 93454
rect 392486 93218 392528 93454
rect 392208 93134 392528 93218
rect 392208 92898 392250 93134
rect 392486 92898 392528 93134
rect 392208 92866 392528 92898
rect 422928 93454 423248 93486
rect 422928 93218 422970 93454
rect 423206 93218 423248 93454
rect 422928 93134 423248 93218
rect 422928 92898 422970 93134
rect 423206 92898 423248 93134
rect 422928 92866 423248 92898
rect 453648 93454 453968 93486
rect 453648 93218 453690 93454
rect 453926 93218 453968 93454
rect 453648 93134 453968 93218
rect 453648 92898 453690 93134
rect 453926 92898 453968 93134
rect 453648 92866 453968 92898
rect 484368 93454 484688 93486
rect 484368 93218 484410 93454
rect 484646 93218 484688 93454
rect 484368 93134 484688 93218
rect 484368 92898 484410 93134
rect 484646 92898 484688 93134
rect 484368 92866 484688 92898
rect 515088 93454 515408 93486
rect 515088 93218 515130 93454
rect 515366 93218 515408 93454
rect 515088 93134 515408 93218
rect 515088 92898 515130 93134
rect 515366 92898 515408 93134
rect 515088 92866 515408 92898
rect 545808 93454 546128 93486
rect 545808 93218 545850 93454
rect 546086 93218 546128 93454
rect 545808 93134 546128 93218
rect 545808 92898 545850 93134
rect 546086 92898 546128 93134
rect 545808 92866 546128 92898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect 8208 75454 8528 75486
rect 8208 75218 8250 75454
rect 8486 75218 8528 75454
rect 8208 75134 8528 75218
rect 8208 74898 8250 75134
rect 8486 74898 8528 75134
rect 8208 74866 8528 74898
rect 38928 75454 39248 75486
rect 38928 75218 38970 75454
rect 39206 75218 39248 75454
rect 38928 75134 39248 75218
rect 38928 74898 38970 75134
rect 39206 74898 39248 75134
rect 38928 74866 39248 74898
rect 69648 75454 69968 75486
rect 69648 75218 69690 75454
rect 69926 75218 69968 75454
rect 69648 75134 69968 75218
rect 69648 74898 69690 75134
rect 69926 74898 69968 75134
rect 69648 74866 69968 74898
rect 100368 75454 100688 75486
rect 100368 75218 100410 75454
rect 100646 75218 100688 75454
rect 100368 75134 100688 75218
rect 100368 74898 100410 75134
rect 100646 74898 100688 75134
rect 100368 74866 100688 74898
rect 131088 75454 131408 75486
rect 131088 75218 131130 75454
rect 131366 75218 131408 75454
rect 131088 75134 131408 75218
rect 131088 74898 131130 75134
rect 131366 74898 131408 75134
rect 131088 74866 131408 74898
rect 161808 75454 162128 75486
rect 161808 75218 161850 75454
rect 162086 75218 162128 75454
rect 161808 75134 162128 75218
rect 161808 74898 161850 75134
rect 162086 74898 162128 75134
rect 161808 74866 162128 74898
rect 192528 75454 192848 75486
rect 192528 75218 192570 75454
rect 192806 75218 192848 75454
rect 192528 75134 192848 75218
rect 192528 74898 192570 75134
rect 192806 74898 192848 75134
rect 192528 74866 192848 74898
rect 223248 75454 223568 75486
rect 223248 75218 223290 75454
rect 223526 75218 223568 75454
rect 223248 75134 223568 75218
rect 223248 74898 223290 75134
rect 223526 74898 223568 75134
rect 223248 74866 223568 74898
rect 253968 75454 254288 75486
rect 253968 75218 254010 75454
rect 254246 75218 254288 75454
rect 253968 75134 254288 75218
rect 253968 74898 254010 75134
rect 254246 74898 254288 75134
rect 253968 74866 254288 74898
rect 284688 75454 285008 75486
rect 284688 75218 284730 75454
rect 284966 75218 285008 75454
rect 284688 75134 285008 75218
rect 284688 74898 284730 75134
rect 284966 74898 285008 75134
rect 284688 74866 285008 74898
rect 315408 75454 315728 75486
rect 315408 75218 315450 75454
rect 315686 75218 315728 75454
rect 315408 75134 315728 75218
rect 315408 74898 315450 75134
rect 315686 74898 315728 75134
rect 315408 74866 315728 74898
rect 346128 75454 346448 75486
rect 346128 75218 346170 75454
rect 346406 75218 346448 75454
rect 346128 75134 346448 75218
rect 346128 74898 346170 75134
rect 346406 74898 346448 75134
rect 346128 74866 346448 74898
rect 376848 75454 377168 75486
rect 376848 75218 376890 75454
rect 377126 75218 377168 75454
rect 376848 75134 377168 75218
rect 376848 74898 376890 75134
rect 377126 74898 377168 75134
rect 376848 74866 377168 74898
rect 407568 75454 407888 75486
rect 407568 75218 407610 75454
rect 407846 75218 407888 75454
rect 407568 75134 407888 75218
rect 407568 74898 407610 75134
rect 407846 74898 407888 75134
rect 407568 74866 407888 74898
rect 438288 75454 438608 75486
rect 438288 75218 438330 75454
rect 438566 75218 438608 75454
rect 438288 75134 438608 75218
rect 438288 74898 438330 75134
rect 438566 74898 438608 75134
rect 438288 74866 438608 74898
rect 469008 75454 469328 75486
rect 469008 75218 469050 75454
rect 469286 75218 469328 75454
rect 469008 75134 469328 75218
rect 469008 74898 469050 75134
rect 469286 74898 469328 75134
rect 469008 74866 469328 74898
rect 499728 75454 500048 75486
rect 499728 75218 499770 75454
rect 500006 75218 500048 75454
rect 499728 75134 500048 75218
rect 499728 74898 499770 75134
rect 500006 74898 500048 75134
rect 499728 74866 500048 74898
rect 530448 75454 530768 75486
rect 530448 75218 530490 75454
rect 530726 75218 530768 75454
rect 530448 75134 530768 75218
rect 530448 74898 530490 75134
rect 530726 74898 530768 75134
rect 530448 74866 530768 74898
rect 561168 75454 561488 75486
rect 561168 75218 561210 75454
rect 561446 75218 561488 75454
rect 561168 75134 561488 75218
rect 561168 74898 561210 75134
rect 561446 74898 561488 75134
rect 561168 74866 561488 74898
rect 567234 64894 567854 100338
rect 567234 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 567854 64894
rect 567234 64574 567854 64658
rect 567234 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 567854 64574
rect 23568 57454 23888 57486
rect 23568 57218 23610 57454
rect 23846 57218 23888 57454
rect 23568 57134 23888 57218
rect 23568 56898 23610 57134
rect 23846 56898 23888 57134
rect 23568 56866 23888 56898
rect 54288 57454 54608 57486
rect 54288 57218 54330 57454
rect 54566 57218 54608 57454
rect 54288 57134 54608 57218
rect 54288 56898 54330 57134
rect 54566 56898 54608 57134
rect 54288 56866 54608 56898
rect 85008 57454 85328 57486
rect 85008 57218 85050 57454
rect 85286 57218 85328 57454
rect 85008 57134 85328 57218
rect 85008 56898 85050 57134
rect 85286 56898 85328 57134
rect 85008 56866 85328 56898
rect 115728 57454 116048 57486
rect 115728 57218 115770 57454
rect 116006 57218 116048 57454
rect 115728 57134 116048 57218
rect 115728 56898 115770 57134
rect 116006 56898 116048 57134
rect 115728 56866 116048 56898
rect 146448 57454 146768 57486
rect 146448 57218 146490 57454
rect 146726 57218 146768 57454
rect 146448 57134 146768 57218
rect 146448 56898 146490 57134
rect 146726 56898 146768 57134
rect 146448 56866 146768 56898
rect 177168 57454 177488 57486
rect 177168 57218 177210 57454
rect 177446 57218 177488 57454
rect 177168 57134 177488 57218
rect 177168 56898 177210 57134
rect 177446 56898 177488 57134
rect 177168 56866 177488 56898
rect 207888 57454 208208 57486
rect 207888 57218 207930 57454
rect 208166 57218 208208 57454
rect 207888 57134 208208 57218
rect 207888 56898 207930 57134
rect 208166 56898 208208 57134
rect 207888 56866 208208 56898
rect 238608 57454 238928 57486
rect 238608 57218 238650 57454
rect 238886 57218 238928 57454
rect 238608 57134 238928 57218
rect 238608 56898 238650 57134
rect 238886 56898 238928 57134
rect 238608 56866 238928 56898
rect 269328 57454 269648 57486
rect 269328 57218 269370 57454
rect 269606 57218 269648 57454
rect 269328 57134 269648 57218
rect 269328 56898 269370 57134
rect 269606 56898 269648 57134
rect 269328 56866 269648 56898
rect 300048 57454 300368 57486
rect 300048 57218 300090 57454
rect 300326 57218 300368 57454
rect 300048 57134 300368 57218
rect 300048 56898 300090 57134
rect 300326 56898 300368 57134
rect 300048 56866 300368 56898
rect 330768 57454 331088 57486
rect 330768 57218 330810 57454
rect 331046 57218 331088 57454
rect 330768 57134 331088 57218
rect 330768 56898 330810 57134
rect 331046 56898 331088 57134
rect 330768 56866 331088 56898
rect 361488 57454 361808 57486
rect 361488 57218 361530 57454
rect 361766 57218 361808 57454
rect 361488 57134 361808 57218
rect 361488 56898 361530 57134
rect 361766 56898 361808 57134
rect 361488 56866 361808 56898
rect 392208 57454 392528 57486
rect 392208 57218 392250 57454
rect 392486 57218 392528 57454
rect 392208 57134 392528 57218
rect 392208 56898 392250 57134
rect 392486 56898 392528 57134
rect 392208 56866 392528 56898
rect 422928 57454 423248 57486
rect 422928 57218 422970 57454
rect 423206 57218 423248 57454
rect 422928 57134 423248 57218
rect 422928 56898 422970 57134
rect 423206 56898 423248 57134
rect 422928 56866 423248 56898
rect 453648 57454 453968 57486
rect 453648 57218 453690 57454
rect 453926 57218 453968 57454
rect 453648 57134 453968 57218
rect 453648 56898 453690 57134
rect 453926 56898 453968 57134
rect 453648 56866 453968 56898
rect 484368 57454 484688 57486
rect 484368 57218 484410 57454
rect 484646 57218 484688 57454
rect 484368 57134 484688 57218
rect 484368 56898 484410 57134
rect 484646 56898 484688 57134
rect 484368 56866 484688 56898
rect 515088 57454 515408 57486
rect 515088 57218 515130 57454
rect 515366 57218 515408 57454
rect 515088 57134 515408 57218
rect 515088 56898 515130 57134
rect 515366 56898 515408 57134
rect 515088 56866 515408 56898
rect 545808 57454 546128 57486
rect 545808 57218 545850 57454
rect 546086 57218 546128 57454
rect 545808 57134 546128 57218
rect 545808 56898 545850 57134
rect 546086 56898 546128 57134
rect 545808 56866 546128 56898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect 8208 39454 8528 39486
rect 8208 39218 8250 39454
rect 8486 39218 8528 39454
rect 8208 39134 8528 39218
rect 8208 38898 8250 39134
rect 8486 38898 8528 39134
rect 8208 38866 8528 38898
rect 38928 39454 39248 39486
rect 38928 39218 38970 39454
rect 39206 39218 39248 39454
rect 38928 39134 39248 39218
rect 38928 38898 38970 39134
rect 39206 38898 39248 39134
rect 38928 38866 39248 38898
rect 69648 39454 69968 39486
rect 69648 39218 69690 39454
rect 69926 39218 69968 39454
rect 69648 39134 69968 39218
rect 69648 38898 69690 39134
rect 69926 38898 69968 39134
rect 69648 38866 69968 38898
rect 100368 39454 100688 39486
rect 100368 39218 100410 39454
rect 100646 39218 100688 39454
rect 100368 39134 100688 39218
rect 100368 38898 100410 39134
rect 100646 38898 100688 39134
rect 100368 38866 100688 38898
rect 131088 39454 131408 39486
rect 131088 39218 131130 39454
rect 131366 39218 131408 39454
rect 131088 39134 131408 39218
rect 131088 38898 131130 39134
rect 131366 38898 131408 39134
rect 131088 38866 131408 38898
rect 161808 39454 162128 39486
rect 161808 39218 161850 39454
rect 162086 39218 162128 39454
rect 161808 39134 162128 39218
rect 161808 38898 161850 39134
rect 162086 38898 162128 39134
rect 161808 38866 162128 38898
rect 192528 39454 192848 39486
rect 192528 39218 192570 39454
rect 192806 39218 192848 39454
rect 192528 39134 192848 39218
rect 192528 38898 192570 39134
rect 192806 38898 192848 39134
rect 192528 38866 192848 38898
rect 223248 39454 223568 39486
rect 223248 39218 223290 39454
rect 223526 39218 223568 39454
rect 223248 39134 223568 39218
rect 223248 38898 223290 39134
rect 223526 38898 223568 39134
rect 223248 38866 223568 38898
rect 253968 39454 254288 39486
rect 253968 39218 254010 39454
rect 254246 39218 254288 39454
rect 253968 39134 254288 39218
rect 253968 38898 254010 39134
rect 254246 38898 254288 39134
rect 253968 38866 254288 38898
rect 284688 39454 285008 39486
rect 284688 39218 284730 39454
rect 284966 39218 285008 39454
rect 284688 39134 285008 39218
rect 284688 38898 284730 39134
rect 284966 38898 285008 39134
rect 284688 38866 285008 38898
rect 315408 39454 315728 39486
rect 315408 39218 315450 39454
rect 315686 39218 315728 39454
rect 315408 39134 315728 39218
rect 315408 38898 315450 39134
rect 315686 38898 315728 39134
rect 315408 38866 315728 38898
rect 346128 39454 346448 39486
rect 346128 39218 346170 39454
rect 346406 39218 346448 39454
rect 346128 39134 346448 39218
rect 346128 38898 346170 39134
rect 346406 38898 346448 39134
rect 346128 38866 346448 38898
rect 376848 39454 377168 39486
rect 376848 39218 376890 39454
rect 377126 39218 377168 39454
rect 376848 39134 377168 39218
rect 376848 38898 376890 39134
rect 377126 38898 377168 39134
rect 376848 38866 377168 38898
rect 407568 39454 407888 39486
rect 407568 39218 407610 39454
rect 407846 39218 407888 39454
rect 407568 39134 407888 39218
rect 407568 38898 407610 39134
rect 407846 38898 407888 39134
rect 407568 38866 407888 38898
rect 438288 39454 438608 39486
rect 438288 39218 438330 39454
rect 438566 39218 438608 39454
rect 438288 39134 438608 39218
rect 438288 38898 438330 39134
rect 438566 38898 438608 39134
rect 438288 38866 438608 38898
rect 469008 39454 469328 39486
rect 469008 39218 469050 39454
rect 469286 39218 469328 39454
rect 469008 39134 469328 39218
rect 469008 38898 469050 39134
rect 469286 38898 469328 39134
rect 469008 38866 469328 38898
rect 499728 39454 500048 39486
rect 499728 39218 499770 39454
rect 500006 39218 500048 39454
rect 499728 39134 500048 39218
rect 499728 38898 499770 39134
rect 500006 38898 500048 39134
rect 499728 38866 500048 38898
rect 530448 39454 530768 39486
rect 530448 39218 530490 39454
rect 530726 39218 530768 39454
rect 530448 39134 530768 39218
rect 530448 38898 530490 39134
rect 530726 38898 530768 39134
rect 530448 38866 530768 38898
rect 561168 39454 561488 39486
rect 561168 39218 561210 39454
rect 561446 39218 561488 39454
rect 561168 39134 561488 39218
rect 561168 38898 561210 39134
rect 561446 38898 561488 39134
rect 561168 38866 561488 38898
rect 567234 28894 567854 64338
rect 567234 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 567854 28894
rect 567234 28574 567854 28658
rect 567234 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 567854 28574
rect 23568 21454 23888 21486
rect 23568 21218 23610 21454
rect 23846 21218 23888 21454
rect 23568 21134 23888 21218
rect 23568 20898 23610 21134
rect 23846 20898 23888 21134
rect 23568 20866 23888 20898
rect 54288 21454 54608 21486
rect 54288 21218 54330 21454
rect 54566 21218 54608 21454
rect 54288 21134 54608 21218
rect 54288 20898 54330 21134
rect 54566 20898 54608 21134
rect 54288 20866 54608 20898
rect 85008 21454 85328 21486
rect 85008 21218 85050 21454
rect 85286 21218 85328 21454
rect 85008 21134 85328 21218
rect 85008 20898 85050 21134
rect 85286 20898 85328 21134
rect 85008 20866 85328 20898
rect 115728 21454 116048 21486
rect 115728 21218 115770 21454
rect 116006 21218 116048 21454
rect 115728 21134 116048 21218
rect 115728 20898 115770 21134
rect 116006 20898 116048 21134
rect 115728 20866 116048 20898
rect 146448 21454 146768 21486
rect 146448 21218 146490 21454
rect 146726 21218 146768 21454
rect 146448 21134 146768 21218
rect 146448 20898 146490 21134
rect 146726 20898 146768 21134
rect 146448 20866 146768 20898
rect 177168 21454 177488 21486
rect 177168 21218 177210 21454
rect 177446 21218 177488 21454
rect 177168 21134 177488 21218
rect 177168 20898 177210 21134
rect 177446 20898 177488 21134
rect 177168 20866 177488 20898
rect 207888 21454 208208 21486
rect 207888 21218 207930 21454
rect 208166 21218 208208 21454
rect 207888 21134 208208 21218
rect 207888 20898 207930 21134
rect 208166 20898 208208 21134
rect 207888 20866 208208 20898
rect 238608 21454 238928 21486
rect 238608 21218 238650 21454
rect 238886 21218 238928 21454
rect 238608 21134 238928 21218
rect 238608 20898 238650 21134
rect 238886 20898 238928 21134
rect 238608 20866 238928 20898
rect 269328 21454 269648 21486
rect 269328 21218 269370 21454
rect 269606 21218 269648 21454
rect 269328 21134 269648 21218
rect 269328 20898 269370 21134
rect 269606 20898 269648 21134
rect 269328 20866 269648 20898
rect 300048 21454 300368 21486
rect 300048 21218 300090 21454
rect 300326 21218 300368 21454
rect 300048 21134 300368 21218
rect 300048 20898 300090 21134
rect 300326 20898 300368 21134
rect 300048 20866 300368 20898
rect 330768 21454 331088 21486
rect 330768 21218 330810 21454
rect 331046 21218 331088 21454
rect 330768 21134 331088 21218
rect 330768 20898 330810 21134
rect 331046 20898 331088 21134
rect 330768 20866 331088 20898
rect 361488 21454 361808 21486
rect 361488 21218 361530 21454
rect 361766 21218 361808 21454
rect 361488 21134 361808 21218
rect 361488 20898 361530 21134
rect 361766 20898 361808 21134
rect 361488 20866 361808 20898
rect 392208 21454 392528 21486
rect 392208 21218 392250 21454
rect 392486 21218 392528 21454
rect 392208 21134 392528 21218
rect 392208 20898 392250 21134
rect 392486 20898 392528 21134
rect 392208 20866 392528 20898
rect 422928 21454 423248 21486
rect 422928 21218 422970 21454
rect 423206 21218 423248 21454
rect 422928 21134 423248 21218
rect 422928 20898 422970 21134
rect 423206 20898 423248 21134
rect 422928 20866 423248 20898
rect 453648 21454 453968 21486
rect 453648 21218 453690 21454
rect 453926 21218 453968 21454
rect 453648 21134 453968 21218
rect 453648 20898 453690 21134
rect 453926 20898 453968 21134
rect 453648 20866 453968 20898
rect 484368 21454 484688 21486
rect 484368 21218 484410 21454
rect 484646 21218 484688 21454
rect 484368 21134 484688 21218
rect 484368 20898 484410 21134
rect 484646 20898 484688 21134
rect 484368 20866 484688 20898
rect 515088 21454 515408 21486
rect 515088 21218 515130 21454
rect 515366 21218 515408 21454
rect 515088 21134 515408 21218
rect 515088 20898 515130 21134
rect 515366 20898 515408 21134
rect 515088 20866 515408 20898
rect 545808 21454 546128 21486
rect 545808 21218 545850 21454
rect 546086 21218 546128 21454
rect 545808 21134 546128 21218
rect 545808 20898 545850 21134
rect 546086 20898 546128 21134
rect 545808 20866 546128 20898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect 8208 3454 8528 3486
rect 8208 3218 8250 3454
rect 8486 3218 8528 3454
rect 8208 3134 8528 3218
rect 8208 2898 8250 3134
rect 8486 2898 8528 3134
rect 8208 2866 8528 2898
rect 38928 3454 39248 3486
rect 38928 3218 38970 3454
rect 39206 3218 39248 3454
rect 38928 3134 39248 3218
rect 38928 2898 38970 3134
rect 39206 2898 39248 3134
rect 38928 2866 39248 2898
rect 69648 3454 69968 3486
rect 69648 3218 69690 3454
rect 69926 3218 69968 3454
rect 69648 3134 69968 3218
rect 69648 2898 69690 3134
rect 69926 2898 69968 3134
rect 69648 2866 69968 2898
rect 100368 3454 100688 3486
rect 100368 3218 100410 3454
rect 100646 3218 100688 3454
rect 100368 3134 100688 3218
rect 100368 2898 100410 3134
rect 100646 2898 100688 3134
rect 100368 2866 100688 2898
rect 131088 3454 131408 3486
rect 131088 3218 131130 3454
rect 131366 3218 131408 3454
rect 131088 3134 131408 3218
rect 131088 2898 131130 3134
rect 131366 2898 131408 3134
rect 131088 2866 131408 2898
rect 161808 3454 162128 3486
rect 161808 3218 161850 3454
rect 162086 3218 162128 3454
rect 161808 3134 162128 3218
rect 161808 2898 161850 3134
rect 162086 2898 162128 3134
rect 161808 2866 162128 2898
rect 192528 3454 192848 3486
rect 192528 3218 192570 3454
rect 192806 3218 192848 3454
rect 192528 3134 192848 3218
rect 192528 2898 192570 3134
rect 192806 2898 192848 3134
rect 192528 2866 192848 2898
rect 223248 3454 223568 3486
rect 223248 3218 223290 3454
rect 223526 3218 223568 3454
rect 223248 3134 223568 3218
rect 223248 2898 223290 3134
rect 223526 2898 223568 3134
rect 223248 2866 223568 2898
rect 253968 3454 254288 3486
rect 253968 3218 254010 3454
rect 254246 3218 254288 3454
rect 253968 3134 254288 3218
rect 253968 2898 254010 3134
rect 254246 2898 254288 3134
rect 253968 2866 254288 2898
rect 284688 3454 285008 3486
rect 284688 3218 284730 3454
rect 284966 3218 285008 3454
rect 284688 3134 285008 3218
rect 284688 2898 284730 3134
rect 284966 2898 285008 3134
rect 284688 2866 285008 2898
rect 315408 3454 315728 3486
rect 315408 3218 315450 3454
rect 315686 3218 315728 3454
rect 315408 3134 315728 3218
rect 315408 2898 315450 3134
rect 315686 2898 315728 3134
rect 315408 2866 315728 2898
rect 346128 3454 346448 3486
rect 346128 3218 346170 3454
rect 346406 3218 346448 3454
rect 346128 3134 346448 3218
rect 346128 2898 346170 3134
rect 346406 2898 346448 3134
rect 346128 2866 346448 2898
rect 376848 3454 377168 3486
rect 376848 3218 376890 3454
rect 377126 3218 377168 3454
rect 376848 3134 377168 3218
rect 376848 2898 376890 3134
rect 377126 2898 377168 3134
rect 376848 2866 377168 2898
rect 407568 3454 407888 3486
rect 407568 3218 407610 3454
rect 407846 3218 407888 3454
rect 407568 3134 407888 3218
rect 407568 2898 407610 3134
rect 407846 2898 407888 3134
rect 407568 2866 407888 2898
rect 438288 3454 438608 3486
rect 438288 3218 438330 3454
rect 438566 3218 438608 3454
rect 438288 3134 438608 3218
rect 438288 2898 438330 3134
rect 438566 2898 438608 3134
rect 438288 2866 438608 2898
rect 469008 3454 469328 3486
rect 469008 3218 469050 3454
rect 469286 3218 469328 3454
rect 469008 3134 469328 3218
rect 469008 2898 469050 3134
rect 469286 2898 469328 3134
rect 469008 2866 469328 2898
rect 499728 3454 500048 3486
rect 499728 3218 499770 3454
rect 500006 3218 500048 3454
rect 499728 3134 500048 3218
rect 499728 2898 499770 3134
rect 500006 2898 500048 3134
rect 499728 2866 500048 2898
rect 530448 3454 530768 3486
rect 530448 3218 530490 3454
rect 530726 3218 530768 3454
rect 530448 3134 530768 3218
rect 530448 2898 530490 3134
rect 530726 2898 530768 3134
rect 530448 2866 530768 2898
rect 561168 3454 561488 3486
rect 561168 3218 561210 3454
rect 561446 3218 561488 3454
rect 561168 3134 561488 3218
rect 561168 2898 561210 3134
rect 561446 2898 561488 3134
rect 561168 2866 561488 2898
rect 531267 1460 531333 1461
rect 531267 1396 531268 1460
rect 531332 1396 531333 1460
rect 531267 1395 531333 1396
rect 531270 645 531330 1395
rect 559419 916 559485 917
rect 559419 852 559420 916
rect 559484 852 559485 916
rect 559419 851 559485 852
rect 531267 644 531333 645
rect 531267 580 531268 644
rect 531332 580 531333 644
rect 531267 579 531333 580
rect 559422 509 559482 851
rect 559419 508 559485 509
rect 559419 444 559420 508
rect 559484 444 559485 508
rect 559419 443 559485 444
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 -2000
rect 5514 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 6134 -2266
rect 5514 -2586 6134 -2502
rect 5514 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 6134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 -2000
rect 9234 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 9854 -4186
rect 9234 -4506 9854 -4422
rect 9234 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 9854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 -2000
rect 23514 -3226 24134 -2000
rect 23514 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 24134 -3226
rect 23514 -3546 24134 -3462
rect 23514 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 24134 -3546
rect 23514 -3814 24134 -3782
rect 27234 -5146 27854 -2000
rect 27234 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 27854 -5146
rect 27234 -5466 27854 -5382
rect 27234 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 27854 -5466
rect 27234 -5734 27854 -5702
rect 12954 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 13574 -6106
rect 12954 -6426 13574 -6342
rect 12954 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 13574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 -2000
rect 41514 -2266 42134 -2000
rect 41514 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 42134 -2266
rect 41514 -2586 42134 -2502
rect 41514 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 42134 -2586
rect 41514 -3814 42134 -2822
rect 45234 -4186 45854 -2000
rect 45234 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 45854 -4186
rect 45234 -4506 45854 -4422
rect 45234 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 45854 -4506
rect 45234 -5734 45854 -4742
rect 30954 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 31574 -7066
rect 30954 -7386 31574 -7302
rect 30954 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 31574 -7386
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 -2000
rect 59514 -3226 60134 -2000
rect 59514 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 60134 -3226
rect 59514 -3546 60134 -3462
rect 59514 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 60134 -3546
rect 59514 -3814 60134 -3782
rect 63234 -5146 63854 -2000
rect 63234 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 63854 -5146
rect 63234 -5466 63854 -5382
rect 63234 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 63854 -5466
rect 63234 -5734 63854 -5702
rect 48954 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 49574 -6106
rect 48954 -6426 49574 -6342
rect 48954 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 49574 -6426
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 -2000
rect 77514 -2266 78134 -2000
rect 77514 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 78134 -2266
rect 77514 -2586 78134 -2502
rect 77514 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 78134 -2586
rect 77514 -3814 78134 -2822
rect 81234 -4186 81854 -2000
rect 81234 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 81854 -4186
rect 81234 -4506 81854 -4422
rect 81234 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 81854 -4506
rect 81234 -5734 81854 -4742
rect 66954 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 67574 -7066
rect 66954 -7386 67574 -7302
rect 66954 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 67574 -7386
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 -2000
rect 95514 -3226 96134 -2000
rect 95514 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 96134 -3226
rect 95514 -3546 96134 -3462
rect 95514 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 96134 -3546
rect 95514 -3814 96134 -3782
rect 99234 -5146 99854 -2000
rect 99234 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 99854 -5146
rect 99234 -5466 99854 -5382
rect 99234 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 99854 -5466
rect 99234 -5734 99854 -5702
rect 84954 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 85574 -6106
rect 84954 -6426 85574 -6342
rect 84954 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 85574 -6426
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 -2000
rect 113514 -2266 114134 -2000
rect 113514 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 114134 -2266
rect 113514 -2586 114134 -2502
rect 113514 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 114134 -2586
rect 113514 -3814 114134 -2822
rect 117234 -4186 117854 -2000
rect 117234 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 117854 -4186
rect 117234 -4506 117854 -4422
rect 117234 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 117854 -4506
rect 117234 -5734 117854 -4742
rect 102954 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 103574 -7066
rect 102954 -7386 103574 -7302
rect 102954 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 103574 -7386
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 -2000
rect 131514 -3226 132134 -2000
rect 131514 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 132134 -3226
rect 131514 -3546 132134 -3462
rect 131514 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 132134 -3546
rect 131514 -3814 132134 -3782
rect 135234 -5146 135854 -2000
rect 135234 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 135854 -5146
rect 135234 -5466 135854 -5382
rect 135234 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 135854 -5466
rect 135234 -5734 135854 -5702
rect 120954 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 121574 -6106
rect 120954 -6426 121574 -6342
rect 120954 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 121574 -6426
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 -2000
rect 149514 -2266 150134 -2000
rect 149514 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 150134 -2266
rect 149514 -2586 150134 -2502
rect 149514 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 150134 -2586
rect 149514 -3814 150134 -2822
rect 153234 -4186 153854 -2000
rect 153234 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 153854 -4186
rect 153234 -4506 153854 -4422
rect 153234 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 153854 -4506
rect 153234 -5734 153854 -4742
rect 138954 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 139574 -7066
rect 138954 -7386 139574 -7302
rect 138954 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 139574 -7386
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 -2000
rect 167514 -3226 168134 -2000
rect 167514 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 168134 -3226
rect 167514 -3546 168134 -3462
rect 167514 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 168134 -3546
rect 167514 -3814 168134 -3782
rect 171234 -5146 171854 -2000
rect 171234 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 171854 -5146
rect 171234 -5466 171854 -5382
rect 171234 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 171854 -5466
rect 171234 -5734 171854 -5702
rect 156954 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 157574 -6106
rect 156954 -6426 157574 -6342
rect 156954 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 157574 -6426
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 -2000
rect 185514 -2266 186134 -2000
rect 185514 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 186134 -2266
rect 185514 -2586 186134 -2502
rect 185514 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 186134 -2586
rect 185514 -3814 186134 -2822
rect 189234 -4186 189854 -2000
rect 189234 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 189854 -4186
rect 189234 -4506 189854 -4422
rect 189234 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 189854 -4506
rect 189234 -5734 189854 -4742
rect 174954 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 175574 -7066
rect 174954 -7386 175574 -7302
rect 174954 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 175574 -7386
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 -2000
rect 203514 -3226 204134 -2000
rect 203514 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 204134 -3226
rect 203514 -3546 204134 -3462
rect 203514 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 204134 -3546
rect 203514 -3814 204134 -3782
rect 207234 -5146 207854 -2000
rect 207234 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 207854 -5146
rect 207234 -5466 207854 -5382
rect 207234 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 207854 -5466
rect 207234 -5734 207854 -5702
rect 192954 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 193574 -6106
rect 192954 -6426 193574 -6342
rect 192954 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 193574 -6426
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 -2000
rect 221514 -2266 222134 -2000
rect 221514 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 222134 -2266
rect 221514 -2586 222134 -2502
rect 221514 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 222134 -2586
rect 221514 -3814 222134 -2822
rect 225234 -4186 225854 -2000
rect 225234 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 225854 -4186
rect 225234 -4506 225854 -4422
rect 225234 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 225854 -4506
rect 225234 -5734 225854 -4742
rect 210954 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 211574 -7066
rect 210954 -7386 211574 -7302
rect 210954 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 211574 -7386
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 -2000
rect 239514 -3226 240134 -2000
rect 239514 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 240134 -3226
rect 239514 -3546 240134 -3462
rect 239514 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 240134 -3546
rect 239514 -3814 240134 -3782
rect 243234 -5146 243854 -2000
rect 243234 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 243854 -5146
rect 243234 -5466 243854 -5382
rect 243234 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 243854 -5466
rect 243234 -5734 243854 -5702
rect 228954 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 229574 -6106
rect 228954 -6426 229574 -6342
rect 228954 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 229574 -6426
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 -2000
rect 257514 -2266 258134 -2000
rect 257514 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 258134 -2266
rect 257514 -2586 258134 -2502
rect 257514 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 258134 -2586
rect 257514 -3814 258134 -2822
rect 261234 -4186 261854 -2000
rect 261234 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 261854 -4186
rect 261234 -4506 261854 -4422
rect 261234 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 261854 -4506
rect 261234 -5734 261854 -4742
rect 246954 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 247574 -7066
rect 246954 -7386 247574 -7302
rect 246954 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 247574 -7386
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 -2000
rect 275514 -3226 276134 -2000
rect 275514 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 276134 -3226
rect 275514 -3546 276134 -3462
rect 275514 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 276134 -3546
rect 275514 -3814 276134 -3782
rect 279234 -5146 279854 -2000
rect 279234 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 279854 -5146
rect 279234 -5466 279854 -5382
rect 279234 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 279854 -5466
rect 279234 -5734 279854 -5702
rect 264954 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 265574 -6106
rect 264954 -6426 265574 -6342
rect 264954 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 265574 -6426
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 -2000
rect 293514 -2266 294134 -2000
rect 293514 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 294134 -2266
rect 293514 -2586 294134 -2502
rect 293514 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 294134 -2586
rect 293514 -3814 294134 -2822
rect 297234 -4186 297854 -2000
rect 297234 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 297854 -4186
rect 297234 -4506 297854 -4422
rect 297234 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 297854 -4506
rect 297234 -5734 297854 -4742
rect 282954 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 283574 -7066
rect 282954 -7386 283574 -7302
rect 282954 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 283574 -7386
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 -2000
rect 311514 -3226 312134 -2000
rect 311514 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 312134 -3226
rect 311514 -3546 312134 -3462
rect 311514 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 312134 -3546
rect 311514 -3814 312134 -3782
rect 315234 -5146 315854 -2000
rect 315234 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 315854 -5146
rect 315234 -5466 315854 -5382
rect 315234 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 315854 -5466
rect 315234 -5734 315854 -5702
rect 300954 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 301574 -6106
rect 300954 -6426 301574 -6342
rect 300954 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 301574 -6426
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 -2000
rect 329514 -2266 330134 -2000
rect 329514 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 330134 -2266
rect 329514 -2586 330134 -2502
rect 329514 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 330134 -2586
rect 329514 -3814 330134 -2822
rect 333234 -4186 333854 -2000
rect 333234 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 333854 -4186
rect 333234 -4506 333854 -4422
rect 333234 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 333854 -4506
rect 333234 -5734 333854 -4742
rect 318954 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 319574 -7066
rect 318954 -7386 319574 -7302
rect 318954 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 319574 -7386
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 -2000
rect 347514 -3226 348134 -2000
rect 347514 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 348134 -3226
rect 347514 -3546 348134 -3462
rect 347514 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 348134 -3546
rect 347514 -3814 348134 -3782
rect 351234 -5146 351854 -2000
rect 351234 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 351854 -5146
rect 351234 -5466 351854 -5382
rect 351234 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 351854 -5466
rect 351234 -5734 351854 -5702
rect 336954 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 337574 -6106
rect 336954 -6426 337574 -6342
rect 336954 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 337574 -6426
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 -2000
rect 365514 -2266 366134 -2000
rect 365514 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 366134 -2266
rect 365514 -2586 366134 -2502
rect 365514 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 366134 -2586
rect 365514 -3814 366134 -2822
rect 369234 -4186 369854 -2000
rect 369234 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 369854 -4186
rect 369234 -4506 369854 -4422
rect 369234 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 369854 -4506
rect 369234 -5734 369854 -4742
rect 354954 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 355574 -7066
rect 354954 -7386 355574 -7302
rect 354954 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 355574 -7386
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 -2000
rect 383514 -3226 384134 -2000
rect 383514 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 384134 -3226
rect 383514 -3546 384134 -3462
rect 383514 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 384134 -3546
rect 383514 -3814 384134 -3782
rect 387234 -5146 387854 -2000
rect 387234 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 387854 -5146
rect 387234 -5466 387854 -5382
rect 387234 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 387854 -5466
rect 387234 -5734 387854 -5702
rect 372954 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 373574 -6106
rect 372954 -6426 373574 -6342
rect 372954 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 373574 -6426
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 -2000
rect 401514 -2266 402134 -2000
rect 401514 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 402134 -2266
rect 401514 -2586 402134 -2502
rect 401514 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 402134 -2586
rect 401514 -3814 402134 -2822
rect 405234 -4186 405854 -2000
rect 405234 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 405854 -4186
rect 405234 -4506 405854 -4422
rect 405234 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 405854 -4506
rect 405234 -5734 405854 -4742
rect 390954 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 391574 -7066
rect 390954 -7386 391574 -7302
rect 390954 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 391574 -7386
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 -2000
rect 419514 -3226 420134 -2000
rect 419514 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 420134 -3226
rect 419514 -3546 420134 -3462
rect 419514 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 420134 -3546
rect 419514 -3814 420134 -3782
rect 423234 -5146 423854 -2000
rect 423234 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 423854 -5146
rect 423234 -5466 423854 -5382
rect 423234 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 423854 -5466
rect 423234 -5734 423854 -5702
rect 408954 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 409574 -6106
rect 408954 -6426 409574 -6342
rect 408954 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 409574 -6426
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 -2000
rect 437514 -2266 438134 -2000
rect 437514 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 438134 -2266
rect 437514 -2586 438134 -2502
rect 437514 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 438134 -2586
rect 437514 -3814 438134 -2822
rect 441234 -4186 441854 -2000
rect 441234 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 441854 -4186
rect 441234 -4506 441854 -4422
rect 441234 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 441854 -4506
rect 441234 -5734 441854 -4742
rect 426954 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 427574 -7066
rect 426954 -7386 427574 -7302
rect 426954 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 427574 -7386
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 -2000
rect 455514 -3226 456134 -2000
rect 455514 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 456134 -3226
rect 455514 -3546 456134 -3462
rect 455514 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 456134 -3546
rect 455514 -3814 456134 -3782
rect 459234 -5146 459854 -2000
rect 459234 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 459854 -5146
rect 459234 -5466 459854 -5382
rect 459234 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 459854 -5466
rect 459234 -5734 459854 -5702
rect 444954 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 445574 -6106
rect 444954 -6426 445574 -6342
rect 444954 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 445574 -6426
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 -2000
rect 473514 -2266 474134 -2000
rect 473514 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 474134 -2266
rect 473514 -2586 474134 -2502
rect 473514 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 474134 -2586
rect 473514 -3814 474134 -2822
rect 477234 -4186 477854 -2000
rect 477234 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 477854 -4186
rect 477234 -4506 477854 -4422
rect 477234 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 477854 -4506
rect 477234 -5734 477854 -4742
rect 462954 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 463574 -7066
rect 462954 -7386 463574 -7302
rect 462954 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 463574 -7386
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 -2000
rect 491514 -3226 492134 -2000
rect 491514 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 492134 -3226
rect 491514 -3546 492134 -3462
rect 491514 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 492134 -3546
rect 491514 -3814 492134 -3782
rect 495234 -5146 495854 -2000
rect 495234 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 495854 -5146
rect 495234 -5466 495854 -5382
rect 495234 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 495854 -5466
rect 495234 -5734 495854 -5702
rect 480954 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 481574 -6106
rect 480954 -6426 481574 -6342
rect 480954 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 481574 -6426
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 -2000
rect 509514 -2266 510134 -2000
rect 509514 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 510134 -2266
rect 509514 -2586 510134 -2502
rect 509514 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 510134 -2586
rect 509514 -3814 510134 -2822
rect 513234 -4186 513854 -2000
rect 513234 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 513854 -4186
rect 513234 -4506 513854 -4422
rect 513234 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 513854 -4506
rect 513234 -5734 513854 -4742
rect 498954 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 499574 -7066
rect 498954 -7386 499574 -7302
rect 498954 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 499574 -7386
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 -2000
rect 527514 -3226 528134 -2000
rect 527514 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 528134 -3226
rect 527514 -3546 528134 -3462
rect 527514 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 528134 -3546
rect 527514 -3814 528134 -3782
rect 531234 -5146 531854 -2000
rect 531234 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 531854 -5146
rect 531234 -5466 531854 -5382
rect 531234 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 531854 -5466
rect 531234 -5734 531854 -5702
rect 516954 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 517574 -6106
rect 516954 -6426 517574 -6342
rect 516954 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 517574 -6426
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 -2000
rect 545514 -2266 546134 -2000
rect 545514 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 546134 -2266
rect 545514 -2586 546134 -2502
rect 545514 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 546134 -2586
rect 545514 -3814 546134 -2822
rect 549234 -4186 549854 -2000
rect 549234 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 549854 -4186
rect 549234 -4506 549854 -4422
rect 549234 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 549854 -4506
rect 549234 -5734 549854 -4742
rect 534954 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 535574 -7066
rect 534954 -7386 535574 -7302
rect 534954 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 535574 -7386
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 -2000
rect 563514 -3226 564134 -2000
rect 563514 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 564134 -3226
rect 563514 -3546 564134 -3462
rect 563514 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 564134 -3546
rect 563514 -3814 564134 -3782
rect 567234 -5146 567854 28338
rect 567234 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 567854 -5146
rect 567234 -5466 567854 -5382
rect 567234 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 567854 -5466
rect 567234 -5734 567854 -5702
rect 570954 680614 571574 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 581514 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 582134 706758
rect 581514 706438 582134 706522
rect 581514 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 582134 706438
rect 570954 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 571574 680614
rect 570954 680294 571574 680378
rect 570954 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 571574 680294
rect 570954 644614 571574 680058
rect 570954 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 571574 644614
rect 570954 644294 571574 644378
rect 570954 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 571574 644294
rect 570954 608614 571574 644058
rect 570954 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 571574 608614
rect 570954 608294 571574 608378
rect 570954 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 571574 608294
rect 570954 572614 571574 608058
rect 570954 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 571574 572614
rect 570954 572294 571574 572378
rect 570954 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 571574 572294
rect 570954 536614 571574 572058
rect 570954 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 571574 536614
rect 570954 536294 571574 536378
rect 570954 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 571574 536294
rect 570954 500614 571574 536058
rect 570954 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 571574 500614
rect 570954 500294 571574 500378
rect 570954 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 571574 500294
rect 570954 464614 571574 500058
rect 570954 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 571574 464614
rect 570954 464294 571574 464378
rect 570954 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 571574 464294
rect 570954 428614 571574 464058
rect 570954 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 571574 428614
rect 570954 428294 571574 428378
rect 570954 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 571574 428294
rect 570954 392614 571574 428058
rect 570954 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 571574 392614
rect 570954 392294 571574 392378
rect 570954 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 571574 392294
rect 570954 356614 571574 392058
rect 570954 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 571574 356614
rect 570954 356294 571574 356378
rect 570954 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 571574 356294
rect 570954 320614 571574 356058
rect 570954 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 571574 320614
rect 570954 320294 571574 320378
rect 570954 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 571574 320294
rect 570954 284614 571574 320058
rect 570954 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 571574 284614
rect 570954 284294 571574 284378
rect 570954 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 571574 284294
rect 570954 248614 571574 284058
rect 570954 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 571574 248614
rect 570954 248294 571574 248378
rect 570954 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 571574 248294
rect 570954 212614 571574 248058
rect 570954 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 571574 212614
rect 570954 212294 571574 212378
rect 570954 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 571574 212294
rect 570954 176614 571574 212058
rect 570954 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 571574 176614
rect 570954 176294 571574 176378
rect 570954 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 571574 176294
rect 570954 140614 571574 176058
rect 570954 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 571574 140614
rect 570954 140294 571574 140378
rect 570954 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 571574 140294
rect 570954 104614 571574 140058
rect 570954 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 571574 104614
rect 570954 104294 571574 104378
rect 570954 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 571574 104294
rect 570954 68614 571574 104058
rect 570954 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 571574 68614
rect 570954 68294 571574 68378
rect 570954 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 571574 68294
rect 570954 32614 571574 68058
rect 570954 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 571574 32614
rect 570954 32294 571574 32378
rect 570954 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 571574 32294
rect 552954 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 553574 -6106
rect 552954 -6426 553574 -6342
rect 552954 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 553574 -6426
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 32058
rect 577794 704838 578414 705830
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 581514 691174 582134 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -2266 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 587850 691174
rect 587230 690854 587850 690938
rect 587230 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 587850 690854
rect 587230 655174 587850 690618
rect 587230 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 587850 655174
rect 587230 654854 587850 654938
rect 587230 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 587850 654854
rect 587230 619174 587850 654618
rect 587230 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 587850 619174
rect 587230 618854 587850 618938
rect 587230 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 587850 618854
rect 587230 583174 587850 618618
rect 587230 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 587850 583174
rect 587230 582854 587850 582938
rect 587230 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 587850 582854
rect 587230 547174 587850 582618
rect 587230 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 587850 547174
rect 587230 546854 587850 546938
rect 587230 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 587850 546854
rect 587230 511174 587850 546618
rect 587230 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 587850 511174
rect 587230 510854 587850 510938
rect 587230 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 587850 510854
rect 587230 475174 587850 510618
rect 587230 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 587850 475174
rect 587230 474854 587850 474938
rect 587230 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 587850 474854
rect 587230 439174 587850 474618
rect 587230 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 587850 439174
rect 587230 438854 587850 438938
rect 587230 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 587850 438854
rect 587230 403174 587850 438618
rect 587230 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 587850 403174
rect 587230 402854 587850 402938
rect 587230 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 587850 402854
rect 587230 367174 587850 402618
rect 587230 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 587850 367174
rect 587230 366854 587850 366938
rect 587230 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 587850 366854
rect 587230 331174 587850 366618
rect 587230 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 587850 331174
rect 587230 330854 587850 330938
rect 587230 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 587850 330854
rect 587230 295174 587850 330618
rect 587230 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 587850 295174
rect 587230 294854 587850 294938
rect 587230 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 587850 294854
rect 587230 259174 587850 294618
rect 587230 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 587850 259174
rect 587230 258854 587850 258938
rect 587230 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 587850 258854
rect 587230 223174 587850 258618
rect 587230 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 587850 223174
rect 587230 222854 587850 222938
rect 587230 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 587850 222854
rect 587230 187174 587850 222618
rect 587230 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 587850 187174
rect 587230 186854 587850 186938
rect 587230 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 587850 186854
rect 587230 151174 587850 186618
rect 587230 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 587850 151174
rect 587230 150854 587850 150938
rect 587230 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 587850 150854
rect 587230 115174 587850 150618
rect 587230 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 587850 115174
rect 587230 114854 587850 114938
rect 587230 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 587850 114854
rect 587230 79174 587850 114618
rect 587230 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 587850 79174
rect 587230 78854 587850 78938
rect 587230 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 587850 78854
rect 587230 43174 587850 78618
rect 587230 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 587850 43174
rect 587230 42854 587850 42938
rect 587230 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 587850 42854
rect 587230 7174 587850 42618
rect 587230 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 587850 7174
rect 587230 6854 587850 6938
rect 587230 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 587850 6854
rect 581514 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 582134 -2266
rect 581514 -2586 582134 -2502
rect 581514 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 582134 -2586
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect 588190 672854 588810 672938
rect 588190 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect 588190 637174 588810 672618
rect 588190 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect 588190 636854 588810 636938
rect 588190 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect 588190 601174 588810 636618
rect 588190 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect 588190 600854 588810 600938
rect 588190 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect 588190 565174 588810 600618
rect 588190 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect 588190 564854 588810 564938
rect 588190 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect 588190 529174 588810 564618
rect 588190 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect 588190 528854 588810 528938
rect 588190 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect 588190 493174 588810 528618
rect 588190 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect 588190 492854 588810 492938
rect 588190 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect 588190 457174 588810 492618
rect 588190 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect 588190 456854 588810 456938
rect 588190 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect 588190 421174 588810 456618
rect 588190 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 588190 420854 588810 420938
rect 588190 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 588190 385174 588810 420618
rect 588190 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 588190 384854 588810 384938
rect 588190 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 588190 349174 588810 384618
rect 588190 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 588190 348854 588810 348938
rect 588190 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 588190 313174 588810 348618
rect 588190 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 588190 312854 588810 312938
rect 588190 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 588190 277174 588810 312618
rect 588190 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 588190 276854 588810 276938
rect 588190 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 588190 241174 588810 276618
rect 588190 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 588190 240854 588810 240938
rect 588190 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 588190 205174 588810 240618
rect 588190 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 588190 204854 588810 204938
rect 588190 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 588190 169174 588810 204618
rect 588190 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 588190 168854 588810 168938
rect 588190 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 588190 133174 588810 168618
rect 588190 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 588190 132854 588810 132938
rect 588190 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 588190 97174 588810 132618
rect 588190 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 588190 96854 588810 96938
rect 588190 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 588190 61174 588810 96618
rect 588190 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 588190 60854 588810 60938
rect 588190 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 588190 25174 588810 60618
rect 588190 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect 588190 24854 588810 24938
rect 588190 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect 588190 -3226 588810 24618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 589770 694894
rect 589150 694574 589770 694658
rect 589150 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 589770 694574
rect 589150 658894 589770 694338
rect 589150 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 589770 658894
rect 589150 658574 589770 658658
rect 589150 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 589770 658574
rect 589150 622894 589770 658338
rect 589150 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 589770 622894
rect 589150 622574 589770 622658
rect 589150 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 589770 622574
rect 589150 586894 589770 622338
rect 589150 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 589770 586894
rect 589150 586574 589770 586658
rect 589150 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 589770 586574
rect 589150 550894 589770 586338
rect 589150 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 589770 550894
rect 589150 550574 589770 550658
rect 589150 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 589770 550574
rect 589150 514894 589770 550338
rect 589150 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 589770 514894
rect 589150 514574 589770 514658
rect 589150 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 589770 514574
rect 589150 478894 589770 514338
rect 589150 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 589770 478894
rect 589150 478574 589770 478658
rect 589150 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 589770 478574
rect 589150 442894 589770 478338
rect 589150 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 589770 442894
rect 589150 442574 589770 442658
rect 589150 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 589770 442574
rect 589150 406894 589770 442338
rect 589150 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 589770 406894
rect 589150 406574 589770 406658
rect 589150 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 589770 406574
rect 589150 370894 589770 406338
rect 589150 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 589770 370894
rect 589150 370574 589770 370658
rect 589150 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 589770 370574
rect 589150 334894 589770 370338
rect 589150 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 589770 334894
rect 589150 334574 589770 334658
rect 589150 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 589770 334574
rect 589150 298894 589770 334338
rect 589150 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 589770 298894
rect 589150 298574 589770 298658
rect 589150 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 589770 298574
rect 589150 262894 589770 298338
rect 589150 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 589770 262894
rect 589150 262574 589770 262658
rect 589150 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 589770 262574
rect 589150 226894 589770 262338
rect 589150 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 589770 226894
rect 589150 226574 589770 226658
rect 589150 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 589770 226574
rect 589150 190894 589770 226338
rect 589150 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 589770 190894
rect 589150 190574 589770 190658
rect 589150 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 589770 190574
rect 589150 154894 589770 190338
rect 589150 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 589770 154894
rect 589150 154574 589770 154658
rect 589150 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 589770 154574
rect 589150 118894 589770 154338
rect 589150 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 589770 118894
rect 589150 118574 589770 118658
rect 589150 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 589770 118574
rect 589150 82894 589770 118338
rect 589150 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 589770 82894
rect 589150 82574 589770 82658
rect 589150 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 589770 82574
rect 589150 46894 589770 82338
rect 589150 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 589770 46894
rect 589150 46574 589770 46658
rect 589150 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 589770 46574
rect 589150 10894 589770 46338
rect 589150 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 589770 10894
rect 589150 10574 589770 10658
rect 589150 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 589770 10574
rect 589150 -4186 589770 10338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect 590110 676574 590730 676658
rect 590110 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect 590110 640894 590730 676338
rect 590110 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect 590110 640574 590730 640658
rect 590110 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect 590110 604894 590730 640338
rect 590110 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect 590110 604574 590730 604658
rect 590110 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect 590110 568894 590730 604338
rect 590110 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect 590110 568574 590730 568658
rect 590110 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect 590110 532894 590730 568338
rect 590110 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect 590110 532574 590730 532658
rect 590110 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect 590110 496894 590730 532338
rect 590110 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect 590110 496574 590730 496658
rect 590110 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect 590110 460894 590730 496338
rect 590110 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect 590110 460574 590730 460658
rect 590110 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect 590110 424894 590730 460338
rect 590110 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 590110 424574 590730 424658
rect 590110 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 590110 388894 590730 424338
rect 590110 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 590110 388574 590730 388658
rect 590110 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 590110 352894 590730 388338
rect 590110 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 590110 352574 590730 352658
rect 590110 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 590110 316894 590730 352338
rect 590110 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 590110 316574 590730 316658
rect 590110 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 590110 280894 590730 316338
rect 590110 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 590110 280574 590730 280658
rect 590110 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 590110 244894 590730 280338
rect 590110 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 590110 244574 590730 244658
rect 590110 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 590110 208894 590730 244338
rect 590110 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 590110 208574 590730 208658
rect 590110 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 590110 172894 590730 208338
rect 590110 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 590110 172574 590730 172658
rect 590110 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 590110 136894 590730 172338
rect 590110 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 590110 136574 590730 136658
rect 590110 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 590110 100894 590730 136338
rect 590110 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 590110 100574 590730 100658
rect 590110 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 590110 64894 590730 100338
rect 590110 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 590110 64574 590730 64658
rect 590110 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 590110 28894 590730 64338
rect 590110 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect 590110 28574 590730 28658
rect 590110 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect 590110 -5146 590730 28338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 591690 698614
rect 591070 698294 591690 698378
rect 591070 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 591690 698294
rect 591070 662614 591690 698058
rect 591070 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 591690 662614
rect 591070 662294 591690 662378
rect 591070 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 591690 662294
rect 591070 626614 591690 662058
rect 591070 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 591690 626614
rect 591070 626294 591690 626378
rect 591070 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 591690 626294
rect 591070 590614 591690 626058
rect 591070 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 591690 590614
rect 591070 590294 591690 590378
rect 591070 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 591690 590294
rect 591070 554614 591690 590058
rect 591070 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 591690 554614
rect 591070 554294 591690 554378
rect 591070 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 591690 554294
rect 591070 518614 591690 554058
rect 591070 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 591690 518614
rect 591070 518294 591690 518378
rect 591070 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 591690 518294
rect 591070 482614 591690 518058
rect 591070 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 591690 482614
rect 591070 482294 591690 482378
rect 591070 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 591690 482294
rect 591070 446614 591690 482058
rect 591070 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 591690 446614
rect 591070 446294 591690 446378
rect 591070 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 591690 446294
rect 591070 410614 591690 446058
rect 591070 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 591690 410614
rect 591070 410294 591690 410378
rect 591070 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 591690 410294
rect 591070 374614 591690 410058
rect 591070 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 591690 374614
rect 591070 374294 591690 374378
rect 591070 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 591690 374294
rect 591070 338614 591690 374058
rect 591070 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 591690 338614
rect 591070 338294 591690 338378
rect 591070 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 591690 338294
rect 591070 302614 591690 338058
rect 591070 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 591690 302614
rect 591070 302294 591690 302378
rect 591070 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 591690 302294
rect 591070 266614 591690 302058
rect 591070 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 591690 266614
rect 591070 266294 591690 266378
rect 591070 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 591690 266294
rect 591070 230614 591690 266058
rect 591070 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 591690 230614
rect 591070 230294 591690 230378
rect 591070 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 591690 230294
rect 591070 194614 591690 230058
rect 591070 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 591690 194614
rect 591070 194294 591690 194378
rect 591070 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 591690 194294
rect 591070 158614 591690 194058
rect 591070 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 591690 158614
rect 591070 158294 591690 158378
rect 591070 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 591690 158294
rect 591070 122614 591690 158058
rect 591070 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 591690 122614
rect 591070 122294 591690 122378
rect 591070 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 591690 122294
rect 591070 86614 591690 122058
rect 591070 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 591690 86614
rect 591070 86294 591690 86378
rect 591070 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 591690 86294
rect 591070 50614 591690 86058
rect 591070 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 591690 50614
rect 591070 50294 591690 50378
rect 591070 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 591690 50294
rect 591070 14614 591690 50058
rect 591070 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 591690 14614
rect 591070 14294 591690 14378
rect 591070 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 591690 14294
rect 591070 -6106 591690 14058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect 592030 680294 592650 680378
rect 592030 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect 592030 644614 592650 680058
rect 592030 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect 592030 644294 592650 644378
rect 592030 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect 592030 608614 592650 644058
rect 592030 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect 592030 608294 592650 608378
rect 592030 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect 592030 572614 592650 608058
rect 592030 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect 592030 572294 592650 572378
rect 592030 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect 592030 536614 592650 572058
rect 592030 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect 592030 536294 592650 536378
rect 592030 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect 592030 500614 592650 536058
rect 592030 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect 592030 500294 592650 500378
rect 592030 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect 592030 464614 592650 500058
rect 592030 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect 592030 464294 592650 464378
rect 592030 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect 592030 428614 592650 464058
rect 592030 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 592030 428294 592650 428378
rect 592030 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 592030 392614 592650 428058
rect 592030 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 592030 392294 592650 392378
rect 592030 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 592030 356614 592650 392058
rect 592030 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 592030 356294 592650 356378
rect 592030 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 592030 320614 592650 356058
rect 592030 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 592030 320294 592650 320378
rect 592030 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 592030 284614 592650 320058
rect 592030 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 592030 284294 592650 284378
rect 592030 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 592030 248614 592650 284058
rect 592030 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 592030 248294 592650 248378
rect 592030 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 592030 212614 592650 248058
rect 592030 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 592030 212294 592650 212378
rect 592030 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 592030 176614 592650 212058
rect 592030 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 592030 176294 592650 176378
rect 592030 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 592030 140614 592650 176058
rect 592030 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 592030 140294 592650 140378
rect 592030 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 592030 104614 592650 140058
rect 592030 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 592030 104294 592650 104378
rect 592030 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 592030 68614 592650 104058
rect 592030 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 592030 68294 592650 68378
rect 592030 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 592030 32614 592650 68058
rect 592030 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect 592030 32294 592650 32378
rect 592030 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect 570954 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 571574 -7066
rect 570954 -7386 571574 -7302
rect 570954 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 571574 -7386
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 680378 -8458 680614
rect -8374 680378 -8138 680614
rect -8694 680058 -8458 680294
rect -8374 680058 -8138 680294
rect -8694 644378 -8458 644614
rect -8374 644378 -8138 644614
rect -8694 644058 -8458 644294
rect -8374 644058 -8138 644294
rect -8694 608378 -8458 608614
rect -8374 608378 -8138 608614
rect -8694 608058 -8458 608294
rect -8374 608058 -8138 608294
rect -8694 572378 -8458 572614
rect -8374 572378 -8138 572614
rect -8694 572058 -8458 572294
rect -8374 572058 -8138 572294
rect -8694 536378 -8458 536614
rect -8374 536378 -8138 536614
rect -8694 536058 -8458 536294
rect -8374 536058 -8138 536294
rect -8694 500378 -8458 500614
rect -8374 500378 -8138 500614
rect -8694 500058 -8458 500294
rect -8374 500058 -8138 500294
rect -8694 464378 -8458 464614
rect -8374 464378 -8138 464614
rect -8694 464058 -8458 464294
rect -8374 464058 -8138 464294
rect -8694 428378 -8458 428614
rect -8374 428378 -8138 428614
rect -8694 428058 -8458 428294
rect -8374 428058 -8138 428294
rect -8694 392378 -8458 392614
rect -8374 392378 -8138 392614
rect -8694 392058 -8458 392294
rect -8374 392058 -8138 392294
rect -8694 356378 -8458 356614
rect -8374 356378 -8138 356614
rect -8694 356058 -8458 356294
rect -8374 356058 -8138 356294
rect -8694 320378 -8458 320614
rect -8374 320378 -8138 320614
rect -8694 320058 -8458 320294
rect -8374 320058 -8138 320294
rect -8694 284378 -8458 284614
rect -8374 284378 -8138 284614
rect -8694 284058 -8458 284294
rect -8374 284058 -8138 284294
rect -8694 248378 -8458 248614
rect -8374 248378 -8138 248614
rect -8694 248058 -8458 248294
rect -8374 248058 -8138 248294
rect -8694 212378 -8458 212614
rect -8374 212378 -8138 212614
rect -8694 212058 -8458 212294
rect -8374 212058 -8138 212294
rect -8694 176378 -8458 176614
rect -8374 176378 -8138 176614
rect -8694 176058 -8458 176294
rect -8374 176058 -8138 176294
rect -8694 140378 -8458 140614
rect -8374 140378 -8138 140614
rect -8694 140058 -8458 140294
rect -8374 140058 -8138 140294
rect -8694 104378 -8458 104614
rect -8374 104378 -8138 104614
rect -8694 104058 -8458 104294
rect -8374 104058 -8138 104294
rect -8694 68378 -8458 68614
rect -8374 68378 -8138 68614
rect -8694 68058 -8458 68294
rect -8374 68058 -8138 68294
rect -8694 32378 -8458 32614
rect -8374 32378 -8138 32614
rect -8694 32058 -8458 32294
rect -8374 32058 -8138 32294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12986 710362 13222 710598
rect 13306 710362 13542 710598
rect 12986 710042 13222 710278
rect 13306 710042 13542 710278
rect -7734 698378 -7498 698614
rect -7414 698378 -7178 698614
rect -7734 698058 -7498 698294
rect -7414 698058 -7178 698294
rect -7734 662378 -7498 662614
rect -7414 662378 -7178 662614
rect -7734 662058 -7498 662294
rect -7414 662058 -7178 662294
rect -7734 626378 -7498 626614
rect -7414 626378 -7178 626614
rect -7734 626058 -7498 626294
rect -7414 626058 -7178 626294
rect -7734 590378 -7498 590614
rect -7414 590378 -7178 590614
rect -7734 590058 -7498 590294
rect -7414 590058 -7178 590294
rect -7734 554378 -7498 554614
rect -7414 554378 -7178 554614
rect -7734 554058 -7498 554294
rect -7414 554058 -7178 554294
rect -7734 518378 -7498 518614
rect -7414 518378 -7178 518614
rect -7734 518058 -7498 518294
rect -7414 518058 -7178 518294
rect -7734 482378 -7498 482614
rect -7414 482378 -7178 482614
rect -7734 482058 -7498 482294
rect -7414 482058 -7178 482294
rect -7734 446378 -7498 446614
rect -7414 446378 -7178 446614
rect -7734 446058 -7498 446294
rect -7414 446058 -7178 446294
rect -7734 410378 -7498 410614
rect -7414 410378 -7178 410614
rect -7734 410058 -7498 410294
rect -7414 410058 -7178 410294
rect -7734 374378 -7498 374614
rect -7414 374378 -7178 374614
rect -7734 374058 -7498 374294
rect -7414 374058 -7178 374294
rect -7734 338378 -7498 338614
rect -7414 338378 -7178 338614
rect -7734 338058 -7498 338294
rect -7414 338058 -7178 338294
rect -7734 302378 -7498 302614
rect -7414 302378 -7178 302614
rect -7734 302058 -7498 302294
rect -7414 302058 -7178 302294
rect -7734 266378 -7498 266614
rect -7414 266378 -7178 266614
rect -7734 266058 -7498 266294
rect -7414 266058 -7178 266294
rect -7734 230378 -7498 230614
rect -7414 230378 -7178 230614
rect -7734 230058 -7498 230294
rect -7414 230058 -7178 230294
rect -7734 194378 -7498 194614
rect -7414 194378 -7178 194614
rect -7734 194058 -7498 194294
rect -7414 194058 -7178 194294
rect -7734 158378 -7498 158614
rect -7414 158378 -7178 158614
rect -7734 158058 -7498 158294
rect -7414 158058 -7178 158294
rect -7734 122378 -7498 122614
rect -7414 122378 -7178 122614
rect -7734 122058 -7498 122294
rect -7414 122058 -7178 122294
rect -7734 86378 -7498 86614
rect -7414 86378 -7178 86614
rect -7734 86058 -7498 86294
rect -7414 86058 -7178 86294
rect -7734 50378 -7498 50614
rect -7414 50378 -7178 50614
rect -7734 50058 -7498 50294
rect -7414 50058 -7178 50294
rect -7734 14378 -7498 14614
rect -7414 14378 -7178 14614
rect -7734 14058 -7498 14294
rect -7414 14058 -7178 14294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 676658 -6538 676894
rect -6454 676658 -6218 676894
rect -6774 676338 -6538 676574
rect -6454 676338 -6218 676574
rect -6774 640658 -6538 640894
rect -6454 640658 -6218 640894
rect -6774 640338 -6538 640574
rect -6454 640338 -6218 640574
rect -6774 604658 -6538 604894
rect -6454 604658 -6218 604894
rect -6774 604338 -6538 604574
rect -6454 604338 -6218 604574
rect -6774 568658 -6538 568894
rect -6454 568658 -6218 568894
rect -6774 568338 -6538 568574
rect -6454 568338 -6218 568574
rect -6774 532658 -6538 532894
rect -6454 532658 -6218 532894
rect -6774 532338 -6538 532574
rect -6454 532338 -6218 532574
rect -6774 496658 -6538 496894
rect -6454 496658 -6218 496894
rect -6774 496338 -6538 496574
rect -6454 496338 -6218 496574
rect -6774 460658 -6538 460894
rect -6454 460658 -6218 460894
rect -6774 460338 -6538 460574
rect -6454 460338 -6218 460574
rect -6774 424658 -6538 424894
rect -6454 424658 -6218 424894
rect -6774 424338 -6538 424574
rect -6454 424338 -6218 424574
rect -6774 388658 -6538 388894
rect -6454 388658 -6218 388894
rect -6774 388338 -6538 388574
rect -6454 388338 -6218 388574
rect -6774 352658 -6538 352894
rect -6454 352658 -6218 352894
rect -6774 352338 -6538 352574
rect -6454 352338 -6218 352574
rect -6774 316658 -6538 316894
rect -6454 316658 -6218 316894
rect -6774 316338 -6538 316574
rect -6454 316338 -6218 316574
rect -6774 280658 -6538 280894
rect -6454 280658 -6218 280894
rect -6774 280338 -6538 280574
rect -6454 280338 -6218 280574
rect -6774 244658 -6538 244894
rect -6454 244658 -6218 244894
rect -6774 244338 -6538 244574
rect -6454 244338 -6218 244574
rect -6774 208658 -6538 208894
rect -6454 208658 -6218 208894
rect -6774 208338 -6538 208574
rect -6454 208338 -6218 208574
rect -6774 172658 -6538 172894
rect -6454 172658 -6218 172894
rect -6774 172338 -6538 172574
rect -6454 172338 -6218 172574
rect -6774 136658 -6538 136894
rect -6454 136658 -6218 136894
rect -6774 136338 -6538 136574
rect -6454 136338 -6218 136574
rect -6774 100658 -6538 100894
rect -6454 100658 -6218 100894
rect -6774 100338 -6538 100574
rect -6454 100338 -6218 100574
rect -6774 64658 -6538 64894
rect -6454 64658 -6218 64894
rect -6774 64338 -6538 64574
rect -6454 64338 -6218 64574
rect -6774 28658 -6538 28894
rect -6454 28658 -6218 28894
rect -6774 28338 -6538 28574
rect -6454 28338 -6218 28574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 9266 708442 9502 708678
rect 9586 708442 9822 708678
rect 9266 708122 9502 708358
rect 9586 708122 9822 708358
rect -5814 694658 -5578 694894
rect -5494 694658 -5258 694894
rect -5814 694338 -5578 694574
rect -5494 694338 -5258 694574
rect -5814 658658 -5578 658894
rect -5494 658658 -5258 658894
rect -5814 658338 -5578 658574
rect -5494 658338 -5258 658574
rect -5814 622658 -5578 622894
rect -5494 622658 -5258 622894
rect -5814 622338 -5578 622574
rect -5494 622338 -5258 622574
rect -5814 586658 -5578 586894
rect -5494 586658 -5258 586894
rect -5814 586338 -5578 586574
rect -5494 586338 -5258 586574
rect -5814 550658 -5578 550894
rect -5494 550658 -5258 550894
rect -5814 550338 -5578 550574
rect -5494 550338 -5258 550574
rect -5814 514658 -5578 514894
rect -5494 514658 -5258 514894
rect -5814 514338 -5578 514574
rect -5494 514338 -5258 514574
rect -5814 478658 -5578 478894
rect -5494 478658 -5258 478894
rect -5814 478338 -5578 478574
rect -5494 478338 -5258 478574
rect -5814 442658 -5578 442894
rect -5494 442658 -5258 442894
rect -5814 442338 -5578 442574
rect -5494 442338 -5258 442574
rect -5814 406658 -5578 406894
rect -5494 406658 -5258 406894
rect -5814 406338 -5578 406574
rect -5494 406338 -5258 406574
rect -5814 370658 -5578 370894
rect -5494 370658 -5258 370894
rect -5814 370338 -5578 370574
rect -5494 370338 -5258 370574
rect -5814 334658 -5578 334894
rect -5494 334658 -5258 334894
rect -5814 334338 -5578 334574
rect -5494 334338 -5258 334574
rect -5814 298658 -5578 298894
rect -5494 298658 -5258 298894
rect -5814 298338 -5578 298574
rect -5494 298338 -5258 298574
rect -5814 262658 -5578 262894
rect -5494 262658 -5258 262894
rect -5814 262338 -5578 262574
rect -5494 262338 -5258 262574
rect -5814 226658 -5578 226894
rect -5494 226658 -5258 226894
rect -5814 226338 -5578 226574
rect -5494 226338 -5258 226574
rect -5814 190658 -5578 190894
rect -5494 190658 -5258 190894
rect -5814 190338 -5578 190574
rect -5494 190338 -5258 190574
rect -5814 154658 -5578 154894
rect -5494 154658 -5258 154894
rect -5814 154338 -5578 154574
rect -5494 154338 -5258 154574
rect -5814 118658 -5578 118894
rect -5494 118658 -5258 118894
rect -5814 118338 -5578 118574
rect -5494 118338 -5258 118574
rect -5814 82658 -5578 82894
rect -5494 82658 -5258 82894
rect -5814 82338 -5578 82574
rect -5494 82338 -5258 82574
rect -5814 46658 -5578 46894
rect -5494 46658 -5258 46894
rect -5814 46338 -5578 46574
rect -5494 46338 -5258 46574
rect -5814 10658 -5578 10894
rect -5494 10658 -5258 10894
rect -5814 10338 -5578 10574
rect -5494 10338 -5258 10574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 672938 -4618 673174
rect -4534 672938 -4298 673174
rect -4854 672618 -4618 672854
rect -4534 672618 -4298 672854
rect -4854 636938 -4618 637174
rect -4534 636938 -4298 637174
rect -4854 636618 -4618 636854
rect -4534 636618 -4298 636854
rect -4854 600938 -4618 601174
rect -4534 600938 -4298 601174
rect -4854 600618 -4618 600854
rect -4534 600618 -4298 600854
rect -4854 564938 -4618 565174
rect -4534 564938 -4298 565174
rect -4854 564618 -4618 564854
rect -4534 564618 -4298 564854
rect -4854 528938 -4618 529174
rect -4534 528938 -4298 529174
rect -4854 528618 -4618 528854
rect -4534 528618 -4298 528854
rect -4854 492938 -4618 493174
rect -4534 492938 -4298 493174
rect -4854 492618 -4618 492854
rect -4534 492618 -4298 492854
rect -4854 456938 -4618 457174
rect -4534 456938 -4298 457174
rect -4854 456618 -4618 456854
rect -4534 456618 -4298 456854
rect -4854 420938 -4618 421174
rect -4534 420938 -4298 421174
rect -4854 420618 -4618 420854
rect -4534 420618 -4298 420854
rect -4854 384938 -4618 385174
rect -4534 384938 -4298 385174
rect -4854 384618 -4618 384854
rect -4534 384618 -4298 384854
rect -4854 348938 -4618 349174
rect -4534 348938 -4298 349174
rect -4854 348618 -4618 348854
rect -4534 348618 -4298 348854
rect -4854 312938 -4618 313174
rect -4534 312938 -4298 313174
rect -4854 312618 -4618 312854
rect -4534 312618 -4298 312854
rect -4854 276938 -4618 277174
rect -4534 276938 -4298 277174
rect -4854 276618 -4618 276854
rect -4534 276618 -4298 276854
rect -4854 240938 -4618 241174
rect -4534 240938 -4298 241174
rect -4854 240618 -4618 240854
rect -4534 240618 -4298 240854
rect -4854 204938 -4618 205174
rect -4534 204938 -4298 205174
rect -4854 204618 -4618 204854
rect -4534 204618 -4298 204854
rect -4854 168938 -4618 169174
rect -4534 168938 -4298 169174
rect -4854 168618 -4618 168854
rect -4534 168618 -4298 168854
rect -4854 132938 -4618 133174
rect -4534 132938 -4298 133174
rect -4854 132618 -4618 132854
rect -4534 132618 -4298 132854
rect -4854 96938 -4618 97174
rect -4534 96938 -4298 97174
rect -4854 96618 -4618 96854
rect -4534 96618 -4298 96854
rect -4854 60938 -4618 61174
rect -4534 60938 -4298 61174
rect -4854 60618 -4618 60854
rect -4534 60618 -4298 60854
rect -4854 24938 -4618 25174
rect -4534 24938 -4298 25174
rect -4854 24618 -4618 24854
rect -4534 24618 -4298 24854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 5546 706522 5782 706758
rect 5866 706522 6102 706758
rect 5546 706202 5782 706438
rect 5866 706202 6102 706438
rect -3894 690938 -3658 691174
rect -3574 690938 -3338 691174
rect -3894 690618 -3658 690854
rect -3574 690618 -3338 690854
rect -3894 654938 -3658 655174
rect -3574 654938 -3338 655174
rect -3894 654618 -3658 654854
rect -3574 654618 -3338 654854
rect -3894 618938 -3658 619174
rect -3574 618938 -3338 619174
rect -3894 618618 -3658 618854
rect -3574 618618 -3338 618854
rect -3894 582938 -3658 583174
rect -3574 582938 -3338 583174
rect -3894 582618 -3658 582854
rect -3574 582618 -3338 582854
rect -3894 546938 -3658 547174
rect -3574 546938 -3338 547174
rect -3894 546618 -3658 546854
rect -3574 546618 -3338 546854
rect -3894 510938 -3658 511174
rect -3574 510938 -3338 511174
rect -3894 510618 -3658 510854
rect -3574 510618 -3338 510854
rect -3894 474938 -3658 475174
rect -3574 474938 -3338 475174
rect -3894 474618 -3658 474854
rect -3574 474618 -3338 474854
rect -3894 438938 -3658 439174
rect -3574 438938 -3338 439174
rect -3894 438618 -3658 438854
rect -3574 438618 -3338 438854
rect -3894 402938 -3658 403174
rect -3574 402938 -3338 403174
rect -3894 402618 -3658 402854
rect -3574 402618 -3338 402854
rect -3894 366938 -3658 367174
rect -3574 366938 -3338 367174
rect -3894 366618 -3658 366854
rect -3574 366618 -3338 366854
rect -3894 330938 -3658 331174
rect -3574 330938 -3338 331174
rect -3894 330618 -3658 330854
rect -3574 330618 -3338 330854
rect -3894 294938 -3658 295174
rect -3574 294938 -3338 295174
rect -3894 294618 -3658 294854
rect -3574 294618 -3338 294854
rect -3894 258938 -3658 259174
rect -3574 258938 -3338 259174
rect -3894 258618 -3658 258854
rect -3574 258618 -3338 258854
rect -3894 222938 -3658 223174
rect -3574 222938 -3338 223174
rect -3894 222618 -3658 222854
rect -3574 222618 -3338 222854
rect -3894 186938 -3658 187174
rect -3574 186938 -3338 187174
rect -3894 186618 -3658 186854
rect -3574 186618 -3338 186854
rect -3894 150938 -3658 151174
rect -3574 150938 -3338 151174
rect -3894 150618 -3658 150854
rect -3574 150618 -3338 150854
rect -3894 114938 -3658 115174
rect -3574 114938 -3338 115174
rect -3894 114618 -3658 114854
rect -3574 114618 -3338 114854
rect -3894 78938 -3658 79174
rect -3574 78938 -3338 79174
rect -3894 78618 -3658 78854
rect -3574 78618 -3338 78854
rect -3894 42938 -3658 43174
rect -3574 42938 -3338 43174
rect -3894 42618 -3658 42854
rect -3574 42618 -3338 42854
rect -3894 6938 -3658 7174
rect -3574 6938 -3338 7174
rect -3894 6618 -3658 6854
rect -3574 6618 -3338 6854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 30986 711322 31222 711558
rect 31306 711322 31542 711558
rect 30986 711002 31222 711238
rect 31306 711002 31542 711238
rect 27266 709402 27502 709638
rect 27586 709402 27822 709638
rect 27266 709082 27502 709318
rect 27586 709082 27822 709318
rect 23546 707482 23782 707718
rect 23866 707482 24102 707718
rect 23546 707162 23782 707398
rect 23866 707162 24102 707398
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 48986 710362 49222 710598
rect 49306 710362 49542 710598
rect 48986 710042 49222 710278
rect 49306 710042 49542 710278
rect 45266 708442 45502 708678
rect 45586 708442 45822 708678
rect 45266 708122 45502 708358
rect 45586 708122 45822 708358
rect 41546 706522 41782 706758
rect 41866 706522 42102 706758
rect 41546 706202 41782 706438
rect 41866 706202 42102 706438
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 66986 711322 67222 711558
rect 67306 711322 67542 711558
rect 66986 711002 67222 711238
rect 67306 711002 67542 711238
rect 63266 709402 63502 709638
rect 63586 709402 63822 709638
rect 63266 709082 63502 709318
rect 63586 709082 63822 709318
rect 59546 707482 59782 707718
rect 59866 707482 60102 707718
rect 59546 707162 59782 707398
rect 59866 707162 60102 707398
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 84986 710362 85222 710598
rect 85306 710362 85542 710598
rect 84986 710042 85222 710278
rect 85306 710042 85542 710278
rect 81266 708442 81502 708678
rect 81586 708442 81822 708678
rect 81266 708122 81502 708358
rect 81586 708122 81822 708358
rect 77546 706522 77782 706758
rect 77866 706522 78102 706758
rect 77546 706202 77782 706438
rect 77866 706202 78102 706438
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 102986 711322 103222 711558
rect 103306 711322 103542 711558
rect 102986 711002 103222 711238
rect 103306 711002 103542 711238
rect 99266 709402 99502 709638
rect 99586 709402 99822 709638
rect 99266 709082 99502 709318
rect 99586 709082 99822 709318
rect 95546 707482 95782 707718
rect 95866 707482 96102 707718
rect 95546 707162 95782 707398
rect 95866 707162 96102 707398
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 120986 710362 121222 710598
rect 121306 710362 121542 710598
rect 120986 710042 121222 710278
rect 121306 710042 121542 710278
rect 117266 708442 117502 708678
rect 117586 708442 117822 708678
rect 117266 708122 117502 708358
rect 117586 708122 117822 708358
rect 113546 706522 113782 706758
rect 113866 706522 114102 706758
rect 113546 706202 113782 706438
rect 113866 706202 114102 706438
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 138986 711322 139222 711558
rect 139306 711322 139542 711558
rect 138986 711002 139222 711238
rect 139306 711002 139542 711238
rect 135266 709402 135502 709638
rect 135586 709402 135822 709638
rect 135266 709082 135502 709318
rect 135586 709082 135822 709318
rect 131546 707482 131782 707718
rect 131866 707482 132102 707718
rect 131546 707162 131782 707398
rect 131866 707162 132102 707398
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 156986 710362 157222 710598
rect 157306 710362 157542 710598
rect 156986 710042 157222 710278
rect 157306 710042 157542 710278
rect 153266 708442 153502 708678
rect 153586 708442 153822 708678
rect 153266 708122 153502 708358
rect 153586 708122 153822 708358
rect 149546 706522 149782 706758
rect 149866 706522 150102 706758
rect 149546 706202 149782 706438
rect 149866 706202 150102 706438
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 174986 711322 175222 711558
rect 175306 711322 175542 711558
rect 174986 711002 175222 711238
rect 175306 711002 175542 711238
rect 171266 709402 171502 709638
rect 171586 709402 171822 709638
rect 171266 709082 171502 709318
rect 171586 709082 171822 709318
rect 167546 707482 167782 707718
rect 167866 707482 168102 707718
rect 167546 707162 167782 707398
rect 167866 707162 168102 707398
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 192986 710362 193222 710598
rect 193306 710362 193542 710598
rect 192986 710042 193222 710278
rect 193306 710042 193542 710278
rect 189266 708442 189502 708678
rect 189586 708442 189822 708678
rect 189266 708122 189502 708358
rect 189586 708122 189822 708358
rect 185546 706522 185782 706758
rect 185866 706522 186102 706758
rect 185546 706202 185782 706438
rect 185866 706202 186102 706438
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 210986 711322 211222 711558
rect 211306 711322 211542 711558
rect 210986 711002 211222 711238
rect 211306 711002 211542 711238
rect 207266 709402 207502 709638
rect 207586 709402 207822 709638
rect 207266 709082 207502 709318
rect 207586 709082 207822 709318
rect 203546 707482 203782 707718
rect 203866 707482 204102 707718
rect 203546 707162 203782 707398
rect 203866 707162 204102 707398
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 228986 710362 229222 710598
rect 229306 710362 229542 710598
rect 228986 710042 229222 710278
rect 229306 710042 229542 710278
rect 225266 708442 225502 708678
rect 225586 708442 225822 708678
rect 225266 708122 225502 708358
rect 225586 708122 225822 708358
rect 221546 706522 221782 706758
rect 221866 706522 222102 706758
rect 221546 706202 221782 706438
rect 221866 706202 222102 706438
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 246986 711322 247222 711558
rect 247306 711322 247542 711558
rect 246986 711002 247222 711238
rect 247306 711002 247542 711238
rect 243266 709402 243502 709638
rect 243586 709402 243822 709638
rect 243266 709082 243502 709318
rect 243586 709082 243822 709318
rect 239546 707482 239782 707718
rect 239866 707482 240102 707718
rect 239546 707162 239782 707398
rect 239866 707162 240102 707398
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 264986 710362 265222 710598
rect 265306 710362 265542 710598
rect 264986 710042 265222 710278
rect 265306 710042 265542 710278
rect 261266 708442 261502 708678
rect 261586 708442 261822 708678
rect 261266 708122 261502 708358
rect 261586 708122 261822 708358
rect 257546 706522 257782 706758
rect 257866 706522 258102 706758
rect 257546 706202 257782 706438
rect 257866 706202 258102 706438
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 282986 711322 283222 711558
rect 283306 711322 283542 711558
rect 282986 711002 283222 711238
rect 283306 711002 283542 711238
rect 279266 709402 279502 709638
rect 279586 709402 279822 709638
rect 279266 709082 279502 709318
rect 279586 709082 279822 709318
rect 275546 707482 275782 707718
rect 275866 707482 276102 707718
rect 275546 707162 275782 707398
rect 275866 707162 276102 707398
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 300986 710362 301222 710598
rect 301306 710362 301542 710598
rect 300986 710042 301222 710278
rect 301306 710042 301542 710278
rect 297266 708442 297502 708678
rect 297586 708442 297822 708678
rect 297266 708122 297502 708358
rect 297586 708122 297822 708358
rect 293546 706522 293782 706758
rect 293866 706522 294102 706758
rect 293546 706202 293782 706438
rect 293866 706202 294102 706438
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 318986 711322 319222 711558
rect 319306 711322 319542 711558
rect 318986 711002 319222 711238
rect 319306 711002 319542 711238
rect 315266 709402 315502 709638
rect 315586 709402 315822 709638
rect 315266 709082 315502 709318
rect 315586 709082 315822 709318
rect 311546 707482 311782 707718
rect 311866 707482 312102 707718
rect 311546 707162 311782 707398
rect 311866 707162 312102 707398
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 336986 710362 337222 710598
rect 337306 710362 337542 710598
rect 336986 710042 337222 710278
rect 337306 710042 337542 710278
rect 333266 708442 333502 708678
rect 333586 708442 333822 708678
rect 333266 708122 333502 708358
rect 333586 708122 333822 708358
rect 329546 706522 329782 706758
rect 329866 706522 330102 706758
rect 329546 706202 329782 706438
rect 329866 706202 330102 706438
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 354986 711322 355222 711558
rect 355306 711322 355542 711558
rect 354986 711002 355222 711238
rect 355306 711002 355542 711238
rect 351266 709402 351502 709638
rect 351586 709402 351822 709638
rect 351266 709082 351502 709318
rect 351586 709082 351822 709318
rect 347546 707482 347782 707718
rect 347866 707482 348102 707718
rect 347546 707162 347782 707398
rect 347866 707162 348102 707398
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 372986 710362 373222 710598
rect 373306 710362 373542 710598
rect 372986 710042 373222 710278
rect 373306 710042 373542 710278
rect 369266 708442 369502 708678
rect 369586 708442 369822 708678
rect 369266 708122 369502 708358
rect 369586 708122 369822 708358
rect 365546 706522 365782 706758
rect 365866 706522 366102 706758
rect 365546 706202 365782 706438
rect 365866 706202 366102 706438
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 390986 711322 391222 711558
rect 391306 711322 391542 711558
rect 390986 711002 391222 711238
rect 391306 711002 391542 711238
rect 387266 709402 387502 709638
rect 387586 709402 387822 709638
rect 387266 709082 387502 709318
rect 387586 709082 387822 709318
rect 383546 707482 383782 707718
rect 383866 707482 384102 707718
rect 383546 707162 383782 707398
rect 383866 707162 384102 707398
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 408986 710362 409222 710598
rect 409306 710362 409542 710598
rect 408986 710042 409222 710278
rect 409306 710042 409542 710278
rect 405266 708442 405502 708678
rect 405586 708442 405822 708678
rect 405266 708122 405502 708358
rect 405586 708122 405822 708358
rect 401546 706522 401782 706758
rect 401866 706522 402102 706758
rect 401546 706202 401782 706438
rect 401866 706202 402102 706438
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 426986 711322 427222 711558
rect 427306 711322 427542 711558
rect 426986 711002 427222 711238
rect 427306 711002 427542 711238
rect 423266 709402 423502 709638
rect 423586 709402 423822 709638
rect 423266 709082 423502 709318
rect 423586 709082 423822 709318
rect 419546 707482 419782 707718
rect 419866 707482 420102 707718
rect 419546 707162 419782 707398
rect 419866 707162 420102 707398
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 444986 710362 445222 710598
rect 445306 710362 445542 710598
rect 444986 710042 445222 710278
rect 445306 710042 445542 710278
rect 441266 708442 441502 708678
rect 441586 708442 441822 708678
rect 441266 708122 441502 708358
rect 441586 708122 441822 708358
rect 437546 706522 437782 706758
rect 437866 706522 438102 706758
rect 437546 706202 437782 706438
rect 437866 706202 438102 706438
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 462986 711322 463222 711558
rect 463306 711322 463542 711558
rect 462986 711002 463222 711238
rect 463306 711002 463542 711238
rect 459266 709402 459502 709638
rect 459586 709402 459822 709638
rect 459266 709082 459502 709318
rect 459586 709082 459822 709318
rect 455546 707482 455782 707718
rect 455866 707482 456102 707718
rect 455546 707162 455782 707398
rect 455866 707162 456102 707398
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 480986 710362 481222 710598
rect 481306 710362 481542 710598
rect 480986 710042 481222 710278
rect 481306 710042 481542 710278
rect 477266 708442 477502 708678
rect 477586 708442 477822 708678
rect 477266 708122 477502 708358
rect 477586 708122 477822 708358
rect 473546 706522 473782 706758
rect 473866 706522 474102 706758
rect 473546 706202 473782 706438
rect 473866 706202 474102 706438
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 498986 711322 499222 711558
rect 499306 711322 499542 711558
rect 498986 711002 499222 711238
rect 499306 711002 499542 711238
rect 495266 709402 495502 709638
rect 495586 709402 495822 709638
rect 495266 709082 495502 709318
rect 495586 709082 495822 709318
rect 491546 707482 491782 707718
rect 491866 707482 492102 707718
rect 491546 707162 491782 707398
rect 491866 707162 492102 707398
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 516986 710362 517222 710598
rect 517306 710362 517542 710598
rect 516986 710042 517222 710278
rect 517306 710042 517542 710278
rect 513266 708442 513502 708678
rect 513586 708442 513822 708678
rect 513266 708122 513502 708358
rect 513586 708122 513822 708358
rect 509546 706522 509782 706758
rect 509866 706522 510102 706758
rect 509546 706202 509782 706438
rect 509866 706202 510102 706438
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 534986 711322 535222 711558
rect 535306 711322 535542 711558
rect 534986 711002 535222 711238
rect 535306 711002 535542 711238
rect 531266 709402 531502 709638
rect 531586 709402 531822 709638
rect 531266 709082 531502 709318
rect 531586 709082 531822 709318
rect 527546 707482 527782 707718
rect 527866 707482 528102 707718
rect 527546 707162 527782 707398
rect 527866 707162 528102 707398
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 552986 710362 553222 710598
rect 553306 710362 553542 710598
rect 552986 710042 553222 710278
rect 553306 710042 553542 710278
rect 549266 708442 549502 708678
rect 549586 708442 549822 708678
rect 549266 708122 549502 708358
rect 549586 708122 549822 708358
rect 545546 706522 545782 706758
rect 545866 706522 546102 706758
rect 545546 706202 545782 706438
rect 545866 706202 546102 706438
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 570986 711322 571222 711558
rect 571306 711322 571542 711558
rect 570986 711002 571222 711238
rect 571306 711002 571542 711238
rect 567266 709402 567502 709638
rect 567586 709402 567822 709638
rect 567266 709082 567502 709318
rect 567586 709082 567822 709318
rect 563546 707482 563782 707718
rect 563866 707482 564102 707718
rect 563546 707162 563782 707398
rect 563866 707162 564102 707398
rect 559826 705562 560062 705798
rect 560146 705562 560382 705798
rect 559826 705242 560062 705478
rect 560146 705242 560382 705478
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect 8250 687218 8486 687454
rect 8250 686898 8486 687134
rect 38970 687218 39206 687454
rect 38970 686898 39206 687134
rect 69690 687218 69926 687454
rect 69690 686898 69926 687134
rect 100410 687218 100646 687454
rect 100410 686898 100646 687134
rect 131130 687218 131366 687454
rect 131130 686898 131366 687134
rect 161850 687218 162086 687454
rect 161850 686898 162086 687134
rect 192570 687218 192806 687454
rect 192570 686898 192806 687134
rect 223290 687218 223526 687454
rect 223290 686898 223526 687134
rect 254010 687218 254246 687454
rect 254010 686898 254246 687134
rect 284730 687218 284966 687454
rect 284730 686898 284966 687134
rect 315450 687218 315686 687454
rect 315450 686898 315686 687134
rect 346170 687218 346406 687454
rect 346170 686898 346406 687134
rect 376890 687218 377126 687454
rect 376890 686898 377126 687134
rect 407610 687218 407846 687454
rect 407610 686898 407846 687134
rect 438330 687218 438566 687454
rect 438330 686898 438566 687134
rect 469050 687218 469286 687454
rect 469050 686898 469286 687134
rect 499770 687218 500006 687454
rect 499770 686898 500006 687134
rect 530490 687218 530726 687454
rect 530490 686898 530726 687134
rect 561210 687218 561446 687454
rect 561210 686898 561446 687134
rect 567266 676658 567502 676894
rect 567586 676658 567822 676894
rect 567266 676338 567502 676574
rect 567586 676338 567822 676574
rect 23610 669218 23846 669454
rect 23610 668898 23846 669134
rect 54330 669218 54566 669454
rect 54330 668898 54566 669134
rect 85050 669218 85286 669454
rect 85050 668898 85286 669134
rect 115770 669218 116006 669454
rect 115770 668898 116006 669134
rect 146490 669218 146726 669454
rect 146490 668898 146726 669134
rect 177210 669218 177446 669454
rect 177210 668898 177446 669134
rect 207930 669218 208166 669454
rect 207930 668898 208166 669134
rect 238650 669218 238886 669454
rect 238650 668898 238886 669134
rect 269370 669218 269606 669454
rect 269370 668898 269606 669134
rect 300090 669218 300326 669454
rect 300090 668898 300326 669134
rect 330810 669218 331046 669454
rect 330810 668898 331046 669134
rect 361530 669218 361766 669454
rect 361530 668898 361766 669134
rect 392250 669218 392486 669454
rect 392250 668898 392486 669134
rect 422970 669218 423206 669454
rect 422970 668898 423206 669134
rect 453690 669218 453926 669454
rect 453690 668898 453926 669134
rect 484410 669218 484646 669454
rect 484410 668898 484646 669134
rect 515130 669218 515366 669454
rect 515130 668898 515366 669134
rect 545850 669218 546086 669454
rect 545850 668898 546086 669134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect 8250 651218 8486 651454
rect 8250 650898 8486 651134
rect 38970 651218 39206 651454
rect 38970 650898 39206 651134
rect 69690 651218 69926 651454
rect 69690 650898 69926 651134
rect 100410 651218 100646 651454
rect 100410 650898 100646 651134
rect 131130 651218 131366 651454
rect 131130 650898 131366 651134
rect 161850 651218 162086 651454
rect 161850 650898 162086 651134
rect 192570 651218 192806 651454
rect 192570 650898 192806 651134
rect 223290 651218 223526 651454
rect 223290 650898 223526 651134
rect 254010 651218 254246 651454
rect 254010 650898 254246 651134
rect 284730 651218 284966 651454
rect 284730 650898 284966 651134
rect 315450 651218 315686 651454
rect 315450 650898 315686 651134
rect 346170 651218 346406 651454
rect 346170 650898 346406 651134
rect 376890 651218 377126 651454
rect 376890 650898 377126 651134
rect 407610 651218 407846 651454
rect 407610 650898 407846 651134
rect 438330 651218 438566 651454
rect 438330 650898 438566 651134
rect 469050 651218 469286 651454
rect 469050 650898 469286 651134
rect 499770 651218 500006 651454
rect 499770 650898 500006 651134
rect 530490 651218 530726 651454
rect 530490 650898 530726 651134
rect 561210 651218 561446 651454
rect 561210 650898 561446 651134
rect 567266 640658 567502 640894
rect 567586 640658 567822 640894
rect 567266 640338 567502 640574
rect 567586 640338 567822 640574
rect 23610 633218 23846 633454
rect 23610 632898 23846 633134
rect 54330 633218 54566 633454
rect 54330 632898 54566 633134
rect 85050 633218 85286 633454
rect 85050 632898 85286 633134
rect 115770 633218 116006 633454
rect 115770 632898 116006 633134
rect 146490 633218 146726 633454
rect 146490 632898 146726 633134
rect 177210 633218 177446 633454
rect 177210 632898 177446 633134
rect 207930 633218 208166 633454
rect 207930 632898 208166 633134
rect 238650 633218 238886 633454
rect 238650 632898 238886 633134
rect 269370 633218 269606 633454
rect 269370 632898 269606 633134
rect 300090 633218 300326 633454
rect 300090 632898 300326 633134
rect 330810 633218 331046 633454
rect 330810 632898 331046 633134
rect 361530 633218 361766 633454
rect 361530 632898 361766 633134
rect 392250 633218 392486 633454
rect 392250 632898 392486 633134
rect 422970 633218 423206 633454
rect 422970 632898 423206 633134
rect 453690 633218 453926 633454
rect 453690 632898 453926 633134
rect 484410 633218 484646 633454
rect 484410 632898 484646 633134
rect 515130 633218 515366 633454
rect 515130 632898 515366 633134
rect 545850 633218 546086 633454
rect 545850 632898 546086 633134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect 8250 615218 8486 615454
rect 8250 614898 8486 615134
rect 38970 615218 39206 615454
rect 38970 614898 39206 615134
rect 69690 615218 69926 615454
rect 69690 614898 69926 615134
rect 100410 615218 100646 615454
rect 100410 614898 100646 615134
rect 131130 615218 131366 615454
rect 131130 614898 131366 615134
rect 161850 615218 162086 615454
rect 161850 614898 162086 615134
rect 192570 615218 192806 615454
rect 192570 614898 192806 615134
rect 223290 615218 223526 615454
rect 223290 614898 223526 615134
rect 254010 615218 254246 615454
rect 254010 614898 254246 615134
rect 284730 615218 284966 615454
rect 284730 614898 284966 615134
rect 315450 615218 315686 615454
rect 315450 614898 315686 615134
rect 346170 615218 346406 615454
rect 346170 614898 346406 615134
rect 376890 615218 377126 615454
rect 376890 614898 377126 615134
rect 407610 615218 407846 615454
rect 407610 614898 407846 615134
rect 438330 615218 438566 615454
rect 438330 614898 438566 615134
rect 469050 615218 469286 615454
rect 469050 614898 469286 615134
rect 499770 615218 500006 615454
rect 499770 614898 500006 615134
rect 530490 615218 530726 615454
rect 530490 614898 530726 615134
rect 561210 615218 561446 615454
rect 561210 614898 561446 615134
rect 567266 604658 567502 604894
rect 567586 604658 567822 604894
rect 567266 604338 567502 604574
rect 567586 604338 567822 604574
rect 23610 597218 23846 597454
rect 23610 596898 23846 597134
rect 54330 597218 54566 597454
rect 54330 596898 54566 597134
rect 85050 597218 85286 597454
rect 85050 596898 85286 597134
rect 115770 597218 116006 597454
rect 115770 596898 116006 597134
rect 146490 597218 146726 597454
rect 146490 596898 146726 597134
rect 177210 597218 177446 597454
rect 177210 596898 177446 597134
rect 207930 597218 208166 597454
rect 207930 596898 208166 597134
rect 238650 597218 238886 597454
rect 238650 596898 238886 597134
rect 269370 597218 269606 597454
rect 269370 596898 269606 597134
rect 300090 597218 300326 597454
rect 300090 596898 300326 597134
rect 330810 597218 331046 597454
rect 330810 596898 331046 597134
rect 361530 597218 361766 597454
rect 361530 596898 361766 597134
rect 392250 597218 392486 597454
rect 392250 596898 392486 597134
rect 422970 597218 423206 597454
rect 422970 596898 423206 597134
rect 453690 597218 453926 597454
rect 453690 596898 453926 597134
rect 484410 597218 484646 597454
rect 484410 596898 484646 597134
rect 515130 597218 515366 597454
rect 515130 596898 515366 597134
rect 545850 597218 546086 597454
rect 545850 596898 546086 597134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect 8250 579218 8486 579454
rect 8250 578898 8486 579134
rect 38970 579218 39206 579454
rect 38970 578898 39206 579134
rect 69690 579218 69926 579454
rect 69690 578898 69926 579134
rect 100410 579218 100646 579454
rect 100410 578898 100646 579134
rect 131130 579218 131366 579454
rect 131130 578898 131366 579134
rect 161850 579218 162086 579454
rect 161850 578898 162086 579134
rect 192570 579218 192806 579454
rect 192570 578898 192806 579134
rect 223290 579218 223526 579454
rect 223290 578898 223526 579134
rect 254010 579218 254246 579454
rect 254010 578898 254246 579134
rect 284730 579218 284966 579454
rect 284730 578898 284966 579134
rect 315450 579218 315686 579454
rect 315450 578898 315686 579134
rect 346170 579218 346406 579454
rect 346170 578898 346406 579134
rect 376890 579218 377126 579454
rect 376890 578898 377126 579134
rect 407610 579218 407846 579454
rect 407610 578898 407846 579134
rect 438330 579218 438566 579454
rect 438330 578898 438566 579134
rect 469050 579218 469286 579454
rect 469050 578898 469286 579134
rect 499770 579218 500006 579454
rect 499770 578898 500006 579134
rect 530490 579218 530726 579454
rect 530490 578898 530726 579134
rect 561210 579218 561446 579454
rect 561210 578898 561446 579134
rect 567266 568658 567502 568894
rect 567586 568658 567822 568894
rect 567266 568338 567502 568574
rect 567586 568338 567822 568574
rect 23610 561218 23846 561454
rect 23610 560898 23846 561134
rect 54330 561218 54566 561454
rect 54330 560898 54566 561134
rect 85050 561218 85286 561454
rect 85050 560898 85286 561134
rect 115770 561218 116006 561454
rect 115770 560898 116006 561134
rect 146490 561218 146726 561454
rect 146490 560898 146726 561134
rect 177210 561218 177446 561454
rect 177210 560898 177446 561134
rect 207930 561218 208166 561454
rect 207930 560898 208166 561134
rect 238650 561218 238886 561454
rect 238650 560898 238886 561134
rect 269370 561218 269606 561454
rect 269370 560898 269606 561134
rect 300090 561218 300326 561454
rect 300090 560898 300326 561134
rect 330810 561218 331046 561454
rect 330810 560898 331046 561134
rect 361530 561218 361766 561454
rect 361530 560898 361766 561134
rect 392250 561218 392486 561454
rect 392250 560898 392486 561134
rect 422970 561218 423206 561454
rect 422970 560898 423206 561134
rect 453690 561218 453926 561454
rect 453690 560898 453926 561134
rect 484410 561218 484646 561454
rect 484410 560898 484646 561134
rect 515130 561218 515366 561454
rect 515130 560898 515366 561134
rect 545850 561218 546086 561454
rect 545850 560898 546086 561134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect 8250 543218 8486 543454
rect 8250 542898 8486 543134
rect 38970 543218 39206 543454
rect 38970 542898 39206 543134
rect 69690 543218 69926 543454
rect 69690 542898 69926 543134
rect 100410 543218 100646 543454
rect 100410 542898 100646 543134
rect 131130 543218 131366 543454
rect 131130 542898 131366 543134
rect 161850 543218 162086 543454
rect 161850 542898 162086 543134
rect 192570 543218 192806 543454
rect 192570 542898 192806 543134
rect 223290 543218 223526 543454
rect 223290 542898 223526 543134
rect 254010 543218 254246 543454
rect 254010 542898 254246 543134
rect 284730 543218 284966 543454
rect 284730 542898 284966 543134
rect 315450 543218 315686 543454
rect 315450 542898 315686 543134
rect 346170 543218 346406 543454
rect 346170 542898 346406 543134
rect 376890 543218 377126 543454
rect 376890 542898 377126 543134
rect 407610 543218 407846 543454
rect 407610 542898 407846 543134
rect 438330 543218 438566 543454
rect 438330 542898 438566 543134
rect 469050 543218 469286 543454
rect 469050 542898 469286 543134
rect 499770 543218 500006 543454
rect 499770 542898 500006 543134
rect 530490 543218 530726 543454
rect 530490 542898 530726 543134
rect 561210 543218 561446 543454
rect 561210 542898 561446 543134
rect 567266 532658 567502 532894
rect 567586 532658 567822 532894
rect 567266 532338 567502 532574
rect 567586 532338 567822 532574
rect 23610 525218 23846 525454
rect 23610 524898 23846 525134
rect 54330 525218 54566 525454
rect 54330 524898 54566 525134
rect 85050 525218 85286 525454
rect 85050 524898 85286 525134
rect 115770 525218 116006 525454
rect 115770 524898 116006 525134
rect 146490 525218 146726 525454
rect 146490 524898 146726 525134
rect 177210 525218 177446 525454
rect 177210 524898 177446 525134
rect 207930 525218 208166 525454
rect 207930 524898 208166 525134
rect 238650 525218 238886 525454
rect 238650 524898 238886 525134
rect 269370 525218 269606 525454
rect 269370 524898 269606 525134
rect 300090 525218 300326 525454
rect 300090 524898 300326 525134
rect 330810 525218 331046 525454
rect 330810 524898 331046 525134
rect 361530 525218 361766 525454
rect 361530 524898 361766 525134
rect 392250 525218 392486 525454
rect 392250 524898 392486 525134
rect 422970 525218 423206 525454
rect 422970 524898 423206 525134
rect 453690 525218 453926 525454
rect 453690 524898 453926 525134
rect 484410 525218 484646 525454
rect 484410 524898 484646 525134
rect 515130 525218 515366 525454
rect 515130 524898 515366 525134
rect 545850 525218 546086 525454
rect 545850 524898 546086 525134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect 8250 507218 8486 507454
rect 8250 506898 8486 507134
rect 38970 507218 39206 507454
rect 38970 506898 39206 507134
rect 69690 507218 69926 507454
rect 69690 506898 69926 507134
rect 100410 507218 100646 507454
rect 100410 506898 100646 507134
rect 131130 507218 131366 507454
rect 131130 506898 131366 507134
rect 161850 507218 162086 507454
rect 161850 506898 162086 507134
rect 192570 507218 192806 507454
rect 192570 506898 192806 507134
rect 223290 507218 223526 507454
rect 223290 506898 223526 507134
rect 254010 507218 254246 507454
rect 254010 506898 254246 507134
rect 284730 507218 284966 507454
rect 284730 506898 284966 507134
rect 315450 507218 315686 507454
rect 315450 506898 315686 507134
rect 346170 507218 346406 507454
rect 346170 506898 346406 507134
rect 376890 507218 377126 507454
rect 376890 506898 377126 507134
rect 407610 507218 407846 507454
rect 407610 506898 407846 507134
rect 438330 507218 438566 507454
rect 438330 506898 438566 507134
rect 469050 507218 469286 507454
rect 469050 506898 469286 507134
rect 499770 507218 500006 507454
rect 499770 506898 500006 507134
rect 530490 507218 530726 507454
rect 530490 506898 530726 507134
rect 561210 507218 561446 507454
rect 561210 506898 561446 507134
rect 567266 496658 567502 496894
rect 567586 496658 567822 496894
rect 567266 496338 567502 496574
rect 567586 496338 567822 496574
rect 23610 489218 23846 489454
rect 23610 488898 23846 489134
rect 54330 489218 54566 489454
rect 54330 488898 54566 489134
rect 85050 489218 85286 489454
rect 85050 488898 85286 489134
rect 115770 489218 116006 489454
rect 115770 488898 116006 489134
rect 146490 489218 146726 489454
rect 146490 488898 146726 489134
rect 177210 489218 177446 489454
rect 177210 488898 177446 489134
rect 207930 489218 208166 489454
rect 207930 488898 208166 489134
rect 238650 489218 238886 489454
rect 238650 488898 238886 489134
rect 269370 489218 269606 489454
rect 269370 488898 269606 489134
rect 300090 489218 300326 489454
rect 300090 488898 300326 489134
rect 330810 489218 331046 489454
rect 330810 488898 331046 489134
rect 361530 489218 361766 489454
rect 361530 488898 361766 489134
rect 392250 489218 392486 489454
rect 392250 488898 392486 489134
rect 422970 489218 423206 489454
rect 422970 488898 423206 489134
rect 453690 489218 453926 489454
rect 453690 488898 453926 489134
rect 484410 489218 484646 489454
rect 484410 488898 484646 489134
rect 515130 489218 515366 489454
rect 515130 488898 515366 489134
rect 545850 489218 546086 489454
rect 545850 488898 546086 489134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect 8250 471218 8486 471454
rect 8250 470898 8486 471134
rect 38970 471218 39206 471454
rect 38970 470898 39206 471134
rect 69690 471218 69926 471454
rect 69690 470898 69926 471134
rect 100410 471218 100646 471454
rect 100410 470898 100646 471134
rect 131130 471218 131366 471454
rect 131130 470898 131366 471134
rect 161850 471218 162086 471454
rect 161850 470898 162086 471134
rect 192570 471218 192806 471454
rect 192570 470898 192806 471134
rect 223290 471218 223526 471454
rect 223290 470898 223526 471134
rect 254010 471218 254246 471454
rect 254010 470898 254246 471134
rect 284730 471218 284966 471454
rect 284730 470898 284966 471134
rect 315450 471218 315686 471454
rect 315450 470898 315686 471134
rect 346170 471218 346406 471454
rect 346170 470898 346406 471134
rect 376890 471218 377126 471454
rect 376890 470898 377126 471134
rect 407610 471218 407846 471454
rect 407610 470898 407846 471134
rect 438330 471218 438566 471454
rect 438330 470898 438566 471134
rect 469050 471218 469286 471454
rect 469050 470898 469286 471134
rect 499770 471218 500006 471454
rect 499770 470898 500006 471134
rect 530490 471218 530726 471454
rect 530490 470898 530726 471134
rect 561210 471218 561446 471454
rect 561210 470898 561446 471134
rect 567266 460658 567502 460894
rect 567586 460658 567822 460894
rect 567266 460338 567502 460574
rect 567586 460338 567822 460574
rect 23610 453218 23846 453454
rect 23610 452898 23846 453134
rect 54330 453218 54566 453454
rect 54330 452898 54566 453134
rect 85050 453218 85286 453454
rect 85050 452898 85286 453134
rect 115770 453218 116006 453454
rect 115770 452898 116006 453134
rect 146490 453218 146726 453454
rect 146490 452898 146726 453134
rect 177210 453218 177446 453454
rect 177210 452898 177446 453134
rect 207930 453218 208166 453454
rect 207930 452898 208166 453134
rect 238650 453218 238886 453454
rect 238650 452898 238886 453134
rect 269370 453218 269606 453454
rect 269370 452898 269606 453134
rect 300090 453218 300326 453454
rect 300090 452898 300326 453134
rect 330810 453218 331046 453454
rect 330810 452898 331046 453134
rect 361530 453218 361766 453454
rect 361530 452898 361766 453134
rect 392250 453218 392486 453454
rect 392250 452898 392486 453134
rect 422970 453218 423206 453454
rect 422970 452898 423206 453134
rect 453690 453218 453926 453454
rect 453690 452898 453926 453134
rect 484410 453218 484646 453454
rect 484410 452898 484646 453134
rect 515130 453218 515366 453454
rect 515130 452898 515366 453134
rect 545850 453218 546086 453454
rect 545850 452898 546086 453134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect 8250 435218 8486 435454
rect 8250 434898 8486 435134
rect 38970 435218 39206 435454
rect 38970 434898 39206 435134
rect 69690 435218 69926 435454
rect 69690 434898 69926 435134
rect 100410 435218 100646 435454
rect 100410 434898 100646 435134
rect 131130 435218 131366 435454
rect 131130 434898 131366 435134
rect 161850 435218 162086 435454
rect 161850 434898 162086 435134
rect 192570 435218 192806 435454
rect 192570 434898 192806 435134
rect 223290 435218 223526 435454
rect 223290 434898 223526 435134
rect 254010 435218 254246 435454
rect 254010 434898 254246 435134
rect 284730 435218 284966 435454
rect 284730 434898 284966 435134
rect 315450 435218 315686 435454
rect 315450 434898 315686 435134
rect 346170 435218 346406 435454
rect 346170 434898 346406 435134
rect 376890 435218 377126 435454
rect 376890 434898 377126 435134
rect 407610 435218 407846 435454
rect 407610 434898 407846 435134
rect 438330 435218 438566 435454
rect 438330 434898 438566 435134
rect 469050 435218 469286 435454
rect 469050 434898 469286 435134
rect 499770 435218 500006 435454
rect 499770 434898 500006 435134
rect 530490 435218 530726 435454
rect 530490 434898 530726 435134
rect 561210 435218 561446 435454
rect 561210 434898 561446 435134
rect 567266 424658 567502 424894
rect 567586 424658 567822 424894
rect 567266 424338 567502 424574
rect 567586 424338 567822 424574
rect 23610 417218 23846 417454
rect 23610 416898 23846 417134
rect 54330 417218 54566 417454
rect 54330 416898 54566 417134
rect 85050 417218 85286 417454
rect 85050 416898 85286 417134
rect 115770 417218 116006 417454
rect 115770 416898 116006 417134
rect 146490 417218 146726 417454
rect 146490 416898 146726 417134
rect 177210 417218 177446 417454
rect 177210 416898 177446 417134
rect 207930 417218 208166 417454
rect 207930 416898 208166 417134
rect 238650 417218 238886 417454
rect 238650 416898 238886 417134
rect 269370 417218 269606 417454
rect 269370 416898 269606 417134
rect 300090 417218 300326 417454
rect 300090 416898 300326 417134
rect 330810 417218 331046 417454
rect 330810 416898 331046 417134
rect 361530 417218 361766 417454
rect 361530 416898 361766 417134
rect 392250 417218 392486 417454
rect 392250 416898 392486 417134
rect 422970 417218 423206 417454
rect 422970 416898 423206 417134
rect 453690 417218 453926 417454
rect 453690 416898 453926 417134
rect 484410 417218 484646 417454
rect 484410 416898 484646 417134
rect 515130 417218 515366 417454
rect 515130 416898 515366 417134
rect 545850 417218 546086 417454
rect 545850 416898 546086 417134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect 8250 399218 8486 399454
rect 8250 398898 8486 399134
rect 38970 399218 39206 399454
rect 38970 398898 39206 399134
rect 69690 399218 69926 399454
rect 69690 398898 69926 399134
rect 100410 399218 100646 399454
rect 100410 398898 100646 399134
rect 131130 399218 131366 399454
rect 131130 398898 131366 399134
rect 161850 399218 162086 399454
rect 161850 398898 162086 399134
rect 192570 399218 192806 399454
rect 192570 398898 192806 399134
rect 223290 399218 223526 399454
rect 223290 398898 223526 399134
rect 254010 399218 254246 399454
rect 254010 398898 254246 399134
rect 284730 399218 284966 399454
rect 284730 398898 284966 399134
rect 315450 399218 315686 399454
rect 315450 398898 315686 399134
rect 346170 399218 346406 399454
rect 346170 398898 346406 399134
rect 376890 399218 377126 399454
rect 376890 398898 377126 399134
rect 407610 399218 407846 399454
rect 407610 398898 407846 399134
rect 438330 399218 438566 399454
rect 438330 398898 438566 399134
rect 469050 399218 469286 399454
rect 469050 398898 469286 399134
rect 499770 399218 500006 399454
rect 499770 398898 500006 399134
rect 530490 399218 530726 399454
rect 530490 398898 530726 399134
rect 561210 399218 561446 399454
rect 561210 398898 561446 399134
rect 567266 388658 567502 388894
rect 567586 388658 567822 388894
rect 567266 388338 567502 388574
rect 567586 388338 567822 388574
rect 23610 381218 23846 381454
rect 23610 380898 23846 381134
rect 54330 381218 54566 381454
rect 54330 380898 54566 381134
rect 85050 381218 85286 381454
rect 85050 380898 85286 381134
rect 115770 381218 116006 381454
rect 115770 380898 116006 381134
rect 146490 381218 146726 381454
rect 146490 380898 146726 381134
rect 177210 381218 177446 381454
rect 177210 380898 177446 381134
rect 207930 381218 208166 381454
rect 207930 380898 208166 381134
rect 238650 381218 238886 381454
rect 238650 380898 238886 381134
rect 269370 381218 269606 381454
rect 269370 380898 269606 381134
rect 300090 381218 300326 381454
rect 300090 380898 300326 381134
rect 330810 381218 331046 381454
rect 330810 380898 331046 381134
rect 361530 381218 361766 381454
rect 361530 380898 361766 381134
rect 392250 381218 392486 381454
rect 392250 380898 392486 381134
rect 422970 381218 423206 381454
rect 422970 380898 423206 381134
rect 453690 381218 453926 381454
rect 453690 380898 453926 381134
rect 484410 381218 484646 381454
rect 484410 380898 484646 381134
rect 515130 381218 515366 381454
rect 515130 380898 515366 381134
rect 545850 381218 546086 381454
rect 545850 380898 546086 381134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect 8250 363218 8486 363454
rect 8250 362898 8486 363134
rect 38970 363218 39206 363454
rect 38970 362898 39206 363134
rect 69690 363218 69926 363454
rect 69690 362898 69926 363134
rect 100410 363218 100646 363454
rect 100410 362898 100646 363134
rect 131130 363218 131366 363454
rect 131130 362898 131366 363134
rect 161850 363218 162086 363454
rect 161850 362898 162086 363134
rect 192570 363218 192806 363454
rect 192570 362898 192806 363134
rect 223290 363218 223526 363454
rect 223290 362898 223526 363134
rect 254010 363218 254246 363454
rect 254010 362898 254246 363134
rect 284730 363218 284966 363454
rect 284730 362898 284966 363134
rect 315450 363218 315686 363454
rect 315450 362898 315686 363134
rect 346170 363218 346406 363454
rect 346170 362898 346406 363134
rect 376890 363218 377126 363454
rect 376890 362898 377126 363134
rect 407610 363218 407846 363454
rect 407610 362898 407846 363134
rect 438330 363218 438566 363454
rect 438330 362898 438566 363134
rect 469050 363218 469286 363454
rect 469050 362898 469286 363134
rect 499770 363218 500006 363454
rect 499770 362898 500006 363134
rect 530490 363218 530726 363454
rect 530490 362898 530726 363134
rect 561210 363218 561446 363454
rect 561210 362898 561446 363134
rect 567266 352658 567502 352894
rect 567586 352658 567822 352894
rect 567266 352338 567502 352574
rect 567586 352338 567822 352574
rect 23610 345218 23846 345454
rect 23610 344898 23846 345134
rect 54330 345218 54566 345454
rect 54330 344898 54566 345134
rect 85050 345218 85286 345454
rect 85050 344898 85286 345134
rect 115770 345218 116006 345454
rect 115770 344898 116006 345134
rect 146490 345218 146726 345454
rect 146490 344898 146726 345134
rect 177210 345218 177446 345454
rect 177210 344898 177446 345134
rect 207930 345218 208166 345454
rect 207930 344898 208166 345134
rect 238650 345218 238886 345454
rect 238650 344898 238886 345134
rect 269370 345218 269606 345454
rect 269370 344898 269606 345134
rect 300090 345218 300326 345454
rect 300090 344898 300326 345134
rect 330810 345218 331046 345454
rect 330810 344898 331046 345134
rect 361530 345218 361766 345454
rect 361530 344898 361766 345134
rect 392250 345218 392486 345454
rect 392250 344898 392486 345134
rect 422970 345218 423206 345454
rect 422970 344898 423206 345134
rect 453690 345218 453926 345454
rect 453690 344898 453926 345134
rect 484410 345218 484646 345454
rect 484410 344898 484646 345134
rect 515130 345218 515366 345454
rect 515130 344898 515366 345134
rect 545850 345218 546086 345454
rect 545850 344898 546086 345134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect 8250 327218 8486 327454
rect 8250 326898 8486 327134
rect 38970 327218 39206 327454
rect 38970 326898 39206 327134
rect 69690 327218 69926 327454
rect 69690 326898 69926 327134
rect 100410 327218 100646 327454
rect 100410 326898 100646 327134
rect 131130 327218 131366 327454
rect 131130 326898 131366 327134
rect 161850 327218 162086 327454
rect 161850 326898 162086 327134
rect 192570 327218 192806 327454
rect 192570 326898 192806 327134
rect 223290 327218 223526 327454
rect 223290 326898 223526 327134
rect 254010 327218 254246 327454
rect 254010 326898 254246 327134
rect 284730 327218 284966 327454
rect 284730 326898 284966 327134
rect 315450 327218 315686 327454
rect 315450 326898 315686 327134
rect 346170 327218 346406 327454
rect 346170 326898 346406 327134
rect 376890 327218 377126 327454
rect 376890 326898 377126 327134
rect 407610 327218 407846 327454
rect 407610 326898 407846 327134
rect 438330 327218 438566 327454
rect 438330 326898 438566 327134
rect 469050 327218 469286 327454
rect 469050 326898 469286 327134
rect 499770 327218 500006 327454
rect 499770 326898 500006 327134
rect 530490 327218 530726 327454
rect 530490 326898 530726 327134
rect 561210 327218 561446 327454
rect 561210 326898 561446 327134
rect 567266 316658 567502 316894
rect 567586 316658 567822 316894
rect 567266 316338 567502 316574
rect 567586 316338 567822 316574
rect 23610 309218 23846 309454
rect 23610 308898 23846 309134
rect 54330 309218 54566 309454
rect 54330 308898 54566 309134
rect 85050 309218 85286 309454
rect 85050 308898 85286 309134
rect 115770 309218 116006 309454
rect 115770 308898 116006 309134
rect 146490 309218 146726 309454
rect 146490 308898 146726 309134
rect 177210 309218 177446 309454
rect 177210 308898 177446 309134
rect 207930 309218 208166 309454
rect 207930 308898 208166 309134
rect 238650 309218 238886 309454
rect 238650 308898 238886 309134
rect 269370 309218 269606 309454
rect 269370 308898 269606 309134
rect 300090 309218 300326 309454
rect 300090 308898 300326 309134
rect 330810 309218 331046 309454
rect 330810 308898 331046 309134
rect 361530 309218 361766 309454
rect 361530 308898 361766 309134
rect 392250 309218 392486 309454
rect 392250 308898 392486 309134
rect 422970 309218 423206 309454
rect 422970 308898 423206 309134
rect 453690 309218 453926 309454
rect 453690 308898 453926 309134
rect 484410 309218 484646 309454
rect 484410 308898 484646 309134
rect 515130 309218 515366 309454
rect 515130 308898 515366 309134
rect 545850 309218 546086 309454
rect 545850 308898 546086 309134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect 8250 291218 8486 291454
rect 8250 290898 8486 291134
rect 38970 291218 39206 291454
rect 38970 290898 39206 291134
rect 69690 291218 69926 291454
rect 69690 290898 69926 291134
rect 100410 291218 100646 291454
rect 100410 290898 100646 291134
rect 131130 291218 131366 291454
rect 131130 290898 131366 291134
rect 161850 291218 162086 291454
rect 161850 290898 162086 291134
rect 192570 291218 192806 291454
rect 192570 290898 192806 291134
rect 223290 291218 223526 291454
rect 223290 290898 223526 291134
rect 254010 291218 254246 291454
rect 254010 290898 254246 291134
rect 284730 291218 284966 291454
rect 284730 290898 284966 291134
rect 315450 291218 315686 291454
rect 315450 290898 315686 291134
rect 346170 291218 346406 291454
rect 346170 290898 346406 291134
rect 376890 291218 377126 291454
rect 376890 290898 377126 291134
rect 407610 291218 407846 291454
rect 407610 290898 407846 291134
rect 438330 291218 438566 291454
rect 438330 290898 438566 291134
rect 469050 291218 469286 291454
rect 469050 290898 469286 291134
rect 499770 291218 500006 291454
rect 499770 290898 500006 291134
rect 530490 291218 530726 291454
rect 530490 290898 530726 291134
rect 561210 291218 561446 291454
rect 561210 290898 561446 291134
rect 567266 280658 567502 280894
rect 567586 280658 567822 280894
rect 567266 280338 567502 280574
rect 567586 280338 567822 280574
rect 23610 273218 23846 273454
rect 23610 272898 23846 273134
rect 54330 273218 54566 273454
rect 54330 272898 54566 273134
rect 85050 273218 85286 273454
rect 85050 272898 85286 273134
rect 115770 273218 116006 273454
rect 115770 272898 116006 273134
rect 146490 273218 146726 273454
rect 146490 272898 146726 273134
rect 177210 273218 177446 273454
rect 177210 272898 177446 273134
rect 207930 273218 208166 273454
rect 207930 272898 208166 273134
rect 238650 273218 238886 273454
rect 238650 272898 238886 273134
rect 269370 273218 269606 273454
rect 269370 272898 269606 273134
rect 300090 273218 300326 273454
rect 300090 272898 300326 273134
rect 330810 273218 331046 273454
rect 330810 272898 331046 273134
rect 361530 273218 361766 273454
rect 361530 272898 361766 273134
rect 392250 273218 392486 273454
rect 392250 272898 392486 273134
rect 422970 273218 423206 273454
rect 422970 272898 423206 273134
rect 453690 273218 453926 273454
rect 453690 272898 453926 273134
rect 484410 273218 484646 273454
rect 484410 272898 484646 273134
rect 515130 273218 515366 273454
rect 515130 272898 515366 273134
rect 545850 273218 546086 273454
rect 545850 272898 546086 273134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect 8250 255218 8486 255454
rect 8250 254898 8486 255134
rect 38970 255218 39206 255454
rect 38970 254898 39206 255134
rect 69690 255218 69926 255454
rect 69690 254898 69926 255134
rect 100410 255218 100646 255454
rect 100410 254898 100646 255134
rect 131130 255218 131366 255454
rect 131130 254898 131366 255134
rect 161850 255218 162086 255454
rect 161850 254898 162086 255134
rect 192570 255218 192806 255454
rect 192570 254898 192806 255134
rect 223290 255218 223526 255454
rect 223290 254898 223526 255134
rect 254010 255218 254246 255454
rect 254010 254898 254246 255134
rect 284730 255218 284966 255454
rect 284730 254898 284966 255134
rect 315450 255218 315686 255454
rect 315450 254898 315686 255134
rect 346170 255218 346406 255454
rect 346170 254898 346406 255134
rect 376890 255218 377126 255454
rect 376890 254898 377126 255134
rect 407610 255218 407846 255454
rect 407610 254898 407846 255134
rect 438330 255218 438566 255454
rect 438330 254898 438566 255134
rect 469050 255218 469286 255454
rect 469050 254898 469286 255134
rect 499770 255218 500006 255454
rect 499770 254898 500006 255134
rect 530490 255218 530726 255454
rect 530490 254898 530726 255134
rect 561210 255218 561446 255454
rect 561210 254898 561446 255134
rect 567266 244658 567502 244894
rect 567586 244658 567822 244894
rect 567266 244338 567502 244574
rect 567586 244338 567822 244574
rect 23610 237218 23846 237454
rect 23610 236898 23846 237134
rect 54330 237218 54566 237454
rect 54330 236898 54566 237134
rect 85050 237218 85286 237454
rect 85050 236898 85286 237134
rect 115770 237218 116006 237454
rect 115770 236898 116006 237134
rect 146490 237218 146726 237454
rect 146490 236898 146726 237134
rect 177210 237218 177446 237454
rect 177210 236898 177446 237134
rect 207930 237218 208166 237454
rect 207930 236898 208166 237134
rect 238650 237218 238886 237454
rect 238650 236898 238886 237134
rect 269370 237218 269606 237454
rect 269370 236898 269606 237134
rect 300090 237218 300326 237454
rect 300090 236898 300326 237134
rect 330810 237218 331046 237454
rect 330810 236898 331046 237134
rect 361530 237218 361766 237454
rect 361530 236898 361766 237134
rect 392250 237218 392486 237454
rect 392250 236898 392486 237134
rect 422970 237218 423206 237454
rect 422970 236898 423206 237134
rect 453690 237218 453926 237454
rect 453690 236898 453926 237134
rect 484410 237218 484646 237454
rect 484410 236898 484646 237134
rect 515130 237218 515366 237454
rect 515130 236898 515366 237134
rect 545850 237218 546086 237454
rect 545850 236898 546086 237134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect 8250 219218 8486 219454
rect 8250 218898 8486 219134
rect 38970 219218 39206 219454
rect 38970 218898 39206 219134
rect 69690 219218 69926 219454
rect 69690 218898 69926 219134
rect 100410 219218 100646 219454
rect 100410 218898 100646 219134
rect 131130 219218 131366 219454
rect 131130 218898 131366 219134
rect 161850 219218 162086 219454
rect 161850 218898 162086 219134
rect 192570 219218 192806 219454
rect 192570 218898 192806 219134
rect 223290 219218 223526 219454
rect 223290 218898 223526 219134
rect 254010 219218 254246 219454
rect 254010 218898 254246 219134
rect 284730 219218 284966 219454
rect 284730 218898 284966 219134
rect 315450 219218 315686 219454
rect 315450 218898 315686 219134
rect 346170 219218 346406 219454
rect 346170 218898 346406 219134
rect 376890 219218 377126 219454
rect 376890 218898 377126 219134
rect 407610 219218 407846 219454
rect 407610 218898 407846 219134
rect 438330 219218 438566 219454
rect 438330 218898 438566 219134
rect 469050 219218 469286 219454
rect 469050 218898 469286 219134
rect 499770 219218 500006 219454
rect 499770 218898 500006 219134
rect 530490 219218 530726 219454
rect 530490 218898 530726 219134
rect 561210 219218 561446 219454
rect 561210 218898 561446 219134
rect 567266 208658 567502 208894
rect 567586 208658 567822 208894
rect 567266 208338 567502 208574
rect 567586 208338 567822 208574
rect 23610 201218 23846 201454
rect 23610 200898 23846 201134
rect 54330 201218 54566 201454
rect 54330 200898 54566 201134
rect 85050 201218 85286 201454
rect 85050 200898 85286 201134
rect 115770 201218 116006 201454
rect 115770 200898 116006 201134
rect 146490 201218 146726 201454
rect 146490 200898 146726 201134
rect 177210 201218 177446 201454
rect 177210 200898 177446 201134
rect 207930 201218 208166 201454
rect 207930 200898 208166 201134
rect 238650 201218 238886 201454
rect 238650 200898 238886 201134
rect 269370 201218 269606 201454
rect 269370 200898 269606 201134
rect 300090 201218 300326 201454
rect 300090 200898 300326 201134
rect 330810 201218 331046 201454
rect 330810 200898 331046 201134
rect 361530 201218 361766 201454
rect 361530 200898 361766 201134
rect 392250 201218 392486 201454
rect 392250 200898 392486 201134
rect 422970 201218 423206 201454
rect 422970 200898 423206 201134
rect 453690 201218 453926 201454
rect 453690 200898 453926 201134
rect 484410 201218 484646 201454
rect 484410 200898 484646 201134
rect 515130 201218 515366 201454
rect 515130 200898 515366 201134
rect 545850 201218 546086 201454
rect 545850 200898 546086 201134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect 8250 183218 8486 183454
rect 8250 182898 8486 183134
rect 38970 183218 39206 183454
rect 38970 182898 39206 183134
rect 69690 183218 69926 183454
rect 69690 182898 69926 183134
rect 100410 183218 100646 183454
rect 100410 182898 100646 183134
rect 131130 183218 131366 183454
rect 131130 182898 131366 183134
rect 161850 183218 162086 183454
rect 161850 182898 162086 183134
rect 192570 183218 192806 183454
rect 192570 182898 192806 183134
rect 223290 183218 223526 183454
rect 223290 182898 223526 183134
rect 254010 183218 254246 183454
rect 254010 182898 254246 183134
rect 284730 183218 284966 183454
rect 284730 182898 284966 183134
rect 315450 183218 315686 183454
rect 315450 182898 315686 183134
rect 346170 183218 346406 183454
rect 346170 182898 346406 183134
rect 376890 183218 377126 183454
rect 376890 182898 377126 183134
rect 407610 183218 407846 183454
rect 407610 182898 407846 183134
rect 438330 183218 438566 183454
rect 438330 182898 438566 183134
rect 469050 183218 469286 183454
rect 469050 182898 469286 183134
rect 499770 183218 500006 183454
rect 499770 182898 500006 183134
rect 530490 183218 530726 183454
rect 530490 182898 530726 183134
rect 561210 183218 561446 183454
rect 561210 182898 561446 183134
rect 567266 172658 567502 172894
rect 567586 172658 567822 172894
rect 567266 172338 567502 172574
rect 567586 172338 567822 172574
rect 23610 165218 23846 165454
rect 23610 164898 23846 165134
rect 54330 165218 54566 165454
rect 54330 164898 54566 165134
rect 85050 165218 85286 165454
rect 85050 164898 85286 165134
rect 115770 165218 116006 165454
rect 115770 164898 116006 165134
rect 146490 165218 146726 165454
rect 146490 164898 146726 165134
rect 177210 165218 177446 165454
rect 177210 164898 177446 165134
rect 207930 165218 208166 165454
rect 207930 164898 208166 165134
rect 238650 165218 238886 165454
rect 238650 164898 238886 165134
rect 269370 165218 269606 165454
rect 269370 164898 269606 165134
rect 300090 165218 300326 165454
rect 300090 164898 300326 165134
rect 330810 165218 331046 165454
rect 330810 164898 331046 165134
rect 361530 165218 361766 165454
rect 361530 164898 361766 165134
rect 392250 165218 392486 165454
rect 392250 164898 392486 165134
rect 422970 165218 423206 165454
rect 422970 164898 423206 165134
rect 453690 165218 453926 165454
rect 453690 164898 453926 165134
rect 484410 165218 484646 165454
rect 484410 164898 484646 165134
rect 515130 165218 515366 165454
rect 515130 164898 515366 165134
rect 545850 165218 546086 165454
rect 545850 164898 546086 165134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect 8250 147218 8486 147454
rect 8250 146898 8486 147134
rect 38970 147218 39206 147454
rect 38970 146898 39206 147134
rect 69690 147218 69926 147454
rect 69690 146898 69926 147134
rect 100410 147218 100646 147454
rect 100410 146898 100646 147134
rect 131130 147218 131366 147454
rect 131130 146898 131366 147134
rect 161850 147218 162086 147454
rect 161850 146898 162086 147134
rect 192570 147218 192806 147454
rect 192570 146898 192806 147134
rect 223290 147218 223526 147454
rect 223290 146898 223526 147134
rect 254010 147218 254246 147454
rect 254010 146898 254246 147134
rect 284730 147218 284966 147454
rect 284730 146898 284966 147134
rect 315450 147218 315686 147454
rect 315450 146898 315686 147134
rect 346170 147218 346406 147454
rect 346170 146898 346406 147134
rect 376890 147218 377126 147454
rect 376890 146898 377126 147134
rect 407610 147218 407846 147454
rect 407610 146898 407846 147134
rect 438330 147218 438566 147454
rect 438330 146898 438566 147134
rect 469050 147218 469286 147454
rect 469050 146898 469286 147134
rect 499770 147218 500006 147454
rect 499770 146898 500006 147134
rect 530490 147218 530726 147454
rect 530490 146898 530726 147134
rect 561210 147218 561446 147454
rect 561210 146898 561446 147134
rect 567266 136658 567502 136894
rect 567586 136658 567822 136894
rect 567266 136338 567502 136574
rect 567586 136338 567822 136574
rect 23610 129218 23846 129454
rect 23610 128898 23846 129134
rect 54330 129218 54566 129454
rect 54330 128898 54566 129134
rect 85050 129218 85286 129454
rect 85050 128898 85286 129134
rect 115770 129218 116006 129454
rect 115770 128898 116006 129134
rect 146490 129218 146726 129454
rect 146490 128898 146726 129134
rect 177210 129218 177446 129454
rect 177210 128898 177446 129134
rect 207930 129218 208166 129454
rect 207930 128898 208166 129134
rect 238650 129218 238886 129454
rect 238650 128898 238886 129134
rect 269370 129218 269606 129454
rect 269370 128898 269606 129134
rect 300090 129218 300326 129454
rect 300090 128898 300326 129134
rect 330810 129218 331046 129454
rect 330810 128898 331046 129134
rect 361530 129218 361766 129454
rect 361530 128898 361766 129134
rect 392250 129218 392486 129454
rect 392250 128898 392486 129134
rect 422970 129218 423206 129454
rect 422970 128898 423206 129134
rect 453690 129218 453926 129454
rect 453690 128898 453926 129134
rect 484410 129218 484646 129454
rect 484410 128898 484646 129134
rect 515130 129218 515366 129454
rect 515130 128898 515366 129134
rect 545850 129218 546086 129454
rect 545850 128898 546086 129134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect 8250 111218 8486 111454
rect 8250 110898 8486 111134
rect 38970 111218 39206 111454
rect 38970 110898 39206 111134
rect 69690 111218 69926 111454
rect 69690 110898 69926 111134
rect 100410 111218 100646 111454
rect 100410 110898 100646 111134
rect 131130 111218 131366 111454
rect 131130 110898 131366 111134
rect 161850 111218 162086 111454
rect 161850 110898 162086 111134
rect 192570 111218 192806 111454
rect 192570 110898 192806 111134
rect 223290 111218 223526 111454
rect 223290 110898 223526 111134
rect 254010 111218 254246 111454
rect 254010 110898 254246 111134
rect 284730 111218 284966 111454
rect 284730 110898 284966 111134
rect 315450 111218 315686 111454
rect 315450 110898 315686 111134
rect 346170 111218 346406 111454
rect 346170 110898 346406 111134
rect 376890 111218 377126 111454
rect 376890 110898 377126 111134
rect 407610 111218 407846 111454
rect 407610 110898 407846 111134
rect 438330 111218 438566 111454
rect 438330 110898 438566 111134
rect 469050 111218 469286 111454
rect 469050 110898 469286 111134
rect 499770 111218 500006 111454
rect 499770 110898 500006 111134
rect 530490 111218 530726 111454
rect 530490 110898 530726 111134
rect 561210 111218 561446 111454
rect 561210 110898 561446 111134
rect 567266 100658 567502 100894
rect 567586 100658 567822 100894
rect 567266 100338 567502 100574
rect 567586 100338 567822 100574
rect 23610 93218 23846 93454
rect 23610 92898 23846 93134
rect 54330 93218 54566 93454
rect 54330 92898 54566 93134
rect 85050 93218 85286 93454
rect 85050 92898 85286 93134
rect 115770 93218 116006 93454
rect 115770 92898 116006 93134
rect 146490 93218 146726 93454
rect 146490 92898 146726 93134
rect 177210 93218 177446 93454
rect 177210 92898 177446 93134
rect 207930 93218 208166 93454
rect 207930 92898 208166 93134
rect 238650 93218 238886 93454
rect 238650 92898 238886 93134
rect 269370 93218 269606 93454
rect 269370 92898 269606 93134
rect 300090 93218 300326 93454
rect 300090 92898 300326 93134
rect 330810 93218 331046 93454
rect 330810 92898 331046 93134
rect 361530 93218 361766 93454
rect 361530 92898 361766 93134
rect 392250 93218 392486 93454
rect 392250 92898 392486 93134
rect 422970 93218 423206 93454
rect 422970 92898 423206 93134
rect 453690 93218 453926 93454
rect 453690 92898 453926 93134
rect 484410 93218 484646 93454
rect 484410 92898 484646 93134
rect 515130 93218 515366 93454
rect 515130 92898 515366 93134
rect 545850 93218 546086 93454
rect 545850 92898 546086 93134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect 8250 75218 8486 75454
rect 8250 74898 8486 75134
rect 38970 75218 39206 75454
rect 38970 74898 39206 75134
rect 69690 75218 69926 75454
rect 69690 74898 69926 75134
rect 100410 75218 100646 75454
rect 100410 74898 100646 75134
rect 131130 75218 131366 75454
rect 131130 74898 131366 75134
rect 161850 75218 162086 75454
rect 161850 74898 162086 75134
rect 192570 75218 192806 75454
rect 192570 74898 192806 75134
rect 223290 75218 223526 75454
rect 223290 74898 223526 75134
rect 254010 75218 254246 75454
rect 254010 74898 254246 75134
rect 284730 75218 284966 75454
rect 284730 74898 284966 75134
rect 315450 75218 315686 75454
rect 315450 74898 315686 75134
rect 346170 75218 346406 75454
rect 346170 74898 346406 75134
rect 376890 75218 377126 75454
rect 376890 74898 377126 75134
rect 407610 75218 407846 75454
rect 407610 74898 407846 75134
rect 438330 75218 438566 75454
rect 438330 74898 438566 75134
rect 469050 75218 469286 75454
rect 469050 74898 469286 75134
rect 499770 75218 500006 75454
rect 499770 74898 500006 75134
rect 530490 75218 530726 75454
rect 530490 74898 530726 75134
rect 561210 75218 561446 75454
rect 561210 74898 561446 75134
rect 567266 64658 567502 64894
rect 567586 64658 567822 64894
rect 567266 64338 567502 64574
rect 567586 64338 567822 64574
rect 23610 57218 23846 57454
rect 23610 56898 23846 57134
rect 54330 57218 54566 57454
rect 54330 56898 54566 57134
rect 85050 57218 85286 57454
rect 85050 56898 85286 57134
rect 115770 57218 116006 57454
rect 115770 56898 116006 57134
rect 146490 57218 146726 57454
rect 146490 56898 146726 57134
rect 177210 57218 177446 57454
rect 177210 56898 177446 57134
rect 207930 57218 208166 57454
rect 207930 56898 208166 57134
rect 238650 57218 238886 57454
rect 238650 56898 238886 57134
rect 269370 57218 269606 57454
rect 269370 56898 269606 57134
rect 300090 57218 300326 57454
rect 300090 56898 300326 57134
rect 330810 57218 331046 57454
rect 330810 56898 331046 57134
rect 361530 57218 361766 57454
rect 361530 56898 361766 57134
rect 392250 57218 392486 57454
rect 392250 56898 392486 57134
rect 422970 57218 423206 57454
rect 422970 56898 423206 57134
rect 453690 57218 453926 57454
rect 453690 56898 453926 57134
rect 484410 57218 484646 57454
rect 484410 56898 484646 57134
rect 515130 57218 515366 57454
rect 515130 56898 515366 57134
rect 545850 57218 546086 57454
rect 545850 56898 546086 57134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect 8250 39218 8486 39454
rect 8250 38898 8486 39134
rect 38970 39218 39206 39454
rect 38970 38898 39206 39134
rect 69690 39218 69926 39454
rect 69690 38898 69926 39134
rect 100410 39218 100646 39454
rect 100410 38898 100646 39134
rect 131130 39218 131366 39454
rect 131130 38898 131366 39134
rect 161850 39218 162086 39454
rect 161850 38898 162086 39134
rect 192570 39218 192806 39454
rect 192570 38898 192806 39134
rect 223290 39218 223526 39454
rect 223290 38898 223526 39134
rect 254010 39218 254246 39454
rect 254010 38898 254246 39134
rect 284730 39218 284966 39454
rect 284730 38898 284966 39134
rect 315450 39218 315686 39454
rect 315450 38898 315686 39134
rect 346170 39218 346406 39454
rect 346170 38898 346406 39134
rect 376890 39218 377126 39454
rect 376890 38898 377126 39134
rect 407610 39218 407846 39454
rect 407610 38898 407846 39134
rect 438330 39218 438566 39454
rect 438330 38898 438566 39134
rect 469050 39218 469286 39454
rect 469050 38898 469286 39134
rect 499770 39218 500006 39454
rect 499770 38898 500006 39134
rect 530490 39218 530726 39454
rect 530490 38898 530726 39134
rect 561210 39218 561446 39454
rect 561210 38898 561446 39134
rect 567266 28658 567502 28894
rect 567586 28658 567822 28894
rect 567266 28338 567502 28574
rect 567586 28338 567822 28574
rect 23610 21218 23846 21454
rect 23610 20898 23846 21134
rect 54330 21218 54566 21454
rect 54330 20898 54566 21134
rect 85050 21218 85286 21454
rect 85050 20898 85286 21134
rect 115770 21218 116006 21454
rect 115770 20898 116006 21134
rect 146490 21218 146726 21454
rect 146490 20898 146726 21134
rect 177210 21218 177446 21454
rect 177210 20898 177446 21134
rect 207930 21218 208166 21454
rect 207930 20898 208166 21134
rect 238650 21218 238886 21454
rect 238650 20898 238886 21134
rect 269370 21218 269606 21454
rect 269370 20898 269606 21134
rect 300090 21218 300326 21454
rect 300090 20898 300326 21134
rect 330810 21218 331046 21454
rect 330810 20898 331046 21134
rect 361530 21218 361766 21454
rect 361530 20898 361766 21134
rect 392250 21218 392486 21454
rect 392250 20898 392486 21134
rect 422970 21218 423206 21454
rect 422970 20898 423206 21134
rect 453690 21218 453926 21454
rect 453690 20898 453926 21134
rect 484410 21218 484646 21454
rect 484410 20898 484646 21134
rect 515130 21218 515366 21454
rect 515130 20898 515366 21134
rect 545850 21218 546086 21454
rect 545850 20898 546086 21134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect 8250 3218 8486 3454
rect 8250 2898 8486 3134
rect 38970 3218 39206 3454
rect 38970 2898 39206 3134
rect 69690 3218 69926 3454
rect 69690 2898 69926 3134
rect 100410 3218 100646 3454
rect 100410 2898 100646 3134
rect 131130 3218 131366 3454
rect 131130 2898 131366 3134
rect 161850 3218 162086 3454
rect 161850 2898 162086 3134
rect 192570 3218 192806 3454
rect 192570 2898 192806 3134
rect 223290 3218 223526 3454
rect 223290 2898 223526 3134
rect 254010 3218 254246 3454
rect 254010 2898 254246 3134
rect 284730 3218 284966 3454
rect 284730 2898 284966 3134
rect 315450 3218 315686 3454
rect 315450 2898 315686 3134
rect 346170 3218 346406 3454
rect 346170 2898 346406 3134
rect 376890 3218 377126 3454
rect 376890 2898 377126 3134
rect 407610 3218 407846 3454
rect 407610 2898 407846 3134
rect 438330 3218 438566 3454
rect 438330 2898 438566 3134
rect 469050 3218 469286 3454
rect 469050 2898 469286 3134
rect 499770 3218 500006 3454
rect 499770 2898 500006 3134
rect 530490 3218 530726 3454
rect 530490 2898 530726 3134
rect 561210 3218 561446 3454
rect 561210 2898 561446 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 5546 -2502 5782 -2266
rect 5866 -2502 6102 -2266
rect 5546 -2822 5782 -2586
rect 5866 -2822 6102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 9266 -4422 9502 -4186
rect 9586 -4422 9822 -4186
rect 9266 -4742 9502 -4506
rect 9586 -4742 9822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 23546 -3462 23782 -3226
rect 23866 -3462 24102 -3226
rect 23546 -3782 23782 -3546
rect 23866 -3782 24102 -3546
rect 27266 -5382 27502 -5146
rect 27586 -5382 27822 -5146
rect 27266 -5702 27502 -5466
rect 27586 -5702 27822 -5466
rect 12986 -6342 13222 -6106
rect 13306 -6342 13542 -6106
rect 12986 -6662 13222 -6426
rect 13306 -6662 13542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 41546 -2502 41782 -2266
rect 41866 -2502 42102 -2266
rect 41546 -2822 41782 -2586
rect 41866 -2822 42102 -2586
rect 45266 -4422 45502 -4186
rect 45586 -4422 45822 -4186
rect 45266 -4742 45502 -4506
rect 45586 -4742 45822 -4506
rect 30986 -7302 31222 -7066
rect 31306 -7302 31542 -7066
rect 30986 -7622 31222 -7386
rect 31306 -7622 31542 -7386
rect 59546 -3462 59782 -3226
rect 59866 -3462 60102 -3226
rect 59546 -3782 59782 -3546
rect 59866 -3782 60102 -3546
rect 63266 -5382 63502 -5146
rect 63586 -5382 63822 -5146
rect 63266 -5702 63502 -5466
rect 63586 -5702 63822 -5466
rect 48986 -6342 49222 -6106
rect 49306 -6342 49542 -6106
rect 48986 -6662 49222 -6426
rect 49306 -6662 49542 -6426
rect 77546 -2502 77782 -2266
rect 77866 -2502 78102 -2266
rect 77546 -2822 77782 -2586
rect 77866 -2822 78102 -2586
rect 81266 -4422 81502 -4186
rect 81586 -4422 81822 -4186
rect 81266 -4742 81502 -4506
rect 81586 -4742 81822 -4506
rect 66986 -7302 67222 -7066
rect 67306 -7302 67542 -7066
rect 66986 -7622 67222 -7386
rect 67306 -7622 67542 -7386
rect 95546 -3462 95782 -3226
rect 95866 -3462 96102 -3226
rect 95546 -3782 95782 -3546
rect 95866 -3782 96102 -3546
rect 99266 -5382 99502 -5146
rect 99586 -5382 99822 -5146
rect 99266 -5702 99502 -5466
rect 99586 -5702 99822 -5466
rect 84986 -6342 85222 -6106
rect 85306 -6342 85542 -6106
rect 84986 -6662 85222 -6426
rect 85306 -6662 85542 -6426
rect 113546 -2502 113782 -2266
rect 113866 -2502 114102 -2266
rect 113546 -2822 113782 -2586
rect 113866 -2822 114102 -2586
rect 117266 -4422 117502 -4186
rect 117586 -4422 117822 -4186
rect 117266 -4742 117502 -4506
rect 117586 -4742 117822 -4506
rect 102986 -7302 103222 -7066
rect 103306 -7302 103542 -7066
rect 102986 -7622 103222 -7386
rect 103306 -7622 103542 -7386
rect 131546 -3462 131782 -3226
rect 131866 -3462 132102 -3226
rect 131546 -3782 131782 -3546
rect 131866 -3782 132102 -3546
rect 135266 -5382 135502 -5146
rect 135586 -5382 135822 -5146
rect 135266 -5702 135502 -5466
rect 135586 -5702 135822 -5466
rect 120986 -6342 121222 -6106
rect 121306 -6342 121542 -6106
rect 120986 -6662 121222 -6426
rect 121306 -6662 121542 -6426
rect 149546 -2502 149782 -2266
rect 149866 -2502 150102 -2266
rect 149546 -2822 149782 -2586
rect 149866 -2822 150102 -2586
rect 153266 -4422 153502 -4186
rect 153586 -4422 153822 -4186
rect 153266 -4742 153502 -4506
rect 153586 -4742 153822 -4506
rect 138986 -7302 139222 -7066
rect 139306 -7302 139542 -7066
rect 138986 -7622 139222 -7386
rect 139306 -7622 139542 -7386
rect 167546 -3462 167782 -3226
rect 167866 -3462 168102 -3226
rect 167546 -3782 167782 -3546
rect 167866 -3782 168102 -3546
rect 171266 -5382 171502 -5146
rect 171586 -5382 171822 -5146
rect 171266 -5702 171502 -5466
rect 171586 -5702 171822 -5466
rect 156986 -6342 157222 -6106
rect 157306 -6342 157542 -6106
rect 156986 -6662 157222 -6426
rect 157306 -6662 157542 -6426
rect 185546 -2502 185782 -2266
rect 185866 -2502 186102 -2266
rect 185546 -2822 185782 -2586
rect 185866 -2822 186102 -2586
rect 189266 -4422 189502 -4186
rect 189586 -4422 189822 -4186
rect 189266 -4742 189502 -4506
rect 189586 -4742 189822 -4506
rect 174986 -7302 175222 -7066
rect 175306 -7302 175542 -7066
rect 174986 -7622 175222 -7386
rect 175306 -7622 175542 -7386
rect 203546 -3462 203782 -3226
rect 203866 -3462 204102 -3226
rect 203546 -3782 203782 -3546
rect 203866 -3782 204102 -3546
rect 207266 -5382 207502 -5146
rect 207586 -5382 207822 -5146
rect 207266 -5702 207502 -5466
rect 207586 -5702 207822 -5466
rect 192986 -6342 193222 -6106
rect 193306 -6342 193542 -6106
rect 192986 -6662 193222 -6426
rect 193306 -6662 193542 -6426
rect 221546 -2502 221782 -2266
rect 221866 -2502 222102 -2266
rect 221546 -2822 221782 -2586
rect 221866 -2822 222102 -2586
rect 225266 -4422 225502 -4186
rect 225586 -4422 225822 -4186
rect 225266 -4742 225502 -4506
rect 225586 -4742 225822 -4506
rect 210986 -7302 211222 -7066
rect 211306 -7302 211542 -7066
rect 210986 -7622 211222 -7386
rect 211306 -7622 211542 -7386
rect 239546 -3462 239782 -3226
rect 239866 -3462 240102 -3226
rect 239546 -3782 239782 -3546
rect 239866 -3782 240102 -3546
rect 243266 -5382 243502 -5146
rect 243586 -5382 243822 -5146
rect 243266 -5702 243502 -5466
rect 243586 -5702 243822 -5466
rect 228986 -6342 229222 -6106
rect 229306 -6342 229542 -6106
rect 228986 -6662 229222 -6426
rect 229306 -6662 229542 -6426
rect 257546 -2502 257782 -2266
rect 257866 -2502 258102 -2266
rect 257546 -2822 257782 -2586
rect 257866 -2822 258102 -2586
rect 261266 -4422 261502 -4186
rect 261586 -4422 261822 -4186
rect 261266 -4742 261502 -4506
rect 261586 -4742 261822 -4506
rect 246986 -7302 247222 -7066
rect 247306 -7302 247542 -7066
rect 246986 -7622 247222 -7386
rect 247306 -7622 247542 -7386
rect 275546 -3462 275782 -3226
rect 275866 -3462 276102 -3226
rect 275546 -3782 275782 -3546
rect 275866 -3782 276102 -3546
rect 279266 -5382 279502 -5146
rect 279586 -5382 279822 -5146
rect 279266 -5702 279502 -5466
rect 279586 -5702 279822 -5466
rect 264986 -6342 265222 -6106
rect 265306 -6342 265542 -6106
rect 264986 -6662 265222 -6426
rect 265306 -6662 265542 -6426
rect 293546 -2502 293782 -2266
rect 293866 -2502 294102 -2266
rect 293546 -2822 293782 -2586
rect 293866 -2822 294102 -2586
rect 297266 -4422 297502 -4186
rect 297586 -4422 297822 -4186
rect 297266 -4742 297502 -4506
rect 297586 -4742 297822 -4506
rect 282986 -7302 283222 -7066
rect 283306 -7302 283542 -7066
rect 282986 -7622 283222 -7386
rect 283306 -7622 283542 -7386
rect 311546 -3462 311782 -3226
rect 311866 -3462 312102 -3226
rect 311546 -3782 311782 -3546
rect 311866 -3782 312102 -3546
rect 315266 -5382 315502 -5146
rect 315586 -5382 315822 -5146
rect 315266 -5702 315502 -5466
rect 315586 -5702 315822 -5466
rect 300986 -6342 301222 -6106
rect 301306 -6342 301542 -6106
rect 300986 -6662 301222 -6426
rect 301306 -6662 301542 -6426
rect 329546 -2502 329782 -2266
rect 329866 -2502 330102 -2266
rect 329546 -2822 329782 -2586
rect 329866 -2822 330102 -2586
rect 333266 -4422 333502 -4186
rect 333586 -4422 333822 -4186
rect 333266 -4742 333502 -4506
rect 333586 -4742 333822 -4506
rect 318986 -7302 319222 -7066
rect 319306 -7302 319542 -7066
rect 318986 -7622 319222 -7386
rect 319306 -7622 319542 -7386
rect 347546 -3462 347782 -3226
rect 347866 -3462 348102 -3226
rect 347546 -3782 347782 -3546
rect 347866 -3782 348102 -3546
rect 351266 -5382 351502 -5146
rect 351586 -5382 351822 -5146
rect 351266 -5702 351502 -5466
rect 351586 -5702 351822 -5466
rect 336986 -6342 337222 -6106
rect 337306 -6342 337542 -6106
rect 336986 -6662 337222 -6426
rect 337306 -6662 337542 -6426
rect 365546 -2502 365782 -2266
rect 365866 -2502 366102 -2266
rect 365546 -2822 365782 -2586
rect 365866 -2822 366102 -2586
rect 369266 -4422 369502 -4186
rect 369586 -4422 369822 -4186
rect 369266 -4742 369502 -4506
rect 369586 -4742 369822 -4506
rect 354986 -7302 355222 -7066
rect 355306 -7302 355542 -7066
rect 354986 -7622 355222 -7386
rect 355306 -7622 355542 -7386
rect 383546 -3462 383782 -3226
rect 383866 -3462 384102 -3226
rect 383546 -3782 383782 -3546
rect 383866 -3782 384102 -3546
rect 387266 -5382 387502 -5146
rect 387586 -5382 387822 -5146
rect 387266 -5702 387502 -5466
rect 387586 -5702 387822 -5466
rect 372986 -6342 373222 -6106
rect 373306 -6342 373542 -6106
rect 372986 -6662 373222 -6426
rect 373306 -6662 373542 -6426
rect 401546 -2502 401782 -2266
rect 401866 -2502 402102 -2266
rect 401546 -2822 401782 -2586
rect 401866 -2822 402102 -2586
rect 405266 -4422 405502 -4186
rect 405586 -4422 405822 -4186
rect 405266 -4742 405502 -4506
rect 405586 -4742 405822 -4506
rect 390986 -7302 391222 -7066
rect 391306 -7302 391542 -7066
rect 390986 -7622 391222 -7386
rect 391306 -7622 391542 -7386
rect 419546 -3462 419782 -3226
rect 419866 -3462 420102 -3226
rect 419546 -3782 419782 -3546
rect 419866 -3782 420102 -3546
rect 423266 -5382 423502 -5146
rect 423586 -5382 423822 -5146
rect 423266 -5702 423502 -5466
rect 423586 -5702 423822 -5466
rect 408986 -6342 409222 -6106
rect 409306 -6342 409542 -6106
rect 408986 -6662 409222 -6426
rect 409306 -6662 409542 -6426
rect 437546 -2502 437782 -2266
rect 437866 -2502 438102 -2266
rect 437546 -2822 437782 -2586
rect 437866 -2822 438102 -2586
rect 441266 -4422 441502 -4186
rect 441586 -4422 441822 -4186
rect 441266 -4742 441502 -4506
rect 441586 -4742 441822 -4506
rect 426986 -7302 427222 -7066
rect 427306 -7302 427542 -7066
rect 426986 -7622 427222 -7386
rect 427306 -7622 427542 -7386
rect 455546 -3462 455782 -3226
rect 455866 -3462 456102 -3226
rect 455546 -3782 455782 -3546
rect 455866 -3782 456102 -3546
rect 459266 -5382 459502 -5146
rect 459586 -5382 459822 -5146
rect 459266 -5702 459502 -5466
rect 459586 -5702 459822 -5466
rect 444986 -6342 445222 -6106
rect 445306 -6342 445542 -6106
rect 444986 -6662 445222 -6426
rect 445306 -6662 445542 -6426
rect 473546 -2502 473782 -2266
rect 473866 -2502 474102 -2266
rect 473546 -2822 473782 -2586
rect 473866 -2822 474102 -2586
rect 477266 -4422 477502 -4186
rect 477586 -4422 477822 -4186
rect 477266 -4742 477502 -4506
rect 477586 -4742 477822 -4506
rect 462986 -7302 463222 -7066
rect 463306 -7302 463542 -7066
rect 462986 -7622 463222 -7386
rect 463306 -7622 463542 -7386
rect 491546 -3462 491782 -3226
rect 491866 -3462 492102 -3226
rect 491546 -3782 491782 -3546
rect 491866 -3782 492102 -3546
rect 495266 -5382 495502 -5146
rect 495586 -5382 495822 -5146
rect 495266 -5702 495502 -5466
rect 495586 -5702 495822 -5466
rect 480986 -6342 481222 -6106
rect 481306 -6342 481542 -6106
rect 480986 -6662 481222 -6426
rect 481306 -6662 481542 -6426
rect 509546 -2502 509782 -2266
rect 509866 -2502 510102 -2266
rect 509546 -2822 509782 -2586
rect 509866 -2822 510102 -2586
rect 513266 -4422 513502 -4186
rect 513586 -4422 513822 -4186
rect 513266 -4742 513502 -4506
rect 513586 -4742 513822 -4506
rect 498986 -7302 499222 -7066
rect 499306 -7302 499542 -7066
rect 498986 -7622 499222 -7386
rect 499306 -7622 499542 -7386
rect 527546 -3462 527782 -3226
rect 527866 -3462 528102 -3226
rect 527546 -3782 527782 -3546
rect 527866 -3782 528102 -3546
rect 531266 -5382 531502 -5146
rect 531586 -5382 531822 -5146
rect 531266 -5702 531502 -5466
rect 531586 -5702 531822 -5466
rect 516986 -6342 517222 -6106
rect 517306 -6342 517542 -6106
rect 516986 -6662 517222 -6426
rect 517306 -6662 517542 -6426
rect 545546 -2502 545782 -2266
rect 545866 -2502 546102 -2266
rect 545546 -2822 545782 -2586
rect 545866 -2822 546102 -2586
rect 549266 -4422 549502 -4186
rect 549586 -4422 549822 -4186
rect 549266 -4742 549502 -4506
rect 549586 -4742 549822 -4506
rect 534986 -7302 535222 -7066
rect 535306 -7302 535542 -7066
rect 534986 -7622 535222 -7386
rect 535306 -7622 535542 -7386
rect 563546 -3462 563782 -3226
rect 563866 -3462 564102 -3226
rect 563546 -3782 563782 -3546
rect 563866 -3782 564102 -3546
rect 567266 -5382 567502 -5146
rect 567586 -5382 567822 -5146
rect 567266 -5702 567502 -5466
rect 567586 -5702 567822 -5466
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 581546 706522 581782 706758
rect 581866 706522 582102 706758
rect 581546 706202 581782 706438
rect 581866 706202 582102 706438
rect 570986 680378 571222 680614
rect 571306 680378 571542 680614
rect 570986 680058 571222 680294
rect 571306 680058 571542 680294
rect 570986 644378 571222 644614
rect 571306 644378 571542 644614
rect 570986 644058 571222 644294
rect 571306 644058 571542 644294
rect 570986 608378 571222 608614
rect 571306 608378 571542 608614
rect 570986 608058 571222 608294
rect 571306 608058 571542 608294
rect 570986 572378 571222 572614
rect 571306 572378 571542 572614
rect 570986 572058 571222 572294
rect 571306 572058 571542 572294
rect 570986 536378 571222 536614
rect 571306 536378 571542 536614
rect 570986 536058 571222 536294
rect 571306 536058 571542 536294
rect 570986 500378 571222 500614
rect 571306 500378 571542 500614
rect 570986 500058 571222 500294
rect 571306 500058 571542 500294
rect 570986 464378 571222 464614
rect 571306 464378 571542 464614
rect 570986 464058 571222 464294
rect 571306 464058 571542 464294
rect 570986 428378 571222 428614
rect 571306 428378 571542 428614
rect 570986 428058 571222 428294
rect 571306 428058 571542 428294
rect 570986 392378 571222 392614
rect 571306 392378 571542 392614
rect 570986 392058 571222 392294
rect 571306 392058 571542 392294
rect 570986 356378 571222 356614
rect 571306 356378 571542 356614
rect 570986 356058 571222 356294
rect 571306 356058 571542 356294
rect 570986 320378 571222 320614
rect 571306 320378 571542 320614
rect 570986 320058 571222 320294
rect 571306 320058 571542 320294
rect 570986 284378 571222 284614
rect 571306 284378 571542 284614
rect 570986 284058 571222 284294
rect 571306 284058 571542 284294
rect 570986 248378 571222 248614
rect 571306 248378 571542 248614
rect 570986 248058 571222 248294
rect 571306 248058 571542 248294
rect 570986 212378 571222 212614
rect 571306 212378 571542 212614
rect 570986 212058 571222 212294
rect 571306 212058 571542 212294
rect 570986 176378 571222 176614
rect 571306 176378 571542 176614
rect 570986 176058 571222 176294
rect 571306 176058 571542 176294
rect 570986 140378 571222 140614
rect 571306 140378 571542 140614
rect 570986 140058 571222 140294
rect 571306 140058 571542 140294
rect 570986 104378 571222 104614
rect 571306 104378 571542 104614
rect 570986 104058 571222 104294
rect 571306 104058 571542 104294
rect 570986 68378 571222 68614
rect 571306 68378 571542 68614
rect 570986 68058 571222 68294
rect 571306 68058 571542 68294
rect 570986 32378 571222 32614
rect 571306 32378 571542 32614
rect 570986 32058 571222 32294
rect 571306 32058 571542 32294
rect 552986 -6342 553222 -6106
rect 553306 -6342 553542 -6106
rect 552986 -6662 553222 -6426
rect 553306 -6662 553542 -6426
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 690938 587498 691174
rect 587582 690938 587818 691174
rect 587262 690618 587498 690854
rect 587582 690618 587818 690854
rect 587262 654938 587498 655174
rect 587582 654938 587818 655174
rect 587262 654618 587498 654854
rect 587582 654618 587818 654854
rect 587262 618938 587498 619174
rect 587582 618938 587818 619174
rect 587262 618618 587498 618854
rect 587582 618618 587818 618854
rect 587262 582938 587498 583174
rect 587582 582938 587818 583174
rect 587262 582618 587498 582854
rect 587582 582618 587818 582854
rect 587262 546938 587498 547174
rect 587582 546938 587818 547174
rect 587262 546618 587498 546854
rect 587582 546618 587818 546854
rect 587262 510938 587498 511174
rect 587582 510938 587818 511174
rect 587262 510618 587498 510854
rect 587582 510618 587818 510854
rect 587262 474938 587498 475174
rect 587582 474938 587818 475174
rect 587262 474618 587498 474854
rect 587582 474618 587818 474854
rect 587262 438938 587498 439174
rect 587582 438938 587818 439174
rect 587262 438618 587498 438854
rect 587582 438618 587818 438854
rect 587262 402938 587498 403174
rect 587582 402938 587818 403174
rect 587262 402618 587498 402854
rect 587582 402618 587818 402854
rect 587262 366938 587498 367174
rect 587582 366938 587818 367174
rect 587262 366618 587498 366854
rect 587582 366618 587818 366854
rect 587262 330938 587498 331174
rect 587582 330938 587818 331174
rect 587262 330618 587498 330854
rect 587582 330618 587818 330854
rect 587262 294938 587498 295174
rect 587582 294938 587818 295174
rect 587262 294618 587498 294854
rect 587582 294618 587818 294854
rect 587262 258938 587498 259174
rect 587582 258938 587818 259174
rect 587262 258618 587498 258854
rect 587582 258618 587818 258854
rect 587262 222938 587498 223174
rect 587582 222938 587818 223174
rect 587262 222618 587498 222854
rect 587582 222618 587818 222854
rect 587262 186938 587498 187174
rect 587582 186938 587818 187174
rect 587262 186618 587498 186854
rect 587582 186618 587818 186854
rect 587262 150938 587498 151174
rect 587582 150938 587818 151174
rect 587262 150618 587498 150854
rect 587582 150618 587818 150854
rect 587262 114938 587498 115174
rect 587582 114938 587818 115174
rect 587262 114618 587498 114854
rect 587582 114618 587818 114854
rect 587262 78938 587498 79174
rect 587582 78938 587818 79174
rect 587262 78618 587498 78854
rect 587582 78618 587818 78854
rect 587262 42938 587498 43174
rect 587582 42938 587818 43174
rect 587262 42618 587498 42854
rect 587582 42618 587818 42854
rect 587262 6938 587498 7174
rect 587582 6938 587818 7174
rect 587262 6618 587498 6854
rect 587582 6618 587818 6854
rect 581546 -2502 581782 -2266
rect 581866 -2502 582102 -2266
rect 581546 -2822 581782 -2586
rect 581866 -2822 582102 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 672938 588458 673174
rect 588542 672938 588778 673174
rect 588222 672618 588458 672854
rect 588542 672618 588778 672854
rect 588222 636938 588458 637174
rect 588542 636938 588778 637174
rect 588222 636618 588458 636854
rect 588542 636618 588778 636854
rect 588222 600938 588458 601174
rect 588542 600938 588778 601174
rect 588222 600618 588458 600854
rect 588542 600618 588778 600854
rect 588222 564938 588458 565174
rect 588542 564938 588778 565174
rect 588222 564618 588458 564854
rect 588542 564618 588778 564854
rect 588222 528938 588458 529174
rect 588542 528938 588778 529174
rect 588222 528618 588458 528854
rect 588542 528618 588778 528854
rect 588222 492938 588458 493174
rect 588542 492938 588778 493174
rect 588222 492618 588458 492854
rect 588542 492618 588778 492854
rect 588222 456938 588458 457174
rect 588542 456938 588778 457174
rect 588222 456618 588458 456854
rect 588542 456618 588778 456854
rect 588222 420938 588458 421174
rect 588542 420938 588778 421174
rect 588222 420618 588458 420854
rect 588542 420618 588778 420854
rect 588222 384938 588458 385174
rect 588542 384938 588778 385174
rect 588222 384618 588458 384854
rect 588542 384618 588778 384854
rect 588222 348938 588458 349174
rect 588542 348938 588778 349174
rect 588222 348618 588458 348854
rect 588542 348618 588778 348854
rect 588222 312938 588458 313174
rect 588542 312938 588778 313174
rect 588222 312618 588458 312854
rect 588542 312618 588778 312854
rect 588222 276938 588458 277174
rect 588542 276938 588778 277174
rect 588222 276618 588458 276854
rect 588542 276618 588778 276854
rect 588222 240938 588458 241174
rect 588542 240938 588778 241174
rect 588222 240618 588458 240854
rect 588542 240618 588778 240854
rect 588222 204938 588458 205174
rect 588542 204938 588778 205174
rect 588222 204618 588458 204854
rect 588542 204618 588778 204854
rect 588222 168938 588458 169174
rect 588542 168938 588778 169174
rect 588222 168618 588458 168854
rect 588542 168618 588778 168854
rect 588222 132938 588458 133174
rect 588542 132938 588778 133174
rect 588222 132618 588458 132854
rect 588542 132618 588778 132854
rect 588222 96938 588458 97174
rect 588542 96938 588778 97174
rect 588222 96618 588458 96854
rect 588542 96618 588778 96854
rect 588222 60938 588458 61174
rect 588542 60938 588778 61174
rect 588222 60618 588458 60854
rect 588542 60618 588778 60854
rect 588222 24938 588458 25174
rect 588542 24938 588778 25174
rect 588222 24618 588458 24854
rect 588542 24618 588778 24854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 694658 589418 694894
rect 589502 694658 589738 694894
rect 589182 694338 589418 694574
rect 589502 694338 589738 694574
rect 589182 658658 589418 658894
rect 589502 658658 589738 658894
rect 589182 658338 589418 658574
rect 589502 658338 589738 658574
rect 589182 622658 589418 622894
rect 589502 622658 589738 622894
rect 589182 622338 589418 622574
rect 589502 622338 589738 622574
rect 589182 586658 589418 586894
rect 589502 586658 589738 586894
rect 589182 586338 589418 586574
rect 589502 586338 589738 586574
rect 589182 550658 589418 550894
rect 589502 550658 589738 550894
rect 589182 550338 589418 550574
rect 589502 550338 589738 550574
rect 589182 514658 589418 514894
rect 589502 514658 589738 514894
rect 589182 514338 589418 514574
rect 589502 514338 589738 514574
rect 589182 478658 589418 478894
rect 589502 478658 589738 478894
rect 589182 478338 589418 478574
rect 589502 478338 589738 478574
rect 589182 442658 589418 442894
rect 589502 442658 589738 442894
rect 589182 442338 589418 442574
rect 589502 442338 589738 442574
rect 589182 406658 589418 406894
rect 589502 406658 589738 406894
rect 589182 406338 589418 406574
rect 589502 406338 589738 406574
rect 589182 370658 589418 370894
rect 589502 370658 589738 370894
rect 589182 370338 589418 370574
rect 589502 370338 589738 370574
rect 589182 334658 589418 334894
rect 589502 334658 589738 334894
rect 589182 334338 589418 334574
rect 589502 334338 589738 334574
rect 589182 298658 589418 298894
rect 589502 298658 589738 298894
rect 589182 298338 589418 298574
rect 589502 298338 589738 298574
rect 589182 262658 589418 262894
rect 589502 262658 589738 262894
rect 589182 262338 589418 262574
rect 589502 262338 589738 262574
rect 589182 226658 589418 226894
rect 589502 226658 589738 226894
rect 589182 226338 589418 226574
rect 589502 226338 589738 226574
rect 589182 190658 589418 190894
rect 589502 190658 589738 190894
rect 589182 190338 589418 190574
rect 589502 190338 589738 190574
rect 589182 154658 589418 154894
rect 589502 154658 589738 154894
rect 589182 154338 589418 154574
rect 589502 154338 589738 154574
rect 589182 118658 589418 118894
rect 589502 118658 589738 118894
rect 589182 118338 589418 118574
rect 589502 118338 589738 118574
rect 589182 82658 589418 82894
rect 589502 82658 589738 82894
rect 589182 82338 589418 82574
rect 589502 82338 589738 82574
rect 589182 46658 589418 46894
rect 589502 46658 589738 46894
rect 589182 46338 589418 46574
rect 589502 46338 589738 46574
rect 589182 10658 589418 10894
rect 589502 10658 589738 10894
rect 589182 10338 589418 10574
rect 589502 10338 589738 10574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 676658 590378 676894
rect 590462 676658 590698 676894
rect 590142 676338 590378 676574
rect 590462 676338 590698 676574
rect 590142 640658 590378 640894
rect 590462 640658 590698 640894
rect 590142 640338 590378 640574
rect 590462 640338 590698 640574
rect 590142 604658 590378 604894
rect 590462 604658 590698 604894
rect 590142 604338 590378 604574
rect 590462 604338 590698 604574
rect 590142 568658 590378 568894
rect 590462 568658 590698 568894
rect 590142 568338 590378 568574
rect 590462 568338 590698 568574
rect 590142 532658 590378 532894
rect 590462 532658 590698 532894
rect 590142 532338 590378 532574
rect 590462 532338 590698 532574
rect 590142 496658 590378 496894
rect 590462 496658 590698 496894
rect 590142 496338 590378 496574
rect 590462 496338 590698 496574
rect 590142 460658 590378 460894
rect 590462 460658 590698 460894
rect 590142 460338 590378 460574
rect 590462 460338 590698 460574
rect 590142 424658 590378 424894
rect 590462 424658 590698 424894
rect 590142 424338 590378 424574
rect 590462 424338 590698 424574
rect 590142 388658 590378 388894
rect 590462 388658 590698 388894
rect 590142 388338 590378 388574
rect 590462 388338 590698 388574
rect 590142 352658 590378 352894
rect 590462 352658 590698 352894
rect 590142 352338 590378 352574
rect 590462 352338 590698 352574
rect 590142 316658 590378 316894
rect 590462 316658 590698 316894
rect 590142 316338 590378 316574
rect 590462 316338 590698 316574
rect 590142 280658 590378 280894
rect 590462 280658 590698 280894
rect 590142 280338 590378 280574
rect 590462 280338 590698 280574
rect 590142 244658 590378 244894
rect 590462 244658 590698 244894
rect 590142 244338 590378 244574
rect 590462 244338 590698 244574
rect 590142 208658 590378 208894
rect 590462 208658 590698 208894
rect 590142 208338 590378 208574
rect 590462 208338 590698 208574
rect 590142 172658 590378 172894
rect 590462 172658 590698 172894
rect 590142 172338 590378 172574
rect 590462 172338 590698 172574
rect 590142 136658 590378 136894
rect 590462 136658 590698 136894
rect 590142 136338 590378 136574
rect 590462 136338 590698 136574
rect 590142 100658 590378 100894
rect 590462 100658 590698 100894
rect 590142 100338 590378 100574
rect 590462 100338 590698 100574
rect 590142 64658 590378 64894
rect 590462 64658 590698 64894
rect 590142 64338 590378 64574
rect 590462 64338 590698 64574
rect 590142 28658 590378 28894
rect 590462 28658 590698 28894
rect 590142 28338 590378 28574
rect 590462 28338 590698 28574
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 698378 591338 698614
rect 591422 698378 591658 698614
rect 591102 698058 591338 698294
rect 591422 698058 591658 698294
rect 591102 662378 591338 662614
rect 591422 662378 591658 662614
rect 591102 662058 591338 662294
rect 591422 662058 591658 662294
rect 591102 626378 591338 626614
rect 591422 626378 591658 626614
rect 591102 626058 591338 626294
rect 591422 626058 591658 626294
rect 591102 590378 591338 590614
rect 591422 590378 591658 590614
rect 591102 590058 591338 590294
rect 591422 590058 591658 590294
rect 591102 554378 591338 554614
rect 591422 554378 591658 554614
rect 591102 554058 591338 554294
rect 591422 554058 591658 554294
rect 591102 518378 591338 518614
rect 591422 518378 591658 518614
rect 591102 518058 591338 518294
rect 591422 518058 591658 518294
rect 591102 482378 591338 482614
rect 591422 482378 591658 482614
rect 591102 482058 591338 482294
rect 591422 482058 591658 482294
rect 591102 446378 591338 446614
rect 591422 446378 591658 446614
rect 591102 446058 591338 446294
rect 591422 446058 591658 446294
rect 591102 410378 591338 410614
rect 591422 410378 591658 410614
rect 591102 410058 591338 410294
rect 591422 410058 591658 410294
rect 591102 374378 591338 374614
rect 591422 374378 591658 374614
rect 591102 374058 591338 374294
rect 591422 374058 591658 374294
rect 591102 338378 591338 338614
rect 591422 338378 591658 338614
rect 591102 338058 591338 338294
rect 591422 338058 591658 338294
rect 591102 302378 591338 302614
rect 591422 302378 591658 302614
rect 591102 302058 591338 302294
rect 591422 302058 591658 302294
rect 591102 266378 591338 266614
rect 591422 266378 591658 266614
rect 591102 266058 591338 266294
rect 591422 266058 591658 266294
rect 591102 230378 591338 230614
rect 591422 230378 591658 230614
rect 591102 230058 591338 230294
rect 591422 230058 591658 230294
rect 591102 194378 591338 194614
rect 591422 194378 591658 194614
rect 591102 194058 591338 194294
rect 591422 194058 591658 194294
rect 591102 158378 591338 158614
rect 591422 158378 591658 158614
rect 591102 158058 591338 158294
rect 591422 158058 591658 158294
rect 591102 122378 591338 122614
rect 591422 122378 591658 122614
rect 591102 122058 591338 122294
rect 591422 122058 591658 122294
rect 591102 86378 591338 86614
rect 591422 86378 591658 86614
rect 591102 86058 591338 86294
rect 591422 86058 591658 86294
rect 591102 50378 591338 50614
rect 591422 50378 591658 50614
rect 591102 50058 591338 50294
rect 591422 50058 591658 50294
rect 591102 14378 591338 14614
rect 591422 14378 591658 14614
rect 591102 14058 591338 14294
rect 591422 14058 591658 14294
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 680378 592298 680614
rect 592382 680378 592618 680614
rect 592062 680058 592298 680294
rect 592382 680058 592618 680294
rect 592062 644378 592298 644614
rect 592382 644378 592618 644614
rect 592062 644058 592298 644294
rect 592382 644058 592618 644294
rect 592062 608378 592298 608614
rect 592382 608378 592618 608614
rect 592062 608058 592298 608294
rect 592382 608058 592618 608294
rect 592062 572378 592298 572614
rect 592382 572378 592618 572614
rect 592062 572058 592298 572294
rect 592382 572058 592618 572294
rect 592062 536378 592298 536614
rect 592382 536378 592618 536614
rect 592062 536058 592298 536294
rect 592382 536058 592618 536294
rect 592062 500378 592298 500614
rect 592382 500378 592618 500614
rect 592062 500058 592298 500294
rect 592382 500058 592618 500294
rect 592062 464378 592298 464614
rect 592382 464378 592618 464614
rect 592062 464058 592298 464294
rect 592382 464058 592618 464294
rect 592062 428378 592298 428614
rect 592382 428378 592618 428614
rect 592062 428058 592298 428294
rect 592382 428058 592618 428294
rect 592062 392378 592298 392614
rect 592382 392378 592618 392614
rect 592062 392058 592298 392294
rect 592382 392058 592618 392294
rect 592062 356378 592298 356614
rect 592382 356378 592618 356614
rect 592062 356058 592298 356294
rect 592382 356058 592618 356294
rect 592062 320378 592298 320614
rect 592382 320378 592618 320614
rect 592062 320058 592298 320294
rect 592382 320058 592618 320294
rect 592062 284378 592298 284614
rect 592382 284378 592618 284614
rect 592062 284058 592298 284294
rect 592382 284058 592618 284294
rect 592062 248378 592298 248614
rect 592382 248378 592618 248614
rect 592062 248058 592298 248294
rect 592382 248058 592618 248294
rect 592062 212378 592298 212614
rect 592382 212378 592618 212614
rect 592062 212058 592298 212294
rect 592382 212058 592618 212294
rect 592062 176378 592298 176614
rect 592382 176378 592618 176614
rect 592062 176058 592298 176294
rect 592382 176058 592618 176294
rect 592062 140378 592298 140614
rect 592382 140378 592618 140614
rect 592062 140058 592298 140294
rect 592382 140058 592618 140294
rect 592062 104378 592298 104614
rect 592382 104378 592618 104614
rect 592062 104058 592298 104294
rect 592382 104058 592618 104294
rect 592062 68378 592298 68614
rect 592382 68378 592618 68614
rect 592062 68058 592298 68294
rect 592382 68058 592618 68294
rect 592062 32378 592298 32614
rect 592382 32378 592618 32614
rect 592062 32058 592298 32294
rect 592382 32058 592618 32294
rect 570986 -7302 571222 -7066
rect 571306 -7302 571542 -7066
rect 570986 -7622 571222 -7386
rect 571306 -7622 571542 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 592650 698294
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 590730 694894
rect -6806 694574 590730 694658
rect -6806 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 590730 694574
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 588810 691174
rect -4886 690854 588810 690938
rect -4886 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 588810 690854
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 8250 687454
rect 8486 687218 38970 687454
rect 39206 687218 69690 687454
rect 69926 687218 100410 687454
rect 100646 687218 131130 687454
rect 131366 687218 161850 687454
rect 162086 687218 192570 687454
rect 192806 687218 223290 687454
rect 223526 687218 254010 687454
rect 254246 687218 284730 687454
rect 284966 687218 315450 687454
rect 315686 687218 346170 687454
rect 346406 687218 376890 687454
rect 377126 687218 407610 687454
rect 407846 687218 438330 687454
rect 438566 687218 469050 687454
rect 469286 687218 499770 687454
rect 500006 687218 530490 687454
rect 530726 687218 561210 687454
rect 561446 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 8250 687134
rect 8486 686898 38970 687134
rect 39206 686898 69690 687134
rect 69926 686898 100410 687134
rect 100646 686898 131130 687134
rect 131366 686898 161850 687134
rect 162086 686898 192570 687134
rect 192806 686898 223290 687134
rect 223526 686898 254010 687134
rect 254246 686898 284730 687134
rect 284966 686898 315450 687134
rect 315686 686898 346170 687134
rect 346406 686898 376890 687134
rect 377126 686898 407610 687134
rect 407846 686898 438330 687134
rect 438566 686898 469050 687134
rect 469286 686898 499770 687134
rect 500006 686898 530490 687134
rect 530726 686898 561210 687134
rect 561446 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect -8726 680294 592650 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect -6806 676574 590730 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect -4886 672854 588810 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 23610 669454
rect 23846 669218 54330 669454
rect 54566 669218 85050 669454
rect 85286 669218 115770 669454
rect 116006 669218 146490 669454
rect 146726 669218 177210 669454
rect 177446 669218 207930 669454
rect 208166 669218 238650 669454
rect 238886 669218 269370 669454
rect 269606 669218 300090 669454
rect 300326 669218 330810 669454
rect 331046 669218 361530 669454
rect 361766 669218 392250 669454
rect 392486 669218 422970 669454
rect 423206 669218 453690 669454
rect 453926 669218 484410 669454
rect 484646 669218 515130 669454
rect 515366 669218 545850 669454
rect 546086 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 23610 669134
rect 23846 668898 54330 669134
rect 54566 668898 85050 669134
rect 85286 668898 115770 669134
rect 116006 668898 146490 669134
rect 146726 668898 177210 669134
rect 177446 668898 207930 669134
rect 208166 668898 238650 669134
rect 238886 668898 269370 669134
rect 269606 668898 300090 669134
rect 300326 668898 330810 669134
rect 331046 668898 361530 669134
rect 361766 668898 392250 669134
rect 392486 668898 422970 669134
rect 423206 668898 453690 669134
rect 453926 668898 484410 669134
rect 484646 668898 515130 669134
rect 515366 668898 545850 669134
rect 546086 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 592650 662294
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 590730 658894
rect -6806 658574 590730 658658
rect -6806 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 590730 658574
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 588810 655174
rect -4886 654854 588810 654938
rect -4886 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 588810 654854
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 8250 651454
rect 8486 651218 38970 651454
rect 39206 651218 69690 651454
rect 69926 651218 100410 651454
rect 100646 651218 131130 651454
rect 131366 651218 161850 651454
rect 162086 651218 192570 651454
rect 192806 651218 223290 651454
rect 223526 651218 254010 651454
rect 254246 651218 284730 651454
rect 284966 651218 315450 651454
rect 315686 651218 346170 651454
rect 346406 651218 376890 651454
rect 377126 651218 407610 651454
rect 407846 651218 438330 651454
rect 438566 651218 469050 651454
rect 469286 651218 499770 651454
rect 500006 651218 530490 651454
rect 530726 651218 561210 651454
rect 561446 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 8250 651134
rect 8486 650898 38970 651134
rect 39206 650898 69690 651134
rect 69926 650898 100410 651134
rect 100646 650898 131130 651134
rect 131366 650898 161850 651134
rect 162086 650898 192570 651134
rect 192806 650898 223290 651134
rect 223526 650898 254010 651134
rect 254246 650898 284730 651134
rect 284966 650898 315450 651134
rect 315686 650898 346170 651134
rect 346406 650898 376890 651134
rect 377126 650898 407610 651134
rect 407846 650898 438330 651134
rect 438566 650898 469050 651134
rect 469286 650898 499770 651134
rect 500006 650898 530490 651134
rect 530726 650898 561210 651134
rect 561446 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect -8726 644294 592650 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect -6806 640574 590730 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect -4886 636854 588810 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 23610 633454
rect 23846 633218 54330 633454
rect 54566 633218 85050 633454
rect 85286 633218 115770 633454
rect 116006 633218 146490 633454
rect 146726 633218 177210 633454
rect 177446 633218 207930 633454
rect 208166 633218 238650 633454
rect 238886 633218 269370 633454
rect 269606 633218 300090 633454
rect 300326 633218 330810 633454
rect 331046 633218 361530 633454
rect 361766 633218 392250 633454
rect 392486 633218 422970 633454
rect 423206 633218 453690 633454
rect 453926 633218 484410 633454
rect 484646 633218 515130 633454
rect 515366 633218 545850 633454
rect 546086 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 23610 633134
rect 23846 632898 54330 633134
rect 54566 632898 85050 633134
rect 85286 632898 115770 633134
rect 116006 632898 146490 633134
rect 146726 632898 177210 633134
rect 177446 632898 207930 633134
rect 208166 632898 238650 633134
rect 238886 632898 269370 633134
rect 269606 632898 300090 633134
rect 300326 632898 330810 633134
rect 331046 632898 361530 633134
rect 361766 632898 392250 633134
rect 392486 632898 422970 633134
rect 423206 632898 453690 633134
rect 453926 632898 484410 633134
rect 484646 632898 515130 633134
rect 515366 632898 545850 633134
rect 546086 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 592650 626294
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 590730 622894
rect -6806 622574 590730 622658
rect -6806 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 590730 622574
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 588810 619174
rect -4886 618854 588810 618938
rect -4886 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 588810 618854
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 8250 615454
rect 8486 615218 38970 615454
rect 39206 615218 69690 615454
rect 69926 615218 100410 615454
rect 100646 615218 131130 615454
rect 131366 615218 161850 615454
rect 162086 615218 192570 615454
rect 192806 615218 223290 615454
rect 223526 615218 254010 615454
rect 254246 615218 284730 615454
rect 284966 615218 315450 615454
rect 315686 615218 346170 615454
rect 346406 615218 376890 615454
rect 377126 615218 407610 615454
rect 407846 615218 438330 615454
rect 438566 615218 469050 615454
rect 469286 615218 499770 615454
rect 500006 615218 530490 615454
rect 530726 615218 561210 615454
rect 561446 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 8250 615134
rect 8486 614898 38970 615134
rect 39206 614898 69690 615134
rect 69926 614898 100410 615134
rect 100646 614898 131130 615134
rect 131366 614898 161850 615134
rect 162086 614898 192570 615134
rect 192806 614898 223290 615134
rect 223526 614898 254010 615134
rect 254246 614898 284730 615134
rect 284966 614898 315450 615134
rect 315686 614898 346170 615134
rect 346406 614898 376890 615134
rect 377126 614898 407610 615134
rect 407846 614898 438330 615134
rect 438566 614898 469050 615134
rect 469286 614898 499770 615134
rect 500006 614898 530490 615134
rect 530726 614898 561210 615134
rect 561446 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect -8726 608294 592650 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect -6806 604574 590730 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect -4886 600854 588810 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 23610 597454
rect 23846 597218 54330 597454
rect 54566 597218 85050 597454
rect 85286 597218 115770 597454
rect 116006 597218 146490 597454
rect 146726 597218 177210 597454
rect 177446 597218 207930 597454
rect 208166 597218 238650 597454
rect 238886 597218 269370 597454
rect 269606 597218 300090 597454
rect 300326 597218 330810 597454
rect 331046 597218 361530 597454
rect 361766 597218 392250 597454
rect 392486 597218 422970 597454
rect 423206 597218 453690 597454
rect 453926 597218 484410 597454
rect 484646 597218 515130 597454
rect 515366 597218 545850 597454
rect 546086 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 23610 597134
rect 23846 596898 54330 597134
rect 54566 596898 85050 597134
rect 85286 596898 115770 597134
rect 116006 596898 146490 597134
rect 146726 596898 177210 597134
rect 177446 596898 207930 597134
rect 208166 596898 238650 597134
rect 238886 596898 269370 597134
rect 269606 596898 300090 597134
rect 300326 596898 330810 597134
rect 331046 596898 361530 597134
rect 361766 596898 392250 597134
rect 392486 596898 422970 597134
rect 423206 596898 453690 597134
rect 453926 596898 484410 597134
rect 484646 596898 515130 597134
rect 515366 596898 545850 597134
rect 546086 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 592650 590294
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 590730 586894
rect -6806 586574 590730 586658
rect -6806 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 590730 586574
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 588810 583174
rect -4886 582854 588810 582938
rect -4886 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 588810 582854
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 8250 579454
rect 8486 579218 38970 579454
rect 39206 579218 69690 579454
rect 69926 579218 100410 579454
rect 100646 579218 131130 579454
rect 131366 579218 161850 579454
rect 162086 579218 192570 579454
rect 192806 579218 223290 579454
rect 223526 579218 254010 579454
rect 254246 579218 284730 579454
rect 284966 579218 315450 579454
rect 315686 579218 346170 579454
rect 346406 579218 376890 579454
rect 377126 579218 407610 579454
rect 407846 579218 438330 579454
rect 438566 579218 469050 579454
rect 469286 579218 499770 579454
rect 500006 579218 530490 579454
rect 530726 579218 561210 579454
rect 561446 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 8250 579134
rect 8486 578898 38970 579134
rect 39206 578898 69690 579134
rect 69926 578898 100410 579134
rect 100646 578898 131130 579134
rect 131366 578898 161850 579134
rect 162086 578898 192570 579134
rect 192806 578898 223290 579134
rect 223526 578898 254010 579134
rect 254246 578898 284730 579134
rect 284966 578898 315450 579134
rect 315686 578898 346170 579134
rect 346406 578898 376890 579134
rect 377126 578898 407610 579134
rect 407846 578898 438330 579134
rect 438566 578898 469050 579134
rect 469286 578898 499770 579134
rect 500006 578898 530490 579134
rect 530726 578898 561210 579134
rect 561446 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect -8726 572294 592650 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect -6806 568574 590730 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect -4886 564854 588810 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect -4886 564586 588810 564618
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 23610 561454
rect 23846 561218 54330 561454
rect 54566 561218 85050 561454
rect 85286 561218 115770 561454
rect 116006 561218 146490 561454
rect 146726 561218 177210 561454
rect 177446 561218 207930 561454
rect 208166 561218 238650 561454
rect 238886 561218 269370 561454
rect 269606 561218 300090 561454
rect 300326 561218 330810 561454
rect 331046 561218 361530 561454
rect 361766 561218 392250 561454
rect 392486 561218 422970 561454
rect 423206 561218 453690 561454
rect 453926 561218 484410 561454
rect 484646 561218 515130 561454
rect 515366 561218 545850 561454
rect 546086 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 23610 561134
rect 23846 560898 54330 561134
rect 54566 560898 85050 561134
rect 85286 560898 115770 561134
rect 116006 560898 146490 561134
rect 146726 560898 177210 561134
rect 177446 560898 207930 561134
rect 208166 560898 238650 561134
rect 238886 560898 269370 561134
rect 269606 560898 300090 561134
rect 300326 560898 330810 561134
rect 331046 560898 361530 561134
rect 361766 560898 392250 561134
rect 392486 560898 422970 561134
rect 423206 560898 453690 561134
rect 453926 560898 484410 561134
rect 484646 560898 515130 561134
rect 515366 560898 545850 561134
rect 546086 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 592650 554294
rect -8726 554026 592650 554058
rect -6806 550894 590730 550926
rect -6806 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 590730 550894
rect -6806 550574 590730 550658
rect -6806 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 590730 550574
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 588810 547174
rect -4886 546854 588810 546938
rect -4886 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 588810 546854
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 8250 543454
rect 8486 543218 38970 543454
rect 39206 543218 69690 543454
rect 69926 543218 100410 543454
rect 100646 543218 131130 543454
rect 131366 543218 161850 543454
rect 162086 543218 192570 543454
rect 192806 543218 223290 543454
rect 223526 543218 254010 543454
rect 254246 543218 284730 543454
rect 284966 543218 315450 543454
rect 315686 543218 346170 543454
rect 346406 543218 376890 543454
rect 377126 543218 407610 543454
rect 407846 543218 438330 543454
rect 438566 543218 469050 543454
rect 469286 543218 499770 543454
rect 500006 543218 530490 543454
rect 530726 543218 561210 543454
rect 561446 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 8250 543134
rect 8486 542898 38970 543134
rect 39206 542898 69690 543134
rect 69926 542898 100410 543134
rect 100646 542898 131130 543134
rect 131366 542898 161850 543134
rect 162086 542898 192570 543134
rect 192806 542898 223290 543134
rect 223526 542898 254010 543134
rect 254246 542898 284730 543134
rect 284966 542898 315450 543134
rect 315686 542898 346170 543134
rect 346406 542898 376890 543134
rect 377126 542898 407610 543134
rect 407846 542898 438330 543134
rect 438566 542898 469050 543134
rect 469286 542898 499770 543134
rect 500006 542898 530490 543134
rect 530726 542898 561210 543134
rect 561446 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect -8726 536294 592650 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect -6806 532574 590730 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect -4886 528854 588810 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 23610 525454
rect 23846 525218 54330 525454
rect 54566 525218 85050 525454
rect 85286 525218 115770 525454
rect 116006 525218 146490 525454
rect 146726 525218 177210 525454
rect 177446 525218 207930 525454
rect 208166 525218 238650 525454
rect 238886 525218 269370 525454
rect 269606 525218 300090 525454
rect 300326 525218 330810 525454
rect 331046 525218 361530 525454
rect 361766 525218 392250 525454
rect 392486 525218 422970 525454
rect 423206 525218 453690 525454
rect 453926 525218 484410 525454
rect 484646 525218 515130 525454
rect 515366 525218 545850 525454
rect 546086 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 23610 525134
rect 23846 524898 54330 525134
rect 54566 524898 85050 525134
rect 85286 524898 115770 525134
rect 116006 524898 146490 525134
rect 146726 524898 177210 525134
rect 177446 524898 207930 525134
rect 208166 524898 238650 525134
rect 238886 524898 269370 525134
rect 269606 524898 300090 525134
rect 300326 524898 330810 525134
rect 331046 524898 361530 525134
rect 361766 524898 392250 525134
rect 392486 524898 422970 525134
rect 423206 524898 453690 525134
rect 453926 524898 484410 525134
rect 484646 524898 515130 525134
rect 515366 524898 545850 525134
rect 546086 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 592650 518294
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 590730 514894
rect -6806 514574 590730 514658
rect -6806 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 590730 514574
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 588810 511174
rect -4886 510854 588810 510938
rect -4886 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 588810 510854
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 8250 507454
rect 8486 507218 38970 507454
rect 39206 507218 69690 507454
rect 69926 507218 100410 507454
rect 100646 507218 131130 507454
rect 131366 507218 161850 507454
rect 162086 507218 192570 507454
rect 192806 507218 223290 507454
rect 223526 507218 254010 507454
rect 254246 507218 284730 507454
rect 284966 507218 315450 507454
rect 315686 507218 346170 507454
rect 346406 507218 376890 507454
rect 377126 507218 407610 507454
rect 407846 507218 438330 507454
rect 438566 507218 469050 507454
rect 469286 507218 499770 507454
rect 500006 507218 530490 507454
rect 530726 507218 561210 507454
rect 561446 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 8250 507134
rect 8486 506898 38970 507134
rect 39206 506898 69690 507134
rect 69926 506898 100410 507134
rect 100646 506898 131130 507134
rect 131366 506898 161850 507134
rect 162086 506898 192570 507134
rect 192806 506898 223290 507134
rect 223526 506898 254010 507134
rect 254246 506898 284730 507134
rect 284966 506898 315450 507134
rect 315686 506898 346170 507134
rect 346406 506898 376890 507134
rect 377126 506898 407610 507134
rect 407846 506898 438330 507134
rect 438566 506898 469050 507134
rect 469286 506898 499770 507134
rect 500006 506898 530490 507134
rect 530726 506898 561210 507134
rect 561446 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect -8726 500294 592650 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect -6806 496574 590730 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect -4886 492854 588810 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 23610 489454
rect 23846 489218 54330 489454
rect 54566 489218 85050 489454
rect 85286 489218 115770 489454
rect 116006 489218 146490 489454
rect 146726 489218 177210 489454
rect 177446 489218 207930 489454
rect 208166 489218 238650 489454
rect 238886 489218 269370 489454
rect 269606 489218 300090 489454
rect 300326 489218 330810 489454
rect 331046 489218 361530 489454
rect 361766 489218 392250 489454
rect 392486 489218 422970 489454
rect 423206 489218 453690 489454
rect 453926 489218 484410 489454
rect 484646 489218 515130 489454
rect 515366 489218 545850 489454
rect 546086 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 23610 489134
rect 23846 488898 54330 489134
rect 54566 488898 85050 489134
rect 85286 488898 115770 489134
rect 116006 488898 146490 489134
rect 146726 488898 177210 489134
rect 177446 488898 207930 489134
rect 208166 488898 238650 489134
rect 238886 488898 269370 489134
rect 269606 488898 300090 489134
rect 300326 488898 330810 489134
rect 331046 488898 361530 489134
rect 361766 488898 392250 489134
rect 392486 488898 422970 489134
rect 423206 488898 453690 489134
rect 453926 488898 484410 489134
rect 484646 488898 515130 489134
rect 515366 488898 545850 489134
rect 546086 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 592650 482294
rect -8726 482026 592650 482058
rect -6806 478894 590730 478926
rect -6806 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 590730 478894
rect -6806 478574 590730 478658
rect -6806 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 590730 478574
rect -6806 478306 590730 478338
rect -4886 475174 588810 475206
rect -4886 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 588810 475174
rect -4886 474854 588810 474938
rect -4886 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 588810 474854
rect -4886 474586 588810 474618
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 8250 471454
rect 8486 471218 38970 471454
rect 39206 471218 69690 471454
rect 69926 471218 100410 471454
rect 100646 471218 131130 471454
rect 131366 471218 161850 471454
rect 162086 471218 192570 471454
rect 192806 471218 223290 471454
rect 223526 471218 254010 471454
rect 254246 471218 284730 471454
rect 284966 471218 315450 471454
rect 315686 471218 346170 471454
rect 346406 471218 376890 471454
rect 377126 471218 407610 471454
rect 407846 471218 438330 471454
rect 438566 471218 469050 471454
rect 469286 471218 499770 471454
rect 500006 471218 530490 471454
rect 530726 471218 561210 471454
rect 561446 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 8250 471134
rect 8486 470898 38970 471134
rect 39206 470898 69690 471134
rect 69926 470898 100410 471134
rect 100646 470898 131130 471134
rect 131366 470898 161850 471134
rect 162086 470898 192570 471134
rect 192806 470898 223290 471134
rect 223526 470898 254010 471134
rect 254246 470898 284730 471134
rect 284966 470898 315450 471134
rect 315686 470898 346170 471134
rect 346406 470898 376890 471134
rect 377126 470898 407610 471134
rect 407846 470898 438330 471134
rect 438566 470898 469050 471134
rect 469286 470898 499770 471134
rect 500006 470898 530490 471134
rect 530726 470898 561210 471134
rect 561446 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect -8726 464294 592650 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect -6806 460574 590730 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect -4886 456854 588810 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 23610 453454
rect 23846 453218 54330 453454
rect 54566 453218 85050 453454
rect 85286 453218 115770 453454
rect 116006 453218 146490 453454
rect 146726 453218 177210 453454
rect 177446 453218 207930 453454
rect 208166 453218 238650 453454
rect 238886 453218 269370 453454
rect 269606 453218 300090 453454
rect 300326 453218 330810 453454
rect 331046 453218 361530 453454
rect 361766 453218 392250 453454
rect 392486 453218 422970 453454
rect 423206 453218 453690 453454
rect 453926 453218 484410 453454
rect 484646 453218 515130 453454
rect 515366 453218 545850 453454
rect 546086 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 23610 453134
rect 23846 452898 54330 453134
rect 54566 452898 85050 453134
rect 85286 452898 115770 453134
rect 116006 452898 146490 453134
rect 146726 452898 177210 453134
rect 177446 452898 207930 453134
rect 208166 452898 238650 453134
rect 238886 452898 269370 453134
rect 269606 452898 300090 453134
rect 300326 452898 330810 453134
rect 331046 452898 361530 453134
rect 361766 452898 392250 453134
rect 392486 452898 422970 453134
rect 423206 452898 453690 453134
rect 453926 452898 484410 453134
rect 484646 452898 515130 453134
rect 515366 452898 545850 453134
rect 546086 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 592650 446294
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 590730 442894
rect -6806 442574 590730 442658
rect -6806 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 590730 442574
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 588810 439174
rect -4886 438854 588810 438938
rect -4886 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 588810 438854
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 8250 435454
rect 8486 435218 38970 435454
rect 39206 435218 69690 435454
rect 69926 435218 100410 435454
rect 100646 435218 131130 435454
rect 131366 435218 161850 435454
rect 162086 435218 192570 435454
rect 192806 435218 223290 435454
rect 223526 435218 254010 435454
rect 254246 435218 284730 435454
rect 284966 435218 315450 435454
rect 315686 435218 346170 435454
rect 346406 435218 376890 435454
rect 377126 435218 407610 435454
rect 407846 435218 438330 435454
rect 438566 435218 469050 435454
rect 469286 435218 499770 435454
rect 500006 435218 530490 435454
rect 530726 435218 561210 435454
rect 561446 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 8250 435134
rect 8486 434898 38970 435134
rect 39206 434898 69690 435134
rect 69926 434898 100410 435134
rect 100646 434898 131130 435134
rect 131366 434898 161850 435134
rect 162086 434898 192570 435134
rect 192806 434898 223290 435134
rect 223526 434898 254010 435134
rect 254246 434898 284730 435134
rect 284966 434898 315450 435134
rect 315686 434898 346170 435134
rect 346406 434898 376890 435134
rect 377126 434898 407610 435134
rect 407846 434898 438330 435134
rect 438566 434898 469050 435134
rect 469286 434898 499770 435134
rect 500006 434898 530490 435134
rect 530726 434898 561210 435134
rect 561446 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect -8726 428294 592650 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect -6806 424574 590730 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect -4886 420854 588810 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 23610 417454
rect 23846 417218 54330 417454
rect 54566 417218 85050 417454
rect 85286 417218 115770 417454
rect 116006 417218 146490 417454
rect 146726 417218 177210 417454
rect 177446 417218 207930 417454
rect 208166 417218 238650 417454
rect 238886 417218 269370 417454
rect 269606 417218 300090 417454
rect 300326 417218 330810 417454
rect 331046 417218 361530 417454
rect 361766 417218 392250 417454
rect 392486 417218 422970 417454
rect 423206 417218 453690 417454
rect 453926 417218 484410 417454
rect 484646 417218 515130 417454
rect 515366 417218 545850 417454
rect 546086 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 23610 417134
rect 23846 416898 54330 417134
rect 54566 416898 85050 417134
rect 85286 416898 115770 417134
rect 116006 416898 146490 417134
rect 146726 416898 177210 417134
rect 177446 416898 207930 417134
rect 208166 416898 238650 417134
rect 238886 416898 269370 417134
rect 269606 416898 300090 417134
rect 300326 416898 330810 417134
rect 331046 416898 361530 417134
rect 361766 416898 392250 417134
rect 392486 416898 422970 417134
rect 423206 416898 453690 417134
rect 453926 416898 484410 417134
rect 484646 416898 515130 417134
rect 515366 416898 545850 417134
rect 546086 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 592650 410294
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 590730 406894
rect -6806 406574 590730 406658
rect -6806 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 590730 406574
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 588810 403174
rect -4886 402854 588810 402938
rect -4886 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 588810 402854
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 8250 399454
rect 8486 399218 38970 399454
rect 39206 399218 69690 399454
rect 69926 399218 100410 399454
rect 100646 399218 131130 399454
rect 131366 399218 161850 399454
rect 162086 399218 192570 399454
rect 192806 399218 223290 399454
rect 223526 399218 254010 399454
rect 254246 399218 284730 399454
rect 284966 399218 315450 399454
rect 315686 399218 346170 399454
rect 346406 399218 376890 399454
rect 377126 399218 407610 399454
rect 407846 399218 438330 399454
rect 438566 399218 469050 399454
rect 469286 399218 499770 399454
rect 500006 399218 530490 399454
rect 530726 399218 561210 399454
rect 561446 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 8250 399134
rect 8486 398898 38970 399134
rect 39206 398898 69690 399134
rect 69926 398898 100410 399134
rect 100646 398898 131130 399134
rect 131366 398898 161850 399134
rect 162086 398898 192570 399134
rect 192806 398898 223290 399134
rect 223526 398898 254010 399134
rect 254246 398898 284730 399134
rect 284966 398898 315450 399134
rect 315686 398898 346170 399134
rect 346406 398898 376890 399134
rect 377126 398898 407610 399134
rect 407846 398898 438330 399134
rect 438566 398898 469050 399134
rect 469286 398898 499770 399134
rect 500006 398898 530490 399134
rect 530726 398898 561210 399134
rect 561446 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect -8726 392294 592650 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect -8726 392026 592650 392058
rect -6806 388894 590730 388926
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect -6806 388574 590730 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect -4886 384854 588810 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 23610 381454
rect 23846 381218 54330 381454
rect 54566 381218 85050 381454
rect 85286 381218 115770 381454
rect 116006 381218 146490 381454
rect 146726 381218 177210 381454
rect 177446 381218 207930 381454
rect 208166 381218 238650 381454
rect 238886 381218 269370 381454
rect 269606 381218 300090 381454
rect 300326 381218 330810 381454
rect 331046 381218 361530 381454
rect 361766 381218 392250 381454
rect 392486 381218 422970 381454
rect 423206 381218 453690 381454
rect 453926 381218 484410 381454
rect 484646 381218 515130 381454
rect 515366 381218 545850 381454
rect 546086 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect -2966 381134 586890 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 23610 381134
rect 23846 380898 54330 381134
rect 54566 380898 85050 381134
rect 85286 380898 115770 381134
rect 116006 380898 146490 381134
rect 146726 380898 177210 381134
rect 177446 380898 207930 381134
rect 208166 380898 238650 381134
rect 238886 380898 269370 381134
rect 269606 380898 300090 381134
rect 300326 380898 330810 381134
rect 331046 380898 361530 381134
rect 361766 380898 392250 381134
rect 392486 380898 422970 381134
rect 423206 380898 453690 381134
rect 453926 380898 484410 381134
rect 484646 380898 515130 381134
rect 515366 380898 545850 381134
rect 546086 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 592650 374294
rect -8726 374026 592650 374058
rect -6806 370894 590730 370926
rect -6806 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 590730 370894
rect -6806 370574 590730 370658
rect -6806 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 590730 370574
rect -6806 370306 590730 370338
rect -4886 367174 588810 367206
rect -4886 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 588810 367174
rect -4886 366854 588810 366938
rect -4886 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 588810 366854
rect -4886 366586 588810 366618
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 8250 363454
rect 8486 363218 38970 363454
rect 39206 363218 69690 363454
rect 69926 363218 100410 363454
rect 100646 363218 131130 363454
rect 131366 363218 161850 363454
rect 162086 363218 192570 363454
rect 192806 363218 223290 363454
rect 223526 363218 254010 363454
rect 254246 363218 284730 363454
rect 284966 363218 315450 363454
rect 315686 363218 346170 363454
rect 346406 363218 376890 363454
rect 377126 363218 407610 363454
rect 407846 363218 438330 363454
rect 438566 363218 469050 363454
rect 469286 363218 499770 363454
rect 500006 363218 530490 363454
rect 530726 363218 561210 363454
rect 561446 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 8250 363134
rect 8486 362898 38970 363134
rect 39206 362898 69690 363134
rect 69926 362898 100410 363134
rect 100646 362898 131130 363134
rect 131366 362898 161850 363134
rect 162086 362898 192570 363134
rect 192806 362898 223290 363134
rect 223526 362898 254010 363134
rect 254246 362898 284730 363134
rect 284966 362898 315450 363134
rect 315686 362898 346170 363134
rect 346406 362898 376890 363134
rect 377126 362898 407610 363134
rect 407846 362898 438330 363134
rect 438566 362898 469050 363134
rect 469286 362898 499770 363134
rect 500006 362898 530490 363134
rect 530726 362898 561210 363134
rect 561446 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect -8726 356614 592650 356646
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect -8726 356294 592650 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect -6806 352574 590730 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect -4886 348854 588810 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect -4886 348586 588810 348618
rect -2966 345454 586890 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 23610 345454
rect 23846 345218 54330 345454
rect 54566 345218 85050 345454
rect 85286 345218 115770 345454
rect 116006 345218 146490 345454
rect 146726 345218 177210 345454
rect 177446 345218 207930 345454
rect 208166 345218 238650 345454
rect 238886 345218 269370 345454
rect 269606 345218 300090 345454
rect 300326 345218 330810 345454
rect 331046 345218 361530 345454
rect 361766 345218 392250 345454
rect 392486 345218 422970 345454
rect 423206 345218 453690 345454
rect 453926 345218 484410 345454
rect 484646 345218 515130 345454
rect 515366 345218 545850 345454
rect 546086 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect -2966 345134 586890 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 23610 345134
rect 23846 344898 54330 345134
rect 54566 344898 85050 345134
rect 85286 344898 115770 345134
rect 116006 344898 146490 345134
rect 146726 344898 177210 345134
rect 177446 344898 207930 345134
rect 208166 344898 238650 345134
rect 238886 344898 269370 345134
rect 269606 344898 300090 345134
rect 300326 344898 330810 345134
rect 331046 344898 361530 345134
rect 361766 344898 392250 345134
rect 392486 344898 422970 345134
rect 423206 344898 453690 345134
rect 453926 344898 484410 345134
rect 484646 344898 515130 345134
rect 515366 344898 545850 345134
rect 546086 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect -2966 344866 586890 344898
rect -8726 338614 592650 338646
rect -8726 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 592650 338294
rect -8726 338026 592650 338058
rect -6806 334894 590730 334926
rect -6806 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 590730 334894
rect -6806 334574 590730 334658
rect -6806 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 590730 334574
rect -6806 334306 590730 334338
rect -4886 331174 588810 331206
rect -4886 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 588810 331174
rect -4886 330854 588810 330938
rect -4886 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 588810 330854
rect -4886 330586 588810 330618
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 8250 327454
rect 8486 327218 38970 327454
rect 39206 327218 69690 327454
rect 69926 327218 100410 327454
rect 100646 327218 131130 327454
rect 131366 327218 161850 327454
rect 162086 327218 192570 327454
rect 192806 327218 223290 327454
rect 223526 327218 254010 327454
rect 254246 327218 284730 327454
rect 284966 327218 315450 327454
rect 315686 327218 346170 327454
rect 346406 327218 376890 327454
rect 377126 327218 407610 327454
rect 407846 327218 438330 327454
rect 438566 327218 469050 327454
rect 469286 327218 499770 327454
rect 500006 327218 530490 327454
rect 530726 327218 561210 327454
rect 561446 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 8250 327134
rect 8486 326898 38970 327134
rect 39206 326898 69690 327134
rect 69926 326898 100410 327134
rect 100646 326898 131130 327134
rect 131366 326898 161850 327134
rect 162086 326898 192570 327134
rect 192806 326898 223290 327134
rect 223526 326898 254010 327134
rect 254246 326898 284730 327134
rect 284966 326898 315450 327134
rect 315686 326898 346170 327134
rect 346406 326898 376890 327134
rect 377126 326898 407610 327134
rect 407846 326898 438330 327134
rect 438566 326898 469050 327134
rect 469286 326898 499770 327134
rect 500006 326898 530490 327134
rect 530726 326898 561210 327134
rect 561446 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect -8726 320294 592650 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect -6806 316574 590730 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect -4886 312854 588810 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 23610 309454
rect 23846 309218 54330 309454
rect 54566 309218 85050 309454
rect 85286 309218 115770 309454
rect 116006 309218 146490 309454
rect 146726 309218 177210 309454
rect 177446 309218 207930 309454
rect 208166 309218 238650 309454
rect 238886 309218 269370 309454
rect 269606 309218 300090 309454
rect 300326 309218 330810 309454
rect 331046 309218 361530 309454
rect 361766 309218 392250 309454
rect 392486 309218 422970 309454
rect 423206 309218 453690 309454
rect 453926 309218 484410 309454
rect 484646 309218 515130 309454
rect 515366 309218 545850 309454
rect 546086 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect -2966 309134 586890 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 23610 309134
rect 23846 308898 54330 309134
rect 54566 308898 85050 309134
rect 85286 308898 115770 309134
rect 116006 308898 146490 309134
rect 146726 308898 177210 309134
rect 177446 308898 207930 309134
rect 208166 308898 238650 309134
rect 238886 308898 269370 309134
rect 269606 308898 300090 309134
rect 300326 308898 330810 309134
rect 331046 308898 361530 309134
rect 361766 308898 392250 309134
rect 392486 308898 422970 309134
rect 423206 308898 453690 309134
rect 453926 308898 484410 309134
rect 484646 308898 515130 309134
rect 515366 308898 545850 309134
rect 546086 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect -2966 308866 586890 308898
rect -8726 302614 592650 302646
rect -8726 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 592650 302294
rect -8726 302026 592650 302058
rect -6806 298894 590730 298926
rect -6806 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 590730 298894
rect -6806 298574 590730 298658
rect -6806 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 590730 298574
rect -6806 298306 590730 298338
rect -4886 295174 588810 295206
rect -4886 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 588810 295174
rect -4886 294854 588810 294938
rect -4886 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 588810 294854
rect -4886 294586 588810 294618
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 8250 291454
rect 8486 291218 38970 291454
rect 39206 291218 69690 291454
rect 69926 291218 100410 291454
rect 100646 291218 131130 291454
rect 131366 291218 161850 291454
rect 162086 291218 192570 291454
rect 192806 291218 223290 291454
rect 223526 291218 254010 291454
rect 254246 291218 284730 291454
rect 284966 291218 315450 291454
rect 315686 291218 346170 291454
rect 346406 291218 376890 291454
rect 377126 291218 407610 291454
rect 407846 291218 438330 291454
rect 438566 291218 469050 291454
rect 469286 291218 499770 291454
rect 500006 291218 530490 291454
rect 530726 291218 561210 291454
rect 561446 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 8250 291134
rect 8486 290898 38970 291134
rect 39206 290898 69690 291134
rect 69926 290898 100410 291134
rect 100646 290898 131130 291134
rect 131366 290898 161850 291134
rect 162086 290898 192570 291134
rect 192806 290898 223290 291134
rect 223526 290898 254010 291134
rect 254246 290898 284730 291134
rect 284966 290898 315450 291134
rect 315686 290898 346170 291134
rect 346406 290898 376890 291134
rect 377126 290898 407610 291134
rect 407846 290898 438330 291134
rect 438566 290898 469050 291134
rect 469286 290898 499770 291134
rect 500006 290898 530490 291134
rect 530726 290898 561210 291134
rect 561446 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect -8726 284294 592650 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect -6806 280574 590730 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect -4886 276854 588810 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect -4886 276586 588810 276618
rect -2966 273454 586890 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 23610 273454
rect 23846 273218 54330 273454
rect 54566 273218 85050 273454
rect 85286 273218 115770 273454
rect 116006 273218 146490 273454
rect 146726 273218 177210 273454
rect 177446 273218 207930 273454
rect 208166 273218 238650 273454
rect 238886 273218 269370 273454
rect 269606 273218 300090 273454
rect 300326 273218 330810 273454
rect 331046 273218 361530 273454
rect 361766 273218 392250 273454
rect 392486 273218 422970 273454
rect 423206 273218 453690 273454
rect 453926 273218 484410 273454
rect 484646 273218 515130 273454
rect 515366 273218 545850 273454
rect 546086 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect -2966 273134 586890 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 23610 273134
rect 23846 272898 54330 273134
rect 54566 272898 85050 273134
rect 85286 272898 115770 273134
rect 116006 272898 146490 273134
rect 146726 272898 177210 273134
rect 177446 272898 207930 273134
rect 208166 272898 238650 273134
rect 238886 272898 269370 273134
rect 269606 272898 300090 273134
rect 300326 272898 330810 273134
rect 331046 272898 361530 273134
rect 361766 272898 392250 273134
rect 392486 272898 422970 273134
rect 423206 272898 453690 273134
rect 453926 272898 484410 273134
rect 484646 272898 515130 273134
rect 515366 272898 545850 273134
rect 546086 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 592650 266294
rect -8726 266026 592650 266058
rect -6806 262894 590730 262926
rect -6806 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 590730 262894
rect -6806 262574 590730 262658
rect -6806 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 590730 262574
rect -6806 262306 590730 262338
rect -4886 259174 588810 259206
rect -4886 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 588810 259174
rect -4886 258854 588810 258938
rect -4886 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 588810 258854
rect -4886 258586 588810 258618
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 8250 255454
rect 8486 255218 38970 255454
rect 39206 255218 69690 255454
rect 69926 255218 100410 255454
rect 100646 255218 131130 255454
rect 131366 255218 161850 255454
rect 162086 255218 192570 255454
rect 192806 255218 223290 255454
rect 223526 255218 254010 255454
rect 254246 255218 284730 255454
rect 284966 255218 315450 255454
rect 315686 255218 346170 255454
rect 346406 255218 376890 255454
rect 377126 255218 407610 255454
rect 407846 255218 438330 255454
rect 438566 255218 469050 255454
rect 469286 255218 499770 255454
rect 500006 255218 530490 255454
rect 530726 255218 561210 255454
rect 561446 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 8250 255134
rect 8486 254898 38970 255134
rect 39206 254898 69690 255134
rect 69926 254898 100410 255134
rect 100646 254898 131130 255134
rect 131366 254898 161850 255134
rect 162086 254898 192570 255134
rect 192806 254898 223290 255134
rect 223526 254898 254010 255134
rect 254246 254898 284730 255134
rect 284966 254898 315450 255134
rect 315686 254898 346170 255134
rect 346406 254898 376890 255134
rect 377126 254898 407610 255134
rect 407846 254898 438330 255134
rect 438566 254898 469050 255134
rect 469286 254898 499770 255134
rect 500006 254898 530490 255134
rect 530726 254898 561210 255134
rect 561446 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -8726 248614 592650 248646
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect -8726 248294 592650 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect -6806 244574 590730 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect -4886 240854 588810 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 23610 237454
rect 23846 237218 54330 237454
rect 54566 237218 85050 237454
rect 85286 237218 115770 237454
rect 116006 237218 146490 237454
rect 146726 237218 177210 237454
rect 177446 237218 207930 237454
rect 208166 237218 238650 237454
rect 238886 237218 269370 237454
rect 269606 237218 300090 237454
rect 300326 237218 330810 237454
rect 331046 237218 361530 237454
rect 361766 237218 392250 237454
rect 392486 237218 422970 237454
rect 423206 237218 453690 237454
rect 453926 237218 484410 237454
rect 484646 237218 515130 237454
rect 515366 237218 545850 237454
rect 546086 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect -2966 237134 586890 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 23610 237134
rect 23846 236898 54330 237134
rect 54566 236898 85050 237134
rect 85286 236898 115770 237134
rect 116006 236898 146490 237134
rect 146726 236898 177210 237134
rect 177446 236898 207930 237134
rect 208166 236898 238650 237134
rect 238886 236898 269370 237134
rect 269606 236898 300090 237134
rect 300326 236898 330810 237134
rect 331046 236898 361530 237134
rect 361766 236898 392250 237134
rect 392486 236898 422970 237134
rect 423206 236898 453690 237134
rect 453926 236898 484410 237134
rect 484646 236898 515130 237134
rect 515366 236898 545850 237134
rect 546086 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 592650 230294
rect -8726 230026 592650 230058
rect -6806 226894 590730 226926
rect -6806 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 590730 226894
rect -6806 226574 590730 226658
rect -6806 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 590730 226574
rect -6806 226306 590730 226338
rect -4886 223174 588810 223206
rect -4886 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 588810 223174
rect -4886 222854 588810 222938
rect -4886 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 588810 222854
rect -4886 222586 588810 222618
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 8250 219454
rect 8486 219218 38970 219454
rect 39206 219218 69690 219454
rect 69926 219218 100410 219454
rect 100646 219218 131130 219454
rect 131366 219218 161850 219454
rect 162086 219218 192570 219454
rect 192806 219218 223290 219454
rect 223526 219218 254010 219454
rect 254246 219218 284730 219454
rect 284966 219218 315450 219454
rect 315686 219218 346170 219454
rect 346406 219218 376890 219454
rect 377126 219218 407610 219454
rect 407846 219218 438330 219454
rect 438566 219218 469050 219454
rect 469286 219218 499770 219454
rect 500006 219218 530490 219454
rect 530726 219218 561210 219454
rect 561446 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 8250 219134
rect 8486 218898 38970 219134
rect 39206 218898 69690 219134
rect 69926 218898 100410 219134
rect 100646 218898 131130 219134
rect 131366 218898 161850 219134
rect 162086 218898 192570 219134
rect 192806 218898 223290 219134
rect 223526 218898 254010 219134
rect 254246 218898 284730 219134
rect 284966 218898 315450 219134
rect 315686 218898 346170 219134
rect 346406 218898 376890 219134
rect 377126 218898 407610 219134
rect 407846 218898 438330 219134
rect 438566 218898 469050 219134
rect 469286 218898 499770 219134
rect 500006 218898 530490 219134
rect 530726 218898 561210 219134
rect 561446 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -8726 212614 592650 212646
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect -8726 212294 592650 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect -6806 208574 590730 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect -4886 204854 588810 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 23610 201454
rect 23846 201218 54330 201454
rect 54566 201218 85050 201454
rect 85286 201218 115770 201454
rect 116006 201218 146490 201454
rect 146726 201218 177210 201454
rect 177446 201218 207930 201454
rect 208166 201218 238650 201454
rect 238886 201218 269370 201454
rect 269606 201218 300090 201454
rect 300326 201218 330810 201454
rect 331046 201218 361530 201454
rect 361766 201218 392250 201454
rect 392486 201218 422970 201454
rect 423206 201218 453690 201454
rect 453926 201218 484410 201454
rect 484646 201218 515130 201454
rect 515366 201218 545850 201454
rect 546086 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect -2966 201134 586890 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 23610 201134
rect 23846 200898 54330 201134
rect 54566 200898 85050 201134
rect 85286 200898 115770 201134
rect 116006 200898 146490 201134
rect 146726 200898 177210 201134
rect 177446 200898 207930 201134
rect 208166 200898 238650 201134
rect 238886 200898 269370 201134
rect 269606 200898 300090 201134
rect 300326 200898 330810 201134
rect 331046 200898 361530 201134
rect 361766 200898 392250 201134
rect 392486 200898 422970 201134
rect 423206 200898 453690 201134
rect 453926 200898 484410 201134
rect 484646 200898 515130 201134
rect 515366 200898 545850 201134
rect 546086 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 592650 194294
rect -8726 194026 592650 194058
rect -6806 190894 590730 190926
rect -6806 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 590730 190894
rect -6806 190574 590730 190658
rect -6806 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 590730 190574
rect -6806 190306 590730 190338
rect -4886 187174 588810 187206
rect -4886 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 588810 187174
rect -4886 186854 588810 186938
rect -4886 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 588810 186854
rect -4886 186586 588810 186618
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 8250 183454
rect 8486 183218 38970 183454
rect 39206 183218 69690 183454
rect 69926 183218 100410 183454
rect 100646 183218 131130 183454
rect 131366 183218 161850 183454
rect 162086 183218 192570 183454
rect 192806 183218 223290 183454
rect 223526 183218 254010 183454
rect 254246 183218 284730 183454
rect 284966 183218 315450 183454
rect 315686 183218 346170 183454
rect 346406 183218 376890 183454
rect 377126 183218 407610 183454
rect 407846 183218 438330 183454
rect 438566 183218 469050 183454
rect 469286 183218 499770 183454
rect 500006 183218 530490 183454
rect 530726 183218 561210 183454
rect 561446 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 8250 183134
rect 8486 182898 38970 183134
rect 39206 182898 69690 183134
rect 69926 182898 100410 183134
rect 100646 182898 131130 183134
rect 131366 182898 161850 183134
rect 162086 182898 192570 183134
rect 192806 182898 223290 183134
rect 223526 182898 254010 183134
rect 254246 182898 284730 183134
rect 284966 182898 315450 183134
rect 315686 182898 346170 183134
rect 346406 182898 376890 183134
rect 377126 182898 407610 183134
rect 407846 182898 438330 183134
rect 438566 182898 469050 183134
rect 469286 182898 499770 183134
rect 500006 182898 530490 183134
rect 530726 182898 561210 183134
rect 561446 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect -8726 176614 592650 176646
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect -8726 176294 592650 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect -8726 176026 592650 176058
rect -6806 172894 590730 172926
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect -6806 172574 590730 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect -6806 172306 590730 172338
rect -4886 169174 588810 169206
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect -4886 168854 588810 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect -4886 168586 588810 168618
rect -2966 165454 586890 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 23610 165454
rect 23846 165218 54330 165454
rect 54566 165218 85050 165454
rect 85286 165218 115770 165454
rect 116006 165218 146490 165454
rect 146726 165218 177210 165454
rect 177446 165218 207930 165454
rect 208166 165218 238650 165454
rect 238886 165218 269370 165454
rect 269606 165218 300090 165454
rect 300326 165218 330810 165454
rect 331046 165218 361530 165454
rect 361766 165218 392250 165454
rect 392486 165218 422970 165454
rect 423206 165218 453690 165454
rect 453926 165218 484410 165454
rect 484646 165218 515130 165454
rect 515366 165218 545850 165454
rect 546086 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect -2966 165134 586890 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 23610 165134
rect 23846 164898 54330 165134
rect 54566 164898 85050 165134
rect 85286 164898 115770 165134
rect 116006 164898 146490 165134
rect 146726 164898 177210 165134
rect 177446 164898 207930 165134
rect 208166 164898 238650 165134
rect 238886 164898 269370 165134
rect 269606 164898 300090 165134
rect 300326 164898 330810 165134
rect 331046 164898 361530 165134
rect 361766 164898 392250 165134
rect 392486 164898 422970 165134
rect 423206 164898 453690 165134
rect 453926 164898 484410 165134
rect 484646 164898 515130 165134
rect 515366 164898 545850 165134
rect 546086 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect -2966 164866 586890 164898
rect -8726 158614 592650 158646
rect -8726 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 592650 158294
rect -8726 158026 592650 158058
rect -6806 154894 590730 154926
rect -6806 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 590730 154894
rect -6806 154574 590730 154658
rect -6806 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 590730 154574
rect -6806 154306 590730 154338
rect -4886 151174 588810 151206
rect -4886 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 588810 151174
rect -4886 150854 588810 150938
rect -4886 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 588810 150854
rect -4886 150586 588810 150618
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 8250 147454
rect 8486 147218 38970 147454
rect 39206 147218 69690 147454
rect 69926 147218 100410 147454
rect 100646 147218 131130 147454
rect 131366 147218 161850 147454
rect 162086 147218 192570 147454
rect 192806 147218 223290 147454
rect 223526 147218 254010 147454
rect 254246 147218 284730 147454
rect 284966 147218 315450 147454
rect 315686 147218 346170 147454
rect 346406 147218 376890 147454
rect 377126 147218 407610 147454
rect 407846 147218 438330 147454
rect 438566 147218 469050 147454
rect 469286 147218 499770 147454
rect 500006 147218 530490 147454
rect 530726 147218 561210 147454
rect 561446 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 8250 147134
rect 8486 146898 38970 147134
rect 39206 146898 69690 147134
rect 69926 146898 100410 147134
rect 100646 146898 131130 147134
rect 131366 146898 161850 147134
rect 162086 146898 192570 147134
rect 192806 146898 223290 147134
rect 223526 146898 254010 147134
rect 254246 146898 284730 147134
rect 284966 146898 315450 147134
rect 315686 146898 346170 147134
rect 346406 146898 376890 147134
rect 377126 146898 407610 147134
rect 407846 146898 438330 147134
rect 438566 146898 469050 147134
rect 469286 146898 499770 147134
rect 500006 146898 530490 147134
rect 530726 146898 561210 147134
rect 561446 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -8726 140614 592650 140646
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect -8726 140294 592650 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect -8726 140026 592650 140058
rect -6806 136894 590730 136926
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect -6806 136574 590730 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect -6806 136306 590730 136338
rect -4886 133174 588810 133206
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect -4886 132854 588810 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect -4886 132586 588810 132618
rect -2966 129454 586890 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 23610 129454
rect 23846 129218 54330 129454
rect 54566 129218 85050 129454
rect 85286 129218 115770 129454
rect 116006 129218 146490 129454
rect 146726 129218 177210 129454
rect 177446 129218 207930 129454
rect 208166 129218 238650 129454
rect 238886 129218 269370 129454
rect 269606 129218 300090 129454
rect 300326 129218 330810 129454
rect 331046 129218 361530 129454
rect 361766 129218 392250 129454
rect 392486 129218 422970 129454
rect 423206 129218 453690 129454
rect 453926 129218 484410 129454
rect 484646 129218 515130 129454
rect 515366 129218 545850 129454
rect 546086 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect -2966 129134 586890 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 23610 129134
rect 23846 128898 54330 129134
rect 54566 128898 85050 129134
rect 85286 128898 115770 129134
rect 116006 128898 146490 129134
rect 146726 128898 177210 129134
rect 177446 128898 207930 129134
rect 208166 128898 238650 129134
rect 238886 128898 269370 129134
rect 269606 128898 300090 129134
rect 300326 128898 330810 129134
rect 331046 128898 361530 129134
rect 361766 128898 392250 129134
rect 392486 128898 422970 129134
rect 423206 128898 453690 129134
rect 453926 128898 484410 129134
rect 484646 128898 515130 129134
rect 515366 128898 545850 129134
rect 546086 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect -2966 128866 586890 128898
rect -8726 122614 592650 122646
rect -8726 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 592650 122294
rect -8726 122026 592650 122058
rect -6806 118894 590730 118926
rect -6806 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 590730 118894
rect -6806 118574 590730 118658
rect -6806 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 590730 118574
rect -6806 118306 590730 118338
rect -4886 115174 588810 115206
rect -4886 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 588810 115174
rect -4886 114854 588810 114938
rect -4886 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 588810 114854
rect -4886 114586 588810 114618
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 8250 111454
rect 8486 111218 38970 111454
rect 39206 111218 69690 111454
rect 69926 111218 100410 111454
rect 100646 111218 131130 111454
rect 131366 111218 161850 111454
rect 162086 111218 192570 111454
rect 192806 111218 223290 111454
rect 223526 111218 254010 111454
rect 254246 111218 284730 111454
rect 284966 111218 315450 111454
rect 315686 111218 346170 111454
rect 346406 111218 376890 111454
rect 377126 111218 407610 111454
rect 407846 111218 438330 111454
rect 438566 111218 469050 111454
rect 469286 111218 499770 111454
rect 500006 111218 530490 111454
rect 530726 111218 561210 111454
rect 561446 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 8250 111134
rect 8486 110898 38970 111134
rect 39206 110898 69690 111134
rect 69926 110898 100410 111134
rect 100646 110898 131130 111134
rect 131366 110898 161850 111134
rect 162086 110898 192570 111134
rect 192806 110898 223290 111134
rect 223526 110898 254010 111134
rect 254246 110898 284730 111134
rect 284966 110898 315450 111134
rect 315686 110898 346170 111134
rect 346406 110898 376890 111134
rect 377126 110898 407610 111134
rect 407846 110898 438330 111134
rect 438566 110898 469050 111134
rect 469286 110898 499770 111134
rect 500006 110898 530490 111134
rect 530726 110898 561210 111134
rect 561446 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -8726 104614 592650 104646
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect -8726 104294 592650 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect -8726 104026 592650 104058
rect -6806 100894 590730 100926
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect -6806 100574 590730 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect -6806 100306 590730 100338
rect -4886 97174 588810 97206
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect -4886 96854 588810 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect -4886 96586 588810 96618
rect -2966 93454 586890 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 23610 93454
rect 23846 93218 54330 93454
rect 54566 93218 85050 93454
rect 85286 93218 115770 93454
rect 116006 93218 146490 93454
rect 146726 93218 177210 93454
rect 177446 93218 207930 93454
rect 208166 93218 238650 93454
rect 238886 93218 269370 93454
rect 269606 93218 300090 93454
rect 300326 93218 330810 93454
rect 331046 93218 361530 93454
rect 361766 93218 392250 93454
rect 392486 93218 422970 93454
rect 423206 93218 453690 93454
rect 453926 93218 484410 93454
rect 484646 93218 515130 93454
rect 515366 93218 545850 93454
rect 546086 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect -2966 93134 586890 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 23610 93134
rect 23846 92898 54330 93134
rect 54566 92898 85050 93134
rect 85286 92898 115770 93134
rect 116006 92898 146490 93134
rect 146726 92898 177210 93134
rect 177446 92898 207930 93134
rect 208166 92898 238650 93134
rect 238886 92898 269370 93134
rect 269606 92898 300090 93134
rect 300326 92898 330810 93134
rect 331046 92898 361530 93134
rect 361766 92898 392250 93134
rect 392486 92898 422970 93134
rect 423206 92898 453690 93134
rect 453926 92898 484410 93134
rect 484646 92898 515130 93134
rect 515366 92898 545850 93134
rect 546086 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect -2966 92866 586890 92898
rect -8726 86614 592650 86646
rect -8726 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 592650 86294
rect -8726 86026 592650 86058
rect -6806 82894 590730 82926
rect -6806 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 590730 82894
rect -6806 82574 590730 82658
rect -6806 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 590730 82574
rect -6806 82306 590730 82338
rect -4886 79174 588810 79206
rect -4886 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 588810 79174
rect -4886 78854 588810 78938
rect -4886 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 588810 78854
rect -4886 78586 588810 78618
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 8250 75454
rect 8486 75218 38970 75454
rect 39206 75218 69690 75454
rect 69926 75218 100410 75454
rect 100646 75218 131130 75454
rect 131366 75218 161850 75454
rect 162086 75218 192570 75454
rect 192806 75218 223290 75454
rect 223526 75218 254010 75454
rect 254246 75218 284730 75454
rect 284966 75218 315450 75454
rect 315686 75218 346170 75454
rect 346406 75218 376890 75454
rect 377126 75218 407610 75454
rect 407846 75218 438330 75454
rect 438566 75218 469050 75454
rect 469286 75218 499770 75454
rect 500006 75218 530490 75454
rect 530726 75218 561210 75454
rect 561446 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 8250 75134
rect 8486 74898 38970 75134
rect 39206 74898 69690 75134
rect 69926 74898 100410 75134
rect 100646 74898 131130 75134
rect 131366 74898 161850 75134
rect 162086 74898 192570 75134
rect 192806 74898 223290 75134
rect 223526 74898 254010 75134
rect 254246 74898 284730 75134
rect 284966 74898 315450 75134
rect 315686 74898 346170 75134
rect 346406 74898 376890 75134
rect 377126 74898 407610 75134
rect 407846 74898 438330 75134
rect 438566 74898 469050 75134
rect 469286 74898 499770 75134
rect 500006 74898 530490 75134
rect 530726 74898 561210 75134
rect 561446 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -8726 68614 592650 68646
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect -8726 68294 592650 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect -8726 68026 592650 68058
rect -6806 64894 590730 64926
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect -6806 64574 590730 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect -6806 64306 590730 64338
rect -4886 61174 588810 61206
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect -4886 60854 588810 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect -4886 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 23610 57454
rect 23846 57218 54330 57454
rect 54566 57218 85050 57454
rect 85286 57218 115770 57454
rect 116006 57218 146490 57454
rect 146726 57218 177210 57454
rect 177446 57218 207930 57454
rect 208166 57218 238650 57454
rect 238886 57218 269370 57454
rect 269606 57218 300090 57454
rect 300326 57218 330810 57454
rect 331046 57218 361530 57454
rect 361766 57218 392250 57454
rect 392486 57218 422970 57454
rect 423206 57218 453690 57454
rect 453926 57218 484410 57454
rect 484646 57218 515130 57454
rect 515366 57218 545850 57454
rect 546086 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 23610 57134
rect 23846 56898 54330 57134
rect 54566 56898 85050 57134
rect 85286 56898 115770 57134
rect 116006 56898 146490 57134
rect 146726 56898 177210 57134
rect 177446 56898 207930 57134
rect 208166 56898 238650 57134
rect 238886 56898 269370 57134
rect 269606 56898 300090 57134
rect 300326 56898 330810 57134
rect 331046 56898 361530 57134
rect 361766 56898 392250 57134
rect 392486 56898 422970 57134
rect 423206 56898 453690 57134
rect 453926 56898 484410 57134
rect 484646 56898 515130 57134
rect 515366 56898 545850 57134
rect 546086 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 592650 50294
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 590730 46894
rect -6806 46574 590730 46658
rect -6806 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 590730 46574
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 588810 43174
rect -4886 42854 588810 42938
rect -4886 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 588810 42854
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 8250 39454
rect 8486 39218 38970 39454
rect 39206 39218 69690 39454
rect 69926 39218 100410 39454
rect 100646 39218 131130 39454
rect 131366 39218 161850 39454
rect 162086 39218 192570 39454
rect 192806 39218 223290 39454
rect 223526 39218 254010 39454
rect 254246 39218 284730 39454
rect 284966 39218 315450 39454
rect 315686 39218 346170 39454
rect 346406 39218 376890 39454
rect 377126 39218 407610 39454
rect 407846 39218 438330 39454
rect 438566 39218 469050 39454
rect 469286 39218 499770 39454
rect 500006 39218 530490 39454
rect 530726 39218 561210 39454
rect 561446 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 8250 39134
rect 8486 38898 38970 39134
rect 39206 38898 69690 39134
rect 69926 38898 100410 39134
rect 100646 38898 131130 39134
rect 131366 38898 161850 39134
rect 162086 38898 192570 39134
rect 192806 38898 223290 39134
rect 223526 38898 254010 39134
rect 254246 38898 284730 39134
rect 284966 38898 315450 39134
rect 315686 38898 346170 39134
rect 346406 38898 376890 39134
rect 377126 38898 407610 39134
rect 407846 38898 438330 39134
rect 438566 38898 469050 39134
rect 469286 38898 499770 39134
rect 500006 38898 530490 39134
rect 530726 38898 561210 39134
rect 561446 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect -8726 32294 592650 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect -6806 28574 590730 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect -4886 24854 588810 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 23610 21454
rect 23846 21218 54330 21454
rect 54566 21218 85050 21454
rect 85286 21218 115770 21454
rect 116006 21218 146490 21454
rect 146726 21218 177210 21454
rect 177446 21218 207930 21454
rect 208166 21218 238650 21454
rect 238886 21218 269370 21454
rect 269606 21218 300090 21454
rect 300326 21218 330810 21454
rect 331046 21218 361530 21454
rect 361766 21218 392250 21454
rect 392486 21218 422970 21454
rect 423206 21218 453690 21454
rect 453926 21218 484410 21454
rect 484646 21218 515130 21454
rect 515366 21218 545850 21454
rect 546086 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 23610 21134
rect 23846 20898 54330 21134
rect 54566 20898 85050 21134
rect 85286 20898 115770 21134
rect 116006 20898 146490 21134
rect 146726 20898 177210 21134
rect 177446 20898 207930 21134
rect 208166 20898 238650 21134
rect 238886 20898 269370 21134
rect 269606 20898 300090 21134
rect 300326 20898 330810 21134
rect 331046 20898 361530 21134
rect 361766 20898 392250 21134
rect 392486 20898 422970 21134
rect 423206 20898 453690 21134
rect 453926 20898 484410 21134
rect 484646 20898 515130 21134
rect 515366 20898 545850 21134
rect 546086 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 592650 14294
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 590730 10894
rect -6806 10574 590730 10658
rect -6806 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 590730 10574
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 588810 7174
rect -4886 6854 588810 6938
rect -4886 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 588810 6854
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 8250 3454
rect 8486 3218 38970 3454
rect 39206 3218 69690 3454
rect 69926 3218 100410 3454
rect 100646 3218 131130 3454
rect 131366 3218 161850 3454
rect 162086 3218 192570 3454
rect 192806 3218 223290 3454
rect 223526 3218 254010 3454
rect 254246 3218 284730 3454
rect 284966 3218 315450 3454
rect 315686 3218 346170 3454
rect 346406 3218 376890 3454
rect 377126 3218 407610 3454
rect 407846 3218 438330 3454
rect 438566 3218 469050 3454
rect 469286 3218 499770 3454
rect 500006 3218 530490 3454
rect 530726 3218 561210 3454
rect 561446 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 8250 3134
rect 8486 2898 38970 3134
rect 39206 2898 69690 3134
rect 69926 2898 100410 3134
rect 100646 2898 131130 3134
rect 131366 2898 161850 3134
rect 162086 2898 192570 3134
rect 192806 2898 223290 3134
rect 223526 2898 254010 3134
rect 254246 2898 284730 3134
rect 284966 2898 315450 3134
rect 315686 2898 346170 3134
rect 346406 2898 376890 3134
rect 377126 2898 407610 3134
rect 407846 2898 438330 3134
rect 438566 2898 469050 3134
rect 469286 2898 499770 3134
rect 500006 2898 530490 3134
rect 530726 2898 561210 3134
rect 561446 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use user_proj  mprj
timestamp 1638672285
transform 1 0 4000 0 1 0
box 566 0 559438 700000
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 702000 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 702000 38414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 702000 74414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 702000 110414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 702000 146414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 702000 182414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 702000 218414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 702000 254414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 702000 290414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 702000 326414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 702000 362414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 702000 398414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 702000 434414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 702000 470414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 702000 506414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 702000 542414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 -3814 6134 -2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 41514 -3814 42134 -2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 77514 -3814 78134 -2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 113514 -3814 114134 -2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 149514 -3814 150134 -2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 185514 -3814 186134 -2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 221514 -3814 222134 -2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 257514 -3814 258134 -2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 293514 -3814 294134 -2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 329514 -3814 330134 -2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 365514 -3814 366134 -2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 401514 -3814 402134 -2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 437514 -3814 438134 -2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 473514 -3814 474134 -2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 509514 -3814 510134 -2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 545514 -3814 546134 -2000 8 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 702000 6134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 702000 42134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 702000 78134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 702000 114134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 702000 150134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 702000 186134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 702000 222134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 702000 258134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 702000 294134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 702000 330134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 702000 366134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 702000 402134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 702000 438134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 702000 474134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 702000 510134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 702000 546134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 581514 -3814 582134 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 -5734 9854 -2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 45234 -5734 45854 -2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 81234 -5734 81854 -2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 117234 -5734 117854 -2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 153234 -5734 153854 -2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 189234 -5734 189854 -2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 225234 -5734 225854 -2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 261234 -5734 261854 -2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 297234 -5734 297854 -2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 333234 -5734 333854 -2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 369234 -5734 369854 -2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 405234 -5734 405854 -2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 441234 -5734 441854 -2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 477234 -5734 477854 -2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 513234 -5734 513854 -2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 549234 -5734 549854 -2000 8 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 702000 9854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 702000 45854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 702000 81854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 702000 117854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 702000 153854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 702000 189854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 702000 225854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 702000 261854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 702000 297854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 702000 333854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 702000 369854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 702000 405854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 702000 441854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 702000 477854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 702000 513854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 702000 549854 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 -7654 13574 -2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 48954 -7654 49574 -2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 84954 -7654 85574 -2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 120954 -7654 121574 -2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 156954 -7654 157574 -2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 192954 -7654 193574 -2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 228954 -7654 229574 -2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 264954 -7654 265574 -2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 300954 -7654 301574 -2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 336954 -7654 337574 -2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 372954 -7654 373574 -2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 408954 -7654 409574 -2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 444954 -7654 445574 -2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 480954 -7654 481574 -2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 516954 -7654 517574 -2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 552954 -7654 553574 -2000 8 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 702000 13574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 702000 49574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 702000 85574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 702000 121574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 702000 157574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 702000 193574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 702000 229574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 702000 265574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 702000 301574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 702000 337574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 702000 373574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 702000 409574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 702000 445574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 702000 481574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 702000 517574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 702000 553574 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 -5734 27854 -2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 -5734 63854 -2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 -5734 99854 -2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 -5734 135854 -2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 -5734 171854 -2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 -5734 207854 -2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 -5734 243854 -2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 -5734 279854 -2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 -5734 315854 -2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 -5734 351854 -2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 -5734 387854 -2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 -5734 423854 -2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 -5734 459854 -2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 -5734 495854 -2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 -5734 531854 -2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 702000 27854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 702000 63854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 702000 99854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 702000 135854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 702000 171854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 702000 207854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 702000 243854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 702000 279854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 702000 315854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 702000 351854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 702000 387854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 702000 423854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 702000 459854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 702000 495854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 702000 531854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 -5734 567854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 -7654 31574 -2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 -7654 67574 -2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 -7654 103574 -2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 -7654 139574 -2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 -7654 175574 -2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 -7654 211574 -2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 -7654 247574 -2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 -7654 283574 -2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 -7654 319574 -2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 -7654 355574 -2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 -7654 391574 -2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 -7654 427574 -2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 -7654 463574 -2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 -7654 499574 -2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 -7654 535574 -2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 702000 31574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 702000 67574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 702000 103574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 702000 139574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 702000 175574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 702000 211574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 702000 247574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 702000 283574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 702000 319574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 702000 355574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 702000 391574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 702000 427574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 702000 463574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 702000 499574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 702000 535574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 -7654 571574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 702000 20414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 702000 56414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 702000 92414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 702000 128414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 702000 164414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 702000 200414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 702000 236414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 702000 272414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 702000 308414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 702000 344414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 702000 380414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 702000 416414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 702000 452414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 702000 488414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 702000 524414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 702000 560414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 -3814 24134 -2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 -3814 60134 -2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 -3814 96134 -2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 -3814 132134 -2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 -3814 168134 -2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 -3814 204134 -2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 -3814 240134 -2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 -3814 276134 -2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 -3814 312134 -2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 -3814 348134 -2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 -3814 384134 -2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 -3814 420134 -2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 -3814 456134 -2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 -3814 492134 -2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 -3814 528134 -2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 -3814 564134 -2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 702000 24134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 702000 60134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 702000 96134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 702000 132134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 702000 168134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 702000 204134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 702000 240134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 702000 276134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 702000 312134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 702000 348134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 702000 384134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 702000 420134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 702000 456134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 702000 492134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 702000 528134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 702000 564134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
