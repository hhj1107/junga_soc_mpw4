magic
tech sky130A
magscale 1 2
timestamp 1641207128
<< obsli1 >>
rect 1104 2159 178267 178449
<< obsm1 >>
rect 842 1164 178650 180736
<< metal2 >>
rect 570 180003 626 180803
rect 1674 180003 1730 180803
rect 2778 180003 2834 180803
rect 3882 180003 3938 180803
rect 4986 180003 5042 180803
rect 6090 180003 6146 180803
rect 7194 180003 7250 180803
rect 8298 180003 8354 180803
rect 9494 180003 9550 180803
rect 10598 180003 10654 180803
rect 11702 180003 11758 180803
rect 12806 180003 12862 180803
rect 13910 180003 13966 180803
rect 15014 180003 15070 180803
rect 16118 180003 16174 180803
rect 17314 180003 17370 180803
rect 18418 180003 18474 180803
rect 19522 180003 19578 180803
rect 20626 180003 20682 180803
rect 21730 180003 21786 180803
rect 22834 180003 22890 180803
rect 23938 180003 23994 180803
rect 25134 180003 25190 180803
rect 26238 180003 26294 180803
rect 27342 180003 27398 180803
rect 28446 180003 28502 180803
rect 29550 180003 29606 180803
rect 30654 180003 30710 180803
rect 31758 180003 31814 180803
rect 32862 180003 32918 180803
rect 34058 180003 34114 180803
rect 35162 180003 35218 180803
rect 36266 180003 36322 180803
rect 37370 180003 37426 180803
rect 38474 180003 38530 180803
rect 39578 180003 39634 180803
rect 40682 180003 40738 180803
rect 41878 180003 41934 180803
rect 42982 180003 43038 180803
rect 44086 180003 44142 180803
rect 45190 180003 45246 180803
rect 46294 180003 46350 180803
rect 47398 180003 47454 180803
rect 48502 180003 48558 180803
rect 49698 180003 49754 180803
rect 50802 180003 50858 180803
rect 51906 180003 51962 180803
rect 53010 180003 53066 180803
rect 54114 180003 54170 180803
rect 55218 180003 55274 180803
rect 56322 180003 56378 180803
rect 57518 180003 57574 180803
rect 58622 180003 58678 180803
rect 59726 180003 59782 180803
rect 60830 180003 60886 180803
rect 61934 180003 61990 180803
rect 63038 180003 63094 180803
rect 64142 180003 64198 180803
rect 65246 180003 65302 180803
rect 66442 180003 66498 180803
rect 67546 180003 67602 180803
rect 68650 180003 68706 180803
rect 69754 180003 69810 180803
rect 70858 180003 70914 180803
rect 71962 180003 72018 180803
rect 73066 180003 73122 180803
rect 74262 180003 74318 180803
rect 75366 180003 75422 180803
rect 76470 180003 76526 180803
rect 77574 180003 77630 180803
rect 78678 180003 78734 180803
rect 79782 180003 79838 180803
rect 80886 180003 80942 180803
rect 82082 180003 82138 180803
rect 83186 180003 83242 180803
rect 84290 180003 84346 180803
rect 85394 180003 85450 180803
rect 86498 180003 86554 180803
rect 87602 180003 87658 180803
rect 88706 180003 88762 180803
rect 89902 180003 89958 180803
rect 91006 180003 91062 180803
rect 92110 180003 92166 180803
rect 93214 180003 93270 180803
rect 94318 180003 94374 180803
rect 95422 180003 95478 180803
rect 96526 180003 96582 180803
rect 97630 180003 97686 180803
rect 98826 180003 98882 180803
rect 99930 180003 99986 180803
rect 101034 180003 101090 180803
rect 102138 180003 102194 180803
rect 103242 180003 103298 180803
rect 104346 180003 104402 180803
rect 105450 180003 105506 180803
rect 106646 180003 106702 180803
rect 107750 180003 107806 180803
rect 108854 180003 108910 180803
rect 109958 180003 110014 180803
rect 111062 180003 111118 180803
rect 112166 180003 112222 180803
rect 113270 180003 113326 180803
rect 114466 180003 114522 180803
rect 115570 180003 115626 180803
rect 116674 180003 116730 180803
rect 117778 180003 117834 180803
rect 118882 180003 118938 180803
rect 119986 180003 120042 180803
rect 121090 180003 121146 180803
rect 122194 180003 122250 180803
rect 123390 180003 123446 180803
rect 124494 180003 124550 180803
rect 125598 180003 125654 180803
rect 126702 180003 126758 180803
rect 127806 180003 127862 180803
rect 128910 180003 128966 180803
rect 130014 180003 130070 180803
rect 131210 180003 131266 180803
rect 132314 180003 132370 180803
rect 133418 180003 133474 180803
rect 134522 180003 134578 180803
rect 135626 180003 135682 180803
rect 136730 180003 136786 180803
rect 137834 180003 137890 180803
rect 139030 180003 139086 180803
rect 140134 180003 140190 180803
rect 141238 180003 141294 180803
rect 142342 180003 142398 180803
rect 143446 180003 143502 180803
rect 144550 180003 144606 180803
rect 145654 180003 145710 180803
rect 146850 180003 146906 180803
rect 147954 180003 148010 180803
rect 149058 180003 149114 180803
rect 150162 180003 150218 180803
rect 151266 180003 151322 180803
rect 152370 180003 152426 180803
rect 153474 180003 153530 180803
rect 154578 180003 154634 180803
rect 155774 180003 155830 180803
rect 156878 180003 156934 180803
rect 157982 180003 158038 180803
rect 159086 180003 159142 180803
rect 160190 180003 160246 180803
rect 161294 180003 161350 180803
rect 162398 180003 162454 180803
rect 163594 180003 163650 180803
rect 164698 180003 164754 180803
rect 165802 180003 165858 180803
rect 166906 180003 166962 180803
rect 168010 180003 168066 180803
rect 169114 180003 169170 180803
rect 170218 180003 170274 180803
rect 171414 180003 171470 180803
rect 172518 180003 172574 180803
rect 173622 180003 173678 180803
rect 174726 180003 174782 180803
rect 175830 180003 175886 180803
rect 176934 180003 176990 180803
rect 178038 180003 178094 180803
rect 570 0 626 800
rect 1766 0 1822 800
rect 3054 0 3110 800
rect 4342 0 4398 800
rect 5630 0 5686 800
rect 6918 0 6974 800
rect 8206 0 8262 800
rect 9494 0 9550 800
rect 10782 0 10838 800
rect 12070 0 12126 800
rect 13358 0 13414 800
rect 14646 0 14702 800
rect 15934 0 15990 800
rect 17222 0 17278 800
rect 18510 0 18566 800
rect 19798 0 19854 800
rect 21086 0 21142 800
rect 22374 0 22430 800
rect 23662 0 23718 800
rect 24950 0 25006 800
rect 26238 0 26294 800
rect 27526 0 27582 800
rect 28814 0 28870 800
rect 30102 0 30158 800
rect 31390 0 31446 800
rect 32678 0 32734 800
rect 33966 0 34022 800
rect 35254 0 35310 800
rect 36542 0 36598 800
rect 37830 0 37886 800
rect 39118 0 39174 800
rect 40406 0 40462 800
rect 41694 0 41750 800
rect 42982 0 43038 800
rect 44270 0 44326 800
rect 45466 0 45522 800
rect 46754 0 46810 800
rect 48042 0 48098 800
rect 49330 0 49386 800
rect 50618 0 50674 800
rect 51906 0 51962 800
rect 53194 0 53250 800
rect 54482 0 54538 800
rect 55770 0 55826 800
rect 57058 0 57114 800
rect 58346 0 58402 800
rect 59634 0 59690 800
rect 60922 0 60978 800
rect 62210 0 62266 800
rect 63498 0 63554 800
rect 64786 0 64842 800
rect 66074 0 66130 800
rect 67362 0 67418 800
rect 68650 0 68706 800
rect 69938 0 69994 800
rect 71226 0 71282 800
rect 72514 0 72570 800
rect 73802 0 73858 800
rect 75090 0 75146 800
rect 76378 0 76434 800
rect 77666 0 77722 800
rect 78954 0 79010 800
rect 80242 0 80298 800
rect 81530 0 81586 800
rect 82818 0 82874 800
rect 84106 0 84162 800
rect 85394 0 85450 800
rect 86682 0 86738 800
rect 87970 0 88026 800
rect 89258 0 89314 800
rect 90454 0 90510 800
rect 91742 0 91798 800
rect 93030 0 93086 800
rect 94318 0 94374 800
rect 95606 0 95662 800
rect 96894 0 96950 800
rect 98182 0 98238 800
rect 99470 0 99526 800
rect 100758 0 100814 800
rect 102046 0 102102 800
rect 103334 0 103390 800
rect 104622 0 104678 800
rect 105910 0 105966 800
rect 107198 0 107254 800
rect 108486 0 108542 800
rect 109774 0 109830 800
rect 111062 0 111118 800
rect 112350 0 112406 800
rect 113638 0 113694 800
rect 114926 0 114982 800
rect 116214 0 116270 800
rect 117502 0 117558 800
rect 118790 0 118846 800
rect 120078 0 120134 800
rect 121366 0 121422 800
rect 122654 0 122710 800
rect 123942 0 123998 800
rect 125230 0 125286 800
rect 126518 0 126574 800
rect 127806 0 127862 800
rect 129094 0 129150 800
rect 130382 0 130438 800
rect 131670 0 131726 800
rect 132958 0 133014 800
rect 134246 0 134302 800
rect 135442 0 135498 800
rect 136730 0 136786 800
rect 138018 0 138074 800
rect 139306 0 139362 800
rect 140594 0 140650 800
rect 141882 0 141938 800
rect 143170 0 143226 800
rect 144458 0 144514 800
rect 145746 0 145802 800
rect 147034 0 147090 800
rect 148322 0 148378 800
rect 149610 0 149666 800
rect 150898 0 150954 800
rect 152186 0 152242 800
rect 153474 0 153530 800
rect 154762 0 154818 800
rect 156050 0 156106 800
rect 157338 0 157394 800
rect 158626 0 158682 800
rect 159914 0 159970 800
rect 161202 0 161258 800
rect 162490 0 162546 800
rect 163778 0 163834 800
rect 165066 0 165122 800
rect 166354 0 166410 800
rect 167642 0 167698 800
rect 168930 0 168986 800
rect 170218 0 170274 800
rect 171506 0 171562 800
rect 172794 0 172850 800
rect 174082 0 174138 800
rect 175370 0 175426 800
rect 176658 0 176714 800
rect 177946 0 178002 800
<< obsm2 >>
rect 18 179947 514 180742
rect 682 179947 1618 180742
rect 1786 179947 2722 180742
rect 2890 179947 3826 180742
rect 3994 179947 4930 180742
rect 5098 179947 6034 180742
rect 6202 179947 7138 180742
rect 7306 179947 8242 180742
rect 8410 179947 9438 180742
rect 9606 179947 10542 180742
rect 10710 179947 11646 180742
rect 11814 179947 12750 180742
rect 12918 179947 13854 180742
rect 14022 179947 14958 180742
rect 15126 179947 16062 180742
rect 16230 179947 17258 180742
rect 17426 179947 18362 180742
rect 18530 179947 19466 180742
rect 19634 179947 20570 180742
rect 20738 179947 21674 180742
rect 21842 179947 22778 180742
rect 22946 179947 23882 180742
rect 24050 179947 25078 180742
rect 25246 179947 26182 180742
rect 26350 179947 27286 180742
rect 27454 179947 28390 180742
rect 28558 179947 29494 180742
rect 29662 179947 30598 180742
rect 30766 179947 31702 180742
rect 31870 179947 32806 180742
rect 32974 179947 34002 180742
rect 34170 179947 35106 180742
rect 35274 179947 36210 180742
rect 36378 179947 37314 180742
rect 37482 179947 38418 180742
rect 38586 179947 39522 180742
rect 39690 179947 40626 180742
rect 40794 179947 41822 180742
rect 41990 179947 42926 180742
rect 43094 179947 44030 180742
rect 44198 179947 45134 180742
rect 45302 179947 46238 180742
rect 46406 179947 47342 180742
rect 47510 179947 48446 180742
rect 48614 179947 49642 180742
rect 49810 179947 50746 180742
rect 50914 179947 51850 180742
rect 52018 179947 52954 180742
rect 53122 179947 54058 180742
rect 54226 179947 55162 180742
rect 55330 179947 56266 180742
rect 56434 179947 57462 180742
rect 57630 179947 58566 180742
rect 58734 179947 59670 180742
rect 59838 179947 60774 180742
rect 60942 179947 61878 180742
rect 62046 179947 62982 180742
rect 63150 179947 64086 180742
rect 64254 179947 65190 180742
rect 65358 179947 66386 180742
rect 66554 179947 67490 180742
rect 67658 179947 68594 180742
rect 68762 179947 69698 180742
rect 69866 179947 70802 180742
rect 70970 179947 71906 180742
rect 72074 179947 73010 180742
rect 73178 179947 74206 180742
rect 74374 179947 75310 180742
rect 75478 179947 76414 180742
rect 76582 179947 77518 180742
rect 77686 179947 78622 180742
rect 78790 179947 79726 180742
rect 79894 179947 80830 180742
rect 80998 179947 82026 180742
rect 82194 179947 83130 180742
rect 83298 179947 84234 180742
rect 84402 179947 85338 180742
rect 85506 179947 86442 180742
rect 86610 179947 87546 180742
rect 87714 179947 88650 180742
rect 88818 179947 89846 180742
rect 90014 179947 90950 180742
rect 91118 179947 92054 180742
rect 92222 179947 93158 180742
rect 93326 179947 94262 180742
rect 94430 179947 95366 180742
rect 95534 179947 96470 180742
rect 96638 179947 97574 180742
rect 97742 179947 98770 180742
rect 98938 179947 99874 180742
rect 100042 179947 100978 180742
rect 101146 179947 102082 180742
rect 102250 179947 103186 180742
rect 103354 179947 104290 180742
rect 104458 179947 105394 180742
rect 105562 179947 106590 180742
rect 106758 179947 107694 180742
rect 107862 179947 108798 180742
rect 108966 179947 109902 180742
rect 110070 179947 111006 180742
rect 111174 179947 112110 180742
rect 112278 179947 113214 180742
rect 113382 179947 114410 180742
rect 114578 179947 115514 180742
rect 115682 179947 116618 180742
rect 116786 179947 117722 180742
rect 117890 179947 118826 180742
rect 118994 179947 119930 180742
rect 120098 179947 121034 180742
rect 121202 179947 122138 180742
rect 122306 179947 123334 180742
rect 123502 179947 124438 180742
rect 124606 179947 125542 180742
rect 125710 179947 126646 180742
rect 126814 179947 127750 180742
rect 127918 179947 128854 180742
rect 129022 179947 129958 180742
rect 130126 179947 131154 180742
rect 131322 179947 132258 180742
rect 132426 179947 133362 180742
rect 133530 179947 134466 180742
rect 134634 179947 135570 180742
rect 135738 179947 136674 180742
rect 136842 179947 137778 180742
rect 137946 179947 138974 180742
rect 139142 179947 140078 180742
rect 140246 179947 141182 180742
rect 141350 179947 142286 180742
rect 142454 179947 143390 180742
rect 143558 179947 144494 180742
rect 144662 179947 145598 180742
rect 145766 179947 146794 180742
rect 146962 179947 147898 180742
rect 148066 179947 149002 180742
rect 149170 179947 150106 180742
rect 150274 179947 151210 180742
rect 151378 179947 152314 180742
rect 152482 179947 153418 180742
rect 153586 179947 154522 180742
rect 154690 179947 155718 180742
rect 155886 179947 156822 180742
rect 156990 179947 157926 180742
rect 158094 179947 159030 180742
rect 159198 179947 160134 180742
rect 160302 179947 161238 180742
rect 161406 179947 162342 180742
rect 162510 179947 163538 180742
rect 163706 179947 164642 180742
rect 164810 179947 165746 180742
rect 165914 179947 166850 180742
rect 167018 179947 167954 180742
rect 168122 179947 169058 180742
rect 169226 179947 170162 180742
rect 170330 179947 171358 180742
rect 171526 179947 172462 180742
rect 172630 179947 173566 180742
rect 173734 179947 174670 180742
rect 174838 179947 175774 180742
rect 175942 179947 176878 180742
rect 177046 179947 177982 180742
rect 178150 179947 178646 180742
rect 18 856 178646 179947
rect 18 734 514 856
rect 682 734 1710 856
rect 1878 734 2998 856
rect 3166 734 4286 856
rect 4454 734 5574 856
rect 5742 734 6862 856
rect 7030 734 8150 856
rect 8318 734 9438 856
rect 9606 734 10726 856
rect 10894 734 12014 856
rect 12182 734 13302 856
rect 13470 734 14590 856
rect 14758 734 15878 856
rect 16046 734 17166 856
rect 17334 734 18454 856
rect 18622 734 19742 856
rect 19910 734 21030 856
rect 21198 734 22318 856
rect 22486 734 23606 856
rect 23774 734 24894 856
rect 25062 734 26182 856
rect 26350 734 27470 856
rect 27638 734 28758 856
rect 28926 734 30046 856
rect 30214 734 31334 856
rect 31502 734 32622 856
rect 32790 734 33910 856
rect 34078 734 35198 856
rect 35366 734 36486 856
rect 36654 734 37774 856
rect 37942 734 39062 856
rect 39230 734 40350 856
rect 40518 734 41638 856
rect 41806 734 42926 856
rect 43094 734 44214 856
rect 44382 734 45410 856
rect 45578 734 46698 856
rect 46866 734 47986 856
rect 48154 734 49274 856
rect 49442 734 50562 856
rect 50730 734 51850 856
rect 52018 734 53138 856
rect 53306 734 54426 856
rect 54594 734 55714 856
rect 55882 734 57002 856
rect 57170 734 58290 856
rect 58458 734 59578 856
rect 59746 734 60866 856
rect 61034 734 62154 856
rect 62322 734 63442 856
rect 63610 734 64730 856
rect 64898 734 66018 856
rect 66186 734 67306 856
rect 67474 734 68594 856
rect 68762 734 69882 856
rect 70050 734 71170 856
rect 71338 734 72458 856
rect 72626 734 73746 856
rect 73914 734 75034 856
rect 75202 734 76322 856
rect 76490 734 77610 856
rect 77778 734 78898 856
rect 79066 734 80186 856
rect 80354 734 81474 856
rect 81642 734 82762 856
rect 82930 734 84050 856
rect 84218 734 85338 856
rect 85506 734 86626 856
rect 86794 734 87914 856
rect 88082 734 89202 856
rect 89370 734 90398 856
rect 90566 734 91686 856
rect 91854 734 92974 856
rect 93142 734 94262 856
rect 94430 734 95550 856
rect 95718 734 96838 856
rect 97006 734 98126 856
rect 98294 734 99414 856
rect 99582 734 100702 856
rect 100870 734 101990 856
rect 102158 734 103278 856
rect 103446 734 104566 856
rect 104734 734 105854 856
rect 106022 734 107142 856
rect 107310 734 108430 856
rect 108598 734 109718 856
rect 109886 734 111006 856
rect 111174 734 112294 856
rect 112462 734 113582 856
rect 113750 734 114870 856
rect 115038 734 116158 856
rect 116326 734 117446 856
rect 117614 734 118734 856
rect 118902 734 120022 856
rect 120190 734 121310 856
rect 121478 734 122598 856
rect 122766 734 123886 856
rect 124054 734 125174 856
rect 125342 734 126462 856
rect 126630 734 127750 856
rect 127918 734 129038 856
rect 129206 734 130326 856
rect 130494 734 131614 856
rect 131782 734 132902 856
rect 133070 734 134190 856
rect 134358 734 135386 856
rect 135554 734 136674 856
rect 136842 734 137962 856
rect 138130 734 139250 856
rect 139418 734 140538 856
rect 140706 734 141826 856
rect 141994 734 143114 856
rect 143282 734 144402 856
rect 144570 734 145690 856
rect 145858 734 146978 856
rect 147146 734 148266 856
rect 148434 734 149554 856
rect 149722 734 150842 856
rect 151010 734 152130 856
rect 152298 734 153418 856
rect 153586 734 154706 856
rect 154874 734 155994 856
rect 156162 734 157282 856
rect 157450 734 158570 856
rect 158738 734 159858 856
rect 160026 734 161146 856
rect 161314 734 162434 856
rect 162602 734 163722 856
rect 163890 734 165010 856
rect 165178 734 166298 856
rect 166466 734 167586 856
rect 167754 734 168874 856
rect 169042 734 170162 856
rect 170330 734 171450 856
rect 171618 734 172738 856
rect 172906 734 174026 856
rect 174194 734 175314 856
rect 175482 734 176602 856
rect 176770 734 177890 856
rect 178058 734 178646 856
<< metal3 >>
rect 177859 178576 178659 178696
rect 0 178304 800 178424
rect 177859 174496 178659 174616
rect 0 173680 800 173800
rect 177859 170552 178659 170672
rect 0 169056 800 169176
rect 177859 166472 178659 166592
rect 0 164432 800 164552
rect 177859 162528 178659 162648
rect 0 159808 800 159928
rect 177859 158448 178659 158568
rect 0 155184 800 155304
rect 177859 154504 178659 154624
rect 0 150560 800 150680
rect 177859 150424 178659 150544
rect 177859 146480 178659 146600
rect 0 145936 800 146056
rect 177859 142400 178659 142520
rect 0 141312 800 141432
rect 177859 138456 178659 138576
rect 0 136688 800 136808
rect 177859 134376 178659 134496
rect 0 132064 800 132184
rect 177859 130432 178659 130552
rect 0 127440 800 127560
rect 177859 126352 178659 126472
rect 0 122816 800 122936
rect 177859 122408 178659 122528
rect 177859 118328 178659 118448
rect 0 118056 800 118176
rect 177859 114248 178659 114368
rect 0 113432 800 113552
rect 177859 110304 178659 110424
rect 0 108808 800 108928
rect 177859 106224 178659 106344
rect 0 104184 800 104304
rect 177859 102280 178659 102400
rect 0 99560 800 99680
rect 177859 98200 178659 98320
rect 0 94936 800 95056
rect 177859 94256 178659 94376
rect 0 90312 800 90432
rect 177859 90176 178659 90296
rect 177859 86232 178659 86352
rect 0 85688 800 85808
rect 177859 82152 178659 82272
rect 0 81064 800 81184
rect 177859 78208 178659 78328
rect 0 76440 800 76560
rect 177859 74128 178659 74248
rect 0 71816 800 71936
rect 177859 70184 178659 70304
rect 0 67192 800 67312
rect 177859 66104 178659 66224
rect 0 62568 800 62688
rect 177859 62160 178659 62280
rect 177859 58080 178659 58200
rect 0 57808 800 57928
rect 177859 54000 178659 54120
rect 0 53184 800 53304
rect 177859 50056 178659 50176
rect 0 48560 800 48680
rect 177859 45976 178659 46096
rect 0 43936 800 44056
rect 177859 42032 178659 42152
rect 0 39312 800 39432
rect 177859 37952 178659 38072
rect 0 34688 800 34808
rect 177859 34008 178659 34128
rect 0 30064 800 30184
rect 177859 29928 178659 30048
rect 177859 25984 178659 26104
rect 0 25440 800 25560
rect 177859 21904 178659 22024
rect 0 20816 800 20936
rect 177859 17960 178659 18080
rect 0 16192 800 16312
rect 177859 13880 178659 14000
rect 0 11568 800 11688
rect 177859 9936 178659 10056
rect 0 6944 800 7064
rect 177859 5856 178659 5976
rect 0 2320 800 2440
rect 177859 1912 178659 2032
<< obsm3 >>
rect 13 178776 178651 180709
rect 13 178504 177779 178776
rect 880 178496 177779 178504
rect 880 178224 178651 178496
rect 13 174696 178651 178224
rect 13 174416 177779 174696
rect 13 173880 178651 174416
rect 880 173600 178651 173880
rect 13 170752 178651 173600
rect 13 170472 177779 170752
rect 13 169256 178651 170472
rect 880 168976 178651 169256
rect 13 166672 178651 168976
rect 13 166392 177779 166672
rect 13 164632 178651 166392
rect 880 164352 178651 164632
rect 13 162728 178651 164352
rect 13 162448 177779 162728
rect 13 160008 178651 162448
rect 880 159728 178651 160008
rect 13 158648 178651 159728
rect 13 158368 177779 158648
rect 13 155384 178651 158368
rect 880 155104 178651 155384
rect 13 154704 178651 155104
rect 13 154424 177779 154704
rect 13 150760 178651 154424
rect 880 150624 178651 150760
rect 880 150480 177779 150624
rect 13 150344 177779 150480
rect 13 146680 178651 150344
rect 13 146400 177779 146680
rect 13 146136 178651 146400
rect 880 145856 178651 146136
rect 13 142600 178651 145856
rect 13 142320 177779 142600
rect 13 141512 178651 142320
rect 880 141232 178651 141512
rect 13 138656 178651 141232
rect 13 138376 177779 138656
rect 13 136888 178651 138376
rect 880 136608 178651 136888
rect 13 134576 178651 136608
rect 13 134296 177779 134576
rect 13 132264 178651 134296
rect 880 131984 178651 132264
rect 13 130632 178651 131984
rect 13 130352 177779 130632
rect 13 127640 178651 130352
rect 880 127360 178651 127640
rect 13 126552 178651 127360
rect 13 126272 177779 126552
rect 13 123016 178651 126272
rect 880 122736 178651 123016
rect 13 122608 178651 122736
rect 13 122328 177779 122608
rect 13 118528 178651 122328
rect 13 118256 177779 118528
rect 880 118248 177779 118256
rect 880 117976 178651 118248
rect 13 114448 178651 117976
rect 13 114168 177779 114448
rect 13 113632 178651 114168
rect 880 113352 178651 113632
rect 13 110504 178651 113352
rect 13 110224 177779 110504
rect 13 109008 178651 110224
rect 880 108728 178651 109008
rect 13 106424 178651 108728
rect 13 106144 177779 106424
rect 13 104384 178651 106144
rect 880 104104 178651 104384
rect 13 102480 178651 104104
rect 13 102200 177779 102480
rect 13 99760 178651 102200
rect 880 99480 178651 99760
rect 13 98400 178651 99480
rect 13 98120 177779 98400
rect 13 95136 178651 98120
rect 880 94856 178651 95136
rect 13 94456 178651 94856
rect 13 94176 177779 94456
rect 13 90512 178651 94176
rect 880 90376 178651 90512
rect 880 90232 177779 90376
rect 13 90096 177779 90232
rect 13 86432 178651 90096
rect 13 86152 177779 86432
rect 13 85888 178651 86152
rect 880 85608 178651 85888
rect 13 82352 178651 85608
rect 13 82072 177779 82352
rect 13 81264 178651 82072
rect 880 80984 178651 81264
rect 13 78408 178651 80984
rect 13 78128 177779 78408
rect 13 76640 178651 78128
rect 880 76360 178651 76640
rect 13 74328 178651 76360
rect 13 74048 177779 74328
rect 13 72016 178651 74048
rect 880 71736 178651 72016
rect 13 70384 178651 71736
rect 13 70104 177779 70384
rect 13 67392 178651 70104
rect 880 67112 178651 67392
rect 13 66304 178651 67112
rect 13 66024 177779 66304
rect 13 62768 178651 66024
rect 880 62488 178651 62768
rect 13 62360 178651 62488
rect 13 62080 177779 62360
rect 13 58280 178651 62080
rect 13 58008 177779 58280
rect 880 58000 177779 58008
rect 880 57728 178651 58000
rect 13 54200 178651 57728
rect 13 53920 177779 54200
rect 13 53384 178651 53920
rect 880 53104 178651 53384
rect 13 50256 178651 53104
rect 13 49976 177779 50256
rect 13 48760 178651 49976
rect 880 48480 178651 48760
rect 13 46176 178651 48480
rect 13 45896 177779 46176
rect 13 44136 178651 45896
rect 880 43856 178651 44136
rect 13 42232 178651 43856
rect 13 41952 177779 42232
rect 13 39512 178651 41952
rect 880 39232 178651 39512
rect 13 38152 178651 39232
rect 13 37872 177779 38152
rect 13 34888 178651 37872
rect 880 34608 178651 34888
rect 13 34208 178651 34608
rect 13 33928 177779 34208
rect 13 30264 178651 33928
rect 880 30128 178651 30264
rect 880 29984 177779 30128
rect 13 29848 177779 29984
rect 13 26184 178651 29848
rect 13 25904 177779 26184
rect 13 25640 178651 25904
rect 880 25360 178651 25640
rect 13 22104 178651 25360
rect 13 21824 177779 22104
rect 13 21016 178651 21824
rect 880 20736 178651 21016
rect 13 18160 178651 20736
rect 13 17880 177779 18160
rect 13 16392 178651 17880
rect 880 16112 178651 16392
rect 13 14080 178651 16112
rect 13 13800 177779 14080
rect 13 11768 178651 13800
rect 880 11488 178651 11768
rect 13 10136 178651 11488
rect 13 9856 177779 10136
rect 13 7144 178651 9856
rect 880 6864 178651 7144
rect 13 6056 178651 6864
rect 13 5776 177779 6056
rect 13 2520 178651 5776
rect 880 2240 178651 2520
rect 13 2112 178651 2240
rect 13 1939 177779 2112
<< metal4 >>
rect 4208 2128 4528 178480
rect 19568 2128 19888 178480
rect 34928 2128 35248 178480
rect 50288 2128 50608 178480
rect 65648 2128 65968 178480
rect 81008 2128 81328 178480
rect 96368 2128 96688 178480
rect 111728 2128 112048 178480
rect 127088 2128 127408 178480
rect 142448 2128 142768 178480
rect 157808 2128 158128 178480
rect 173168 2128 173488 178480
<< obsm4 >>
rect 19379 178560 175845 180709
rect 19379 5339 19488 178560
rect 19968 5339 34848 178560
rect 35328 5339 50208 178560
rect 50688 5339 65568 178560
rect 66048 5339 80928 178560
rect 81408 5339 96288 178560
rect 96768 5339 111648 178560
rect 112128 5339 127008 178560
rect 127488 5339 142368 178560
rect 142848 5339 157728 178560
rect 158208 5339 173088 178560
rect 173568 5339 175845 178560
<< labels >>
rlabel metal2 s 127806 180003 127862 180803 6 clk_i
port 1 nsew signal input
rlabel metal2 s 130014 180003 130070 180803 6 i_dout0[0]
port 2 nsew signal input
rlabel metal2 s 156050 0 156106 800 6 i_dout0[10]
port 3 nsew signal input
rlabel metal2 s 157338 0 157394 800 6 i_dout0[11]
port 4 nsew signal input
rlabel metal3 s 0 113432 800 113552 6 i_dout0[12]
port 5 nsew signal input
rlabel metal2 s 150162 180003 150218 180803 6 i_dout0[13]
port 6 nsew signal input
rlabel metal2 s 161202 0 161258 800 6 i_dout0[14]
port 7 nsew signal input
rlabel metal2 s 152370 180003 152426 180803 6 i_dout0[15]
port 8 nsew signal input
rlabel metal3 s 177859 114248 178659 114368 6 i_dout0[16]
port 9 nsew signal input
rlabel metal2 s 154578 180003 154634 180803 6 i_dout0[17]
port 10 nsew signal input
rlabel metal3 s 177859 118328 178659 118448 6 i_dout0[18]
port 11 nsew signal input
rlabel metal3 s 0 136688 800 136808 6 i_dout0[19]
port 12 nsew signal input
rlabel metal2 s 143170 0 143226 800 6 i_dout0[1]
port 13 nsew signal input
rlabel metal3 s 177859 130432 178659 130552 6 i_dout0[20]
port 14 nsew signal input
rlabel metal2 s 161294 180003 161350 180803 6 i_dout0[21]
port 15 nsew signal input
rlabel metal2 s 168930 0 168986 800 6 i_dout0[22]
port 16 nsew signal input
rlabel metal3 s 0 150560 800 150680 6 i_dout0[23]
port 17 nsew signal input
rlabel metal2 s 170218 0 170274 800 6 i_dout0[24]
port 18 nsew signal input
rlabel metal3 s 177859 154504 178659 154624 6 i_dout0[25]
port 19 nsew signal input
rlabel metal3 s 0 159808 800 159928 6 i_dout0[26]
port 20 nsew signal input
rlabel metal2 s 170218 180003 170274 180803 6 i_dout0[27]
port 21 nsew signal input
rlabel metal3 s 177859 166472 178659 166592 6 i_dout0[28]
port 22 nsew signal input
rlabel metal2 s 175830 180003 175886 180803 6 i_dout0[29]
port 23 nsew signal input
rlabel metal2 s 144458 0 144514 800 6 i_dout0[2]
port 24 nsew signal input
rlabel metal3 s 177859 174496 178659 174616 6 i_dout0[30]
port 25 nsew signal input
rlabel metal3 s 177859 178576 178659 178696 6 i_dout0[31]
port 26 nsew signal input
rlabel metal3 s 0 34688 800 34808 6 i_dout0[3]
port 27 nsew signal input
rlabel metal3 s 177859 42032 178659 42152 6 i_dout0[4]
port 28 nsew signal input
rlabel metal3 s 0 67192 800 67312 6 i_dout0[5]
port 29 nsew signal input
rlabel metal2 s 150898 0 150954 800 6 i_dout0[6]
port 30 nsew signal input
rlabel metal3 s 177859 54000 178659 54120 6 i_dout0[7]
port 31 nsew signal input
rlabel metal2 s 145654 180003 145710 180803 6 i_dout0[8]
port 32 nsew signal input
rlabel metal2 s 147954 180003 148010 180803 6 i_dout0[9]
port 33 nsew signal input
rlabel metal3 s 177859 13880 178659 14000 6 i_dout0_1[0]
port 34 nsew signal input
rlabel metal3 s 0 99560 800 99680 6 i_dout0_1[10]
port 35 nsew signal input
rlabel metal3 s 0 108808 800 108928 6 i_dout0_1[11]
port 36 nsew signal input
rlabel metal3 s 177859 90176 178659 90296 6 i_dout0_1[12]
port 37 nsew signal input
rlabel metal2 s 149058 180003 149114 180803 6 i_dout0_1[13]
port 38 nsew signal input
rlabel metal3 s 0 122816 800 122936 6 i_dout0_1[14]
port 39 nsew signal input
rlabel metal2 s 151266 180003 151322 180803 6 i_dout0_1[15]
port 40 nsew signal input
rlabel metal3 s 177859 110304 178659 110424 6 i_dout0_1[16]
port 41 nsew signal input
rlabel metal2 s 165066 0 165122 800 6 i_dout0_1[17]
port 42 nsew signal input
rlabel metal2 s 156878 180003 156934 180803 6 i_dout0_1[18]
port 43 nsew signal input
rlabel metal3 s 177859 126352 178659 126472 6 i_dout0_1[19]
port 44 nsew signal input
rlabel metal2 s 141882 0 141938 800 6 i_dout0_1[1]
port 45 nsew signal input
rlabel metal3 s 0 141312 800 141432 6 i_dout0_1[20]
port 46 nsew signal input
rlabel metal2 s 167642 0 167698 800 6 i_dout0_1[21]
port 47 nsew signal input
rlabel metal3 s 177859 138456 178659 138576 6 i_dout0_1[22]
port 48 nsew signal input
rlabel metal3 s 177859 142400 178659 142520 6 i_dout0_1[23]
port 49 nsew signal input
rlabel metal3 s 177859 146480 178659 146600 6 i_dout0_1[24]
port 50 nsew signal input
rlabel metal2 s 171506 0 171562 800 6 i_dout0_1[25]
port 51 nsew signal input
rlabel metal3 s 177859 158448 178659 158568 6 i_dout0_1[26]
port 52 nsew signal input
rlabel metal3 s 177859 162528 178659 162648 6 i_dout0_1[27]
port 53 nsew signal input
rlabel metal2 s 173622 180003 173678 180803 6 i_dout0_1[28]
port 54 nsew signal input
rlabel metal3 s 0 164432 800 164552 6 i_dout0_1[29]
port 55 nsew signal input
rlabel metal2 s 135626 180003 135682 180803 6 i_dout0_1[2]
port 56 nsew signal input
rlabel metal2 s 175370 0 175426 800 6 i_dout0_1[30]
port 57 nsew signal input
rlabel metal2 s 176658 0 176714 800 6 i_dout0_1[31]
port 58 nsew signal input
rlabel metal2 s 145746 0 145802 800 6 i_dout0_1[3]
port 59 nsew signal input
rlabel metal2 s 147034 0 147090 800 6 i_dout0_1[4]
port 60 nsew signal input
rlabel metal3 s 0 62568 800 62688 6 i_dout0_1[5]
port 61 nsew signal input
rlabel metal3 s 0 81064 800 81184 6 i_dout0_1[6]
port 62 nsew signal input
rlabel metal2 s 153474 0 153530 800 6 i_dout0_1[7]
port 63 nsew signal input
rlabel metal3 s 177859 70184 178659 70304 6 i_dout0_1[8]
port 64 nsew signal input
rlabel metal3 s 0 90312 800 90432 6 i_dout0_1[9]
port 65 nsew signal input
rlabel metal2 s 570 180003 626 180803 6 io_in[0]
port 66 nsew signal input
rlabel metal2 s 34058 180003 34114 180803 6 io_in[10]
port 67 nsew signal input
rlabel metal2 s 37370 180003 37426 180803 6 io_in[11]
port 68 nsew signal input
rlabel metal2 s 40682 180003 40738 180803 6 io_in[12]
port 69 nsew signal input
rlabel metal2 s 44086 180003 44142 180803 6 io_in[13]
port 70 nsew signal input
rlabel metal2 s 47398 180003 47454 180803 6 io_in[14]
port 71 nsew signal input
rlabel metal2 s 50802 180003 50858 180803 6 io_in[15]
port 72 nsew signal input
rlabel metal2 s 54114 180003 54170 180803 6 io_in[16]
port 73 nsew signal input
rlabel metal2 s 57518 180003 57574 180803 6 io_in[17]
port 74 nsew signal input
rlabel metal2 s 60830 180003 60886 180803 6 io_in[18]
port 75 nsew signal input
rlabel metal2 s 64142 180003 64198 180803 6 io_in[19]
port 76 nsew signal input
rlabel metal2 s 3882 180003 3938 180803 6 io_in[1]
port 77 nsew signal input
rlabel metal2 s 67546 180003 67602 180803 6 io_in[20]
port 78 nsew signal input
rlabel metal2 s 70858 180003 70914 180803 6 io_in[21]
port 79 nsew signal input
rlabel metal2 s 74262 180003 74318 180803 6 io_in[22]
port 80 nsew signal input
rlabel metal2 s 77574 180003 77630 180803 6 io_in[23]
port 81 nsew signal input
rlabel metal2 s 80886 180003 80942 180803 6 io_in[24]
port 82 nsew signal input
rlabel metal2 s 84290 180003 84346 180803 6 io_in[25]
port 83 nsew signal input
rlabel metal2 s 87602 180003 87658 180803 6 io_in[26]
port 84 nsew signal input
rlabel metal2 s 91006 180003 91062 180803 6 io_in[27]
port 85 nsew signal input
rlabel metal2 s 94318 180003 94374 180803 6 io_in[28]
port 86 nsew signal input
rlabel metal2 s 97630 180003 97686 180803 6 io_in[29]
port 87 nsew signal input
rlabel metal2 s 7194 180003 7250 180803 6 io_in[2]
port 88 nsew signal input
rlabel metal2 s 101034 180003 101090 180803 6 io_in[30]
port 89 nsew signal input
rlabel metal2 s 104346 180003 104402 180803 6 io_in[31]
port 90 nsew signal input
rlabel metal2 s 107750 180003 107806 180803 6 io_in[32]
port 91 nsew signal input
rlabel metal2 s 111062 180003 111118 180803 6 io_in[33]
port 92 nsew signal input
rlabel metal2 s 114466 180003 114522 180803 6 io_in[34]
port 93 nsew signal input
rlabel metal2 s 117778 180003 117834 180803 6 io_in[35]
port 94 nsew signal input
rlabel metal2 s 121090 180003 121146 180803 6 io_in[36]
port 95 nsew signal input
rlabel metal2 s 124494 180003 124550 180803 6 io_in[37]
port 96 nsew signal input
rlabel metal2 s 10598 180003 10654 180803 6 io_in[3]
port 97 nsew signal input
rlabel metal2 s 13910 180003 13966 180803 6 io_in[4]
port 98 nsew signal input
rlabel metal2 s 17314 180003 17370 180803 6 io_in[5]
port 99 nsew signal input
rlabel metal2 s 20626 180003 20682 180803 6 io_in[6]
port 100 nsew signal input
rlabel metal2 s 23938 180003 23994 180803 6 io_in[7]
port 101 nsew signal input
rlabel metal2 s 27342 180003 27398 180803 6 io_in[8]
port 102 nsew signal input
rlabel metal2 s 30654 180003 30710 180803 6 io_in[9]
port 103 nsew signal input
rlabel metal2 s 1674 180003 1730 180803 6 io_oeb[0]
port 104 nsew signal output
rlabel metal2 s 35162 180003 35218 180803 6 io_oeb[10]
port 105 nsew signal output
rlabel metal2 s 38474 180003 38530 180803 6 io_oeb[11]
port 106 nsew signal output
rlabel metal2 s 41878 180003 41934 180803 6 io_oeb[12]
port 107 nsew signal output
rlabel metal2 s 45190 180003 45246 180803 6 io_oeb[13]
port 108 nsew signal output
rlabel metal2 s 48502 180003 48558 180803 6 io_oeb[14]
port 109 nsew signal output
rlabel metal2 s 51906 180003 51962 180803 6 io_oeb[15]
port 110 nsew signal output
rlabel metal2 s 55218 180003 55274 180803 6 io_oeb[16]
port 111 nsew signal output
rlabel metal2 s 58622 180003 58678 180803 6 io_oeb[17]
port 112 nsew signal output
rlabel metal2 s 61934 180003 61990 180803 6 io_oeb[18]
port 113 nsew signal output
rlabel metal2 s 65246 180003 65302 180803 6 io_oeb[19]
port 114 nsew signal output
rlabel metal2 s 4986 180003 5042 180803 6 io_oeb[1]
port 115 nsew signal output
rlabel metal2 s 68650 180003 68706 180803 6 io_oeb[20]
port 116 nsew signal output
rlabel metal2 s 71962 180003 72018 180803 6 io_oeb[21]
port 117 nsew signal output
rlabel metal2 s 75366 180003 75422 180803 6 io_oeb[22]
port 118 nsew signal output
rlabel metal2 s 78678 180003 78734 180803 6 io_oeb[23]
port 119 nsew signal output
rlabel metal2 s 82082 180003 82138 180803 6 io_oeb[24]
port 120 nsew signal output
rlabel metal2 s 85394 180003 85450 180803 6 io_oeb[25]
port 121 nsew signal output
rlabel metal2 s 88706 180003 88762 180803 6 io_oeb[26]
port 122 nsew signal output
rlabel metal2 s 92110 180003 92166 180803 6 io_oeb[27]
port 123 nsew signal output
rlabel metal2 s 95422 180003 95478 180803 6 io_oeb[28]
port 124 nsew signal output
rlabel metal2 s 98826 180003 98882 180803 6 io_oeb[29]
port 125 nsew signal output
rlabel metal2 s 8298 180003 8354 180803 6 io_oeb[2]
port 126 nsew signal output
rlabel metal2 s 102138 180003 102194 180803 6 io_oeb[30]
port 127 nsew signal output
rlabel metal2 s 105450 180003 105506 180803 6 io_oeb[31]
port 128 nsew signal output
rlabel metal2 s 108854 180003 108910 180803 6 io_oeb[32]
port 129 nsew signal output
rlabel metal2 s 112166 180003 112222 180803 6 io_oeb[33]
port 130 nsew signal output
rlabel metal2 s 115570 180003 115626 180803 6 io_oeb[34]
port 131 nsew signal output
rlabel metal2 s 118882 180003 118938 180803 6 io_oeb[35]
port 132 nsew signal output
rlabel metal2 s 122194 180003 122250 180803 6 io_oeb[36]
port 133 nsew signal output
rlabel metal2 s 125598 180003 125654 180803 6 io_oeb[37]
port 134 nsew signal output
rlabel metal2 s 11702 180003 11758 180803 6 io_oeb[3]
port 135 nsew signal output
rlabel metal2 s 15014 180003 15070 180803 6 io_oeb[4]
port 136 nsew signal output
rlabel metal2 s 18418 180003 18474 180803 6 io_oeb[5]
port 137 nsew signal output
rlabel metal2 s 21730 180003 21786 180803 6 io_oeb[6]
port 138 nsew signal output
rlabel metal2 s 25134 180003 25190 180803 6 io_oeb[7]
port 139 nsew signal output
rlabel metal2 s 28446 180003 28502 180803 6 io_oeb[8]
port 140 nsew signal output
rlabel metal2 s 31758 180003 31814 180803 6 io_oeb[9]
port 141 nsew signal output
rlabel metal2 s 2778 180003 2834 180803 6 io_out[0]
port 142 nsew signal output
rlabel metal2 s 36266 180003 36322 180803 6 io_out[10]
port 143 nsew signal output
rlabel metal2 s 39578 180003 39634 180803 6 io_out[11]
port 144 nsew signal output
rlabel metal2 s 42982 180003 43038 180803 6 io_out[12]
port 145 nsew signal output
rlabel metal2 s 46294 180003 46350 180803 6 io_out[13]
port 146 nsew signal output
rlabel metal2 s 49698 180003 49754 180803 6 io_out[14]
port 147 nsew signal output
rlabel metal2 s 53010 180003 53066 180803 6 io_out[15]
port 148 nsew signal output
rlabel metal2 s 56322 180003 56378 180803 6 io_out[16]
port 149 nsew signal output
rlabel metal2 s 59726 180003 59782 180803 6 io_out[17]
port 150 nsew signal output
rlabel metal2 s 63038 180003 63094 180803 6 io_out[18]
port 151 nsew signal output
rlabel metal2 s 66442 180003 66498 180803 6 io_out[19]
port 152 nsew signal output
rlabel metal2 s 6090 180003 6146 180803 6 io_out[1]
port 153 nsew signal output
rlabel metal2 s 69754 180003 69810 180803 6 io_out[20]
port 154 nsew signal output
rlabel metal2 s 73066 180003 73122 180803 6 io_out[21]
port 155 nsew signal output
rlabel metal2 s 76470 180003 76526 180803 6 io_out[22]
port 156 nsew signal output
rlabel metal2 s 79782 180003 79838 180803 6 io_out[23]
port 157 nsew signal output
rlabel metal2 s 83186 180003 83242 180803 6 io_out[24]
port 158 nsew signal output
rlabel metal2 s 86498 180003 86554 180803 6 io_out[25]
port 159 nsew signal output
rlabel metal2 s 89902 180003 89958 180803 6 io_out[26]
port 160 nsew signal output
rlabel metal2 s 93214 180003 93270 180803 6 io_out[27]
port 161 nsew signal output
rlabel metal2 s 96526 180003 96582 180803 6 io_out[28]
port 162 nsew signal output
rlabel metal2 s 99930 180003 99986 180803 6 io_out[29]
port 163 nsew signal output
rlabel metal2 s 9494 180003 9550 180803 6 io_out[2]
port 164 nsew signal output
rlabel metal2 s 103242 180003 103298 180803 6 io_out[30]
port 165 nsew signal output
rlabel metal2 s 106646 180003 106702 180803 6 io_out[31]
port 166 nsew signal output
rlabel metal2 s 109958 180003 110014 180803 6 io_out[32]
port 167 nsew signal output
rlabel metal2 s 113270 180003 113326 180803 6 io_out[33]
port 168 nsew signal output
rlabel metal2 s 116674 180003 116730 180803 6 io_out[34]
port 169 nsew signal output
rlabel metal2 s 119986 180003 120042 180803 6 io_out[35]
port 170 nsew signal output
rlabel metal2 s 123390 180003 123446 180803 6 io_out[36]
port 171 nsew signal output
rlabel metal2 s 126702 180003 126758 180803 6 io_out[37]
port 172 nsew signal output
rlabel metal2 s 12806 180003 12862 180803 6 io_out[3]
port 173 nsew signal output
rlabel metal2 s 16118 180003 16174 180803 6 io_out[4]
port 174 nsew signal output
rlabel metal2 s 19522 180003 19578 180803 6 io_out[5]
port 175 nsew signal output
rlabel metal2 s 22834 180003 22890 180803 6 io_out[6]
port 176 nsew signal output
rlabel metal2 s 26238 180003 26294 180803 6 io_out[7]
port 177 nsew signal output
rlabel metal2 s 29550 180003 29606 180803 6 io_out[8]
port 178 nsew signal output
rlabel metal2 s 32862 180003 32918 180803 6 io_out[9]
port 179 nsew signal output
rlabel metal2 s 136730 0 136786 800 6 irq[0]
port 180 nsew signal output
rlabel metal2 s 138018 0 138074 800 6 irq[1]
port 181 nsew signal output
rlabel metal2 s 139306 0 139362 800 6 irq[2]
port 182 nsew signal output
rlabel metal3 s 177859 1912 178659 2032 6 o_csb0
port 183 nsew signal output
rlabel metal2 s 128910 180003 128966 180803 6 o_csb0_1
port 184 nsew signal output
rlabel metal2 s 131210 180003 131266 180803 6 o_din0[0]
port 185 nsew signal output
rlabel metal3 s 177859 82152 178659 82272 6 o_din0[10]
port 186 nsew signal output
rlabel metal3 s 177859 86232 178659 86352 6 o_din0[11]
port 187 nsew signal output
rlabel metal2 s 159914 0 159970 800 6 o_din0[12]
port 188 nsew signal output
rlabel metal3 s 0 118056 800 118176 6 o_din0[13]
port 189 nsew signal output
rlabel metal3 s 177859 106224 178659 106344 6 o_din0[14]
port 190 nsew signal output
rlabel metal2 s 162490 0 162546 800 6 o_din0[15]
port 191 nsew signal output
rlabel metal3 s 0 127440 800 127560 6 o_din0[16]
port 192 nsew signal output
rlabel metal2 s 166354 0 166410 800 6 o_din0[17]
port 193 nsew signal output
rlabel metal3 s 177859 122408 178659 122528 6 o_din0[18]
port 194 nsew signal output
rlabel metal2 s 159086 180003 159142 180803 6 o_din0[19]
port 195 nsew signal output
rlabel metal3 s 177859 25984 178659 26104 6 o_din0[1]
port 196 nsew signal output
rlabel metal3 s 0 145936 800 146056 6 o_din0[20]
port 197 nsew signal output
rlabel metal3 s 177859 134376 178659 134496 6 o_din0[21]
port 198 nsew signal output
rlabel metal2 s 164698 180003 164754 180803 6 o_din0[22]
port 199 nsew signal output
rlabel metal3 s 0 155184 800 155304 6 o_din0[23]
port 200 nsew signal output
rlabel metal2 s 166906 180003 166962 180803 6 o_din0[24]
port 201 nsew signal output
rlabel metal2 s 174082 0 174138 800 6 o_din0[25]
port 202 nsew signal output
rlabel metal2 s 169114 180003 169170 180803 6 o_din0[26]
port 203 nsew signal output
rlabel metal2 s 172518 180003 172574 180803 6 o_din0[27]
port 204 nsew signal output
rlabel metal3 s 177859 170552 178659 170672 6 o_din0[28]
port 205 nsew signal output
rlabel metal3 s 0 169056 800 169176 6 o_din0[29]
port 206 nsew signal output
rlabel metal3 s 0 25440 800 25560 6 o_din0[2]
port 207 nsew signal output
rlabel metal3 s 0 178304 800 178424 6 o_din0[30]
port 208 nsew signal output
rlabel metal2 s 178038 180003 178094 180803 6 o_din0[31]
port 209 nsew signal output
rlabel metal3 s 0 39312 800 39432 6 o_din0[3]
port 210 nsew signal output
rlabel metal2 s 141238 180003 141294 180803 6 o_din0[4]
port 211 nsew signal output
rlabel metal2 s 149610 0 149666 800 6 o_din0[5]
port 212 nsew signal output
rlabel metal3 s 177859 45976 178659 46096 6 o_din0[6]
port 213 nsew signal output
rlabel metal2 s 144550 180003 144606 180803 6 o_din0[7]
port 214 nsew signal output
rlabel metal2 s 154762 0 154818 800 6 o_din0[8]
port 215 nsew signal output
rlabel metal3 s 177859 78208 178659 78328 6 o_din0[9]
port 216 nsew signal output
rlabel metal3 s 177859 17960 178659 18080 6 o_din0_1[0]
port 217 nsew signal output
rlabel metal3 s 0 104184 800 104304 6 o_din0_1[10]
port 218 nsew signal output
rlabel metal2 s 158626 0 158682 800 6 o_din0_1[11]
port 219 nsew signal output
rlabel metal3 s 177859 94256 178659 94376 6 o_din0_1[12]
port 220 nsew signal output
rlabel metal3 s 177859 98200 178659 98320 6 o_din0_1[13]
port 221 nsew signal output
rlabel metal3 s 177859 102280 178659 102400 6 o_din0_1[14]
port 222 nsew signal output
rlabel metal2 s 153474 180003 153530 180803 6 o_din0_1[15]
port 223 nsew signal output
rlabel metal2 s 163778 0 163834 800 6 o_din0_1[16]
port 224 nsew signal output
rlabel metal2 s 155774 180003 155830 180803 6 o_din0_1[17]
port 225 nsew signal output
rlabel metal3 s 0 132064 800 132184 6 o_din0_1[18]
port 226 nsew signal output
rlabel metal2 s 157982 180003 158038 180803 6 o_din0_1[19]
port 227 nsew signal output
rlabel metal2 s 132314 180003 132370 180803 6 o_din0_1[1]
port 228 nsew signal output
rlabel metal2 s 160190 180003 160246 180803 6 o_din0_1[20]
port 229 nsew signal output
rlabel metal2 s 162398 180003 162454 180803 6 o_din0_1[21]
port 230 nsew signal output
rlabel metal2 s 163594 180003 163650 180803 6 o_din0_1[22]
port 231 nsew signal output
rlabel metal2 s 165802 180003 165858 180803 6 o_din0_1[23]
port 232 nsew signal output
rlabel metal3 s 177859 150424 178659 150544 6 o_din0_1[24]
port 233 nsew signal output
rlabel metal2 s 172794 0 172850 800 6 o_din0_1[25]
port 234 nsew signal output
rlabel metal2 s 168010 180003 168066 180803 6 o_din0_1[26]
port 235 nsew signal output
rlabel metal2 s 171414 180003 171470 180803 6 o_din0_1[27]
port 236 nsew signal output
rlabel metal2 s 174726 180003 174782 180803 6 o_din0_1[28]
port 237 nsew signal output
rlabel metal2 s 176934 180003 176990 180803 6 o_din0_1[29]
port 238 nsew signal output
rlabel metal3 s 0 20816 800 20936 6 o_din0_1[2]
port 239 nsew signal output
rlabel metal3 s 0 173680 800 173800 6 o_din0_1[30]
port 240 nsew signal output
rlabel metal2 s 177946 0 178002 800 6 o_din0_1[31]
port 241 nsew signal output
rlabel metal2 s 139030 180003 139086 180803 6 o_din0_1[3]
port 242 nsew signal output
rlabel metal3 s 0 53184 800 53304 6 o_din0_1[4]
port 243 nsew signal output
rlabel metal3 s 0 71816 800 71936 6 o_din0_1[5]
port 244 nsew signal output
rlabel metal2 s 143446 180003 143502 180803 6 o_din0_1[6]
port 245 nsew signal output
rlabel metal3 s 177859 58080 178659 58200 6 o_din0_1[7]
port 246 nsew signal output
rlabel metal3 s 0 85688 800 85808 6 o_din0_1[8]
port 247 nsew signal output
rlabel metal3 s 0 94936 800 95056 6 o_din0_1[9]
port 248 nsew signal output
rlabel metal3 s 0 6944 800 7064 6 o_waddr0[0]
port 249 nsew signal output
rlabel metal2 s 133418 180003 133474 180803 6 o_waddr0[1]
port 250 nsew signal output
rlabel metal2 s 136730 180003 136786 180803 6 o_waddr0[2]
port 251 nsew signal output
rlabel metal3 s 0 48560 800 48680 6 o_waddr0[3]
port 252 nsew signal output
rlabel metal3 s 0 57808 800 57928 6 o_waddr0[4]
port 253 nsew signal output
rlabel metal2 s 142342 180003 142398 180803 6 o_waddr0[5]
port 254 nsew signal output
rlabel metal2 s 152186 0 152242 800 6 o_waddr0[6]
port 255 nsew signal output
rlabel metal3 s 177859 66104 178659 66224 6 o_waddr0[7]
port 256 nsew signal output
rlabel metal3 s 177859 74128 178659 74248 6 o_waddr0[8]
port 257 nsew signal output
rlabel metal2 s 140594 0 140650 800 6 o_waddr0_1[0]
port 258 nsew signal output
rlabel metal3 s 0 16192 800 16312 6 o_waddr0_1[1]
port 259 nsew signal output
rlabel metal3 s 177859 34008 178659 34128 6 o_waddr0_1[2]
port 260 nsew signal output
rlabel metal3 s 0 43936 800 44056 6 o_waddr0_1[3]
port 261 nsew signal output
rlabel metal2 s 148322 0 148378 800 6 o_waddr0_1[4]
port 262 nsew signal output
rlabel metal3 s 0 76440 800 76560 6 o_waddr0_1[5]
port 263 nsew signal output
rlabel metal3 s 177859 50056 178659 50176 6 o_waddr0_1[6]
port 264 nsew signal output
rlabel metal3 s 177859 62160 178659 62280 6 o_waddr0_1[7]
port 265 nsew signal output
rlabel metal2 s 146850 180003 146906 180803 6 o_waddr0_1[8]
port 266 nsew signal output
rlabel metal3 s 177859 5856 178659 5976 6 o_web0
port 267 nsew signal output
rlabel metal3 s 177859 9936 178659 10056 6 o_web0_1
port 268 nsew signal output
rlabel metal3 s 0 11568 800 11688 6 o_wmask0[0]
port 269 nsew signal output
rlabel metal3 s 177859 29928 178659 30048 6 o_wmask0[1]
port 270 nsew signal output
rlabel metal2 s 137834 180003 137890 180803 6 o_wmask0[2]
port 271 nsew signal output
rlabel metal3 s 177859 37952 178659 38072 6 o_wmask0[3]
port 272 nsew signal output
rlabel metal3 s 177859 21904 178659 22024 6 o_wmask0_1[0]
port 273 nsew signal output
rlabel metal2 s 134522 180003 134578 180803 6 o_wmask0_1[1]
port 274 nsew signal output
rlabel metal3 s 0 30064 800 30184 6 o_wmask0_1[2]
port 275 nsew signal output
rlabel metal2 s 140134 180003 140190 180803 6 o_wmask0_1[3]
port 276 nsew signal output
rlabel metal3 s 0 2320 800 2440 6 rst_i
port 277 nsew signal input
rlabel metal4 s 4208 2128 4528 178480 6 vccd1
port 278 nsew power input
rlabel metal4 s 34928 2128 35248 178480 6 vccd1
port 278 nsew power input
rlabel metal4 s 65648 2128 65968 178480 6 vccd1
port 278 nsew power input
rlabel metal4 s 96368 2128 96688 178480 6 vccd1
port 278 nsew power input
rlabel metal4 s 127088 2128 127408 178480 6 vccd1
port 278 nsew power input
rlabel metal4 s 157808 2128 158128 178480 6 vccd1
port 278 nsew power input
rlabel metal4 s 19568 2128 19888 178480 6 vssd1
port 279 nsew ground input
rlabel metal4 s 50288 2128 50608 178480 6 vssd1
port 279 nsew ground input
rlabel metal4 s 81008 2128 81328 178480 6 vssd1
port 279 nsew ground input
rlabel metal4 s 111728 2128 112048 178480 6 vssd1
port 279 nsew ground input
rlabel metal4 s 142448 2128 142768 178480 6 vssd1
port 279 nsew ground input
rlabel metal4 s 173168 2128 173488 178480 6 vssd1
port 279 nsew ground input
rlabel metal2 s 570 0 626 800 6 wb_clk_i
port 280 nsew signal input
rlabel metal2 s 1766 0 1822 800 6 wb_rst_i
port 281 nsew signal input
rlabel metal2 s 3054 0 3110 800 6 wbs_ack_o
port 282 nsew signal output
rlabel metal2 s 8206 0 8262 800 6 wbs_adr_i[0]
port 283 nsew signal input
rlabel metal2 s 51906 0 51962 800 6 wbs_adr_i[10]
port 284 nsew signal input
rlabel metal2 s 55770 0 55826 800 6 wbs_adr_i[11]
port 285 nsew signal input
rlabel metal2 s 59634 0 59690 800 6 wbs_adr_i[12]
port 286 nsew signal input
rlabel metal2 s 63498 0 63554 800 6 wbs_adr_i[13]
port 287 nsew signal input
rlabel metal2 s 67362 0 67418 800 6 wbs_adr_i[14]
port 288 nsew signal input
rlabel metal2 s 71226 0 71282 800 6 wbs_adr_i[15]
port 289 nsew signal input
rlabel metal2 s 75090 0 75146 800 6 wbs_adr_i[16]
port 290 nsew signal input
rlabel metal2 s 78954 0 79010 800 6 wbs_adr_i[17]
port 291 nsew signal input
rlabel metal2 s 82818 0 82874 800 6 wbs_adr_i[18]
port 292 nsew signal input
rlabel metal2 s 86682 0 86738 800 6 wbs_adr_i[19]
port 293 nsew signal input
rlabel metal2 s 13358 0 13414 800 6 wbs_adr_i[1]
port 294 nsew signal input
rlabel metal2 s 90454 0 90510 800 6 wbs_adr_i[20]
port 295 nsew signal input
rlabel metal2 s 94318 0 94374 800 6 wbs_adr_i[21]
port 296 nsew signal input
rlabel metal2 s 98182 0 98238 800 6 wbs_adr_i[22]
port 297 nsew signal input
rlabel metal2 s 102046 0 102102 800 6 wbs_adr_i[23]
port 298 nsew signal input
rlabel metal2 s 105910 0 105966 800 6 wbs_adr_i[24]
port 299 nsew signal input
rlabel metal2 s 109774 0 109830 800 6 wbs_adr_i[25]
port 300 nsew signal input
rlabel metal2 s 113638 0 113694 800 6 wbs_adr_i[26]
port 301 nsew signal input
rlabel metal2 s 117502 0 117558 800 6 wbs_adr_i[27]
port 302 nsew signal input
rlabel metal2 s 121366 0 121422 800 6 wbs_adr_i[28]
port 303 nsew signal input
rlabel metal2 s 125230 0 125286 800 6 wbs_adr_i[29]
port 304 nsew signal input
rlabel metal2 s 18510 0 18566 800 6 wbs_adr_i[2]
port 305 nsew signal input
rlabel metal2 s 129094 0 129150 800 6 wbs_adr_i[30]
port 306 nsew signal input
rlabel metal2 s 132958 0 133014 800 6 wbs_adr_i[31]
port 307 nsew signal input
rlabel metal2 s 23662 0 23718 800 6 wbs_adr_i[3]
port 308 nsew signal input
rlabel metal2 s 28814 0 28870 800 6 wbs_adr_i[4]
port 309 nsew signal input
rlabel metal2 s 32678 0 32734 800 6 wbs_adr_i[5]
port 310 nsew signal input
rlabel metal2 s 36542 0 36598 800 6 wbs_adr_i[6]
port 311 nsew signal input
rlabel metal2 s 40406 0 40462 800 6 wbs_adr_i[7]
port 312 nsew signal input
rlabel metal2 s 44270 0 44326 800 6 wbs_adr_i[8]
port 313 nsew signal input
rlabel metal2 s 48042 0 48098 800 6 wbs_adr_i[9]
port 314 nsew signal input
rlabel metal2 s 4342 0 4398 800 6 wbs_cyc_i
port 315 nsew signal input
rlabel metal2 s 9494 0 9550 800 6 wbs_dat_i[0]
port 316 nsew signal input
rlabel metal2 s 53194 0 53250 800 6 wbs_dat_i[10]
port 317 nsew signal input
rlabel metal2 s 57058 0 57114 800 6 wbs_dat_i[11]
port 318 nsew signal input
rlabel metal2 s 60922 0 60978 800 6 wbs_dat_i[12]
port 319 nsew signal input
rlabel metal2 s 64786 0 64842 800 6 wbs_dat_i[13]
port 320 nsew signal input
rlabel metal2 s 68650 0 68706 800 6 wbs_dat_i[14]
port 321 nsew signal input
rlabel metal2 s 72514 0 72570 800 6 wbs_dat_i[15]
port 322 nsew signal input
rlabel metal2 s 76378 0 76434 800 6 wbs_dat_i[16]
port 323 nsew signal input
rlabel metal2 s 80242 0 80298 800 6 wbs_dat_i[17]
port 324 nsew signal input
rlabel metal2 s 84106 0 84162 800 6 wbs_dat_i[18]
port 325 nsew signal input
rlabel metal2 s 87970 0 88026 800 6 wbs_dat_i[19]
port 326 nsew signal input
rlabel metal2 s 14646 0 14702 800 6 wbs_dat_i[1]
port 327 nsew signal input
rlabel metal2 s 91742 0 91798 800 6 wbs_dat_i[20]
port 328 nsew signal input
rlabel metal2 s 95606 0 95662 800 6 wbs_dat_i[21]
port 329 nsew signal input
rlabel metal2 s 99470 0 99526 800 6 wbs_dat_i[22]
port 330 nsew signal input
rlabel metal2 s 103334 0 103390 800 6 wbs_dat_i[23]
port 331 nsew signal input
rlabel metal2 s 107198 0 107254 800 6 wbs_dat_i[24]
port 332 nsew signal input
rlabel metal2 s 111062 0 111118 800 6 wbs_dat_i[25]
port 333 nsew signal input
rlabel metal2 s 114926 0 114982 800 6 wbs_dat_i[26]
port 334 nsew signal input
rlabel metal2 s 118790 0 118846 800 6 wbs_dat_i[27]
port 335 nsew signal input
rlabel metal2 s 122654 0 122710 800 6 wbs_dat_i[28]
port 336 nsew signal input
rlabel metal2 s 126518 0 126574 800 6 wbs_dat_i[29]
port 337 nsew signal input
rlabel metal2 s 19798 0 19854 800 6 wbs_dat_i[2]
port 338 nsew signal input
rlabel metal2 s 130382 0 130438 800 6 wbs_dat_i[30]
port 339 nsew signal input
rlabel metal2 s 134246 0 134302 800 6 wbs_dat_i[31]
port 340 nsew signal input
rlabel metal2 s 24950 0 25006 800 6 wbs_dat_i[3]
port 341 nsew signal input
rlabel metal2 s 30102 0 30158 800 6 wbs_dat_i[4]
port 342 nsew signal input
rlabel metal2 s 33966 0 34022 800 6 wbs_dat_i[5]
port 343 nsew signal input
rlabel metal2 s 37830 0 37886 800 6 wbs_dat_i[6]
port 344 nsew signal input
rlabel metal2 s 41694 0 41750 800 6 wbs_dat_i[7]
port 345 nsew signal input
rlabel metal2 s 45466 0 45522 800 6 wbs_dat_i[8]
port 346 nsew signal input
rlabel metal2 s 49330 0 49386 800 6 wbs_dat_i[9]
port 347 nsew signal input
rlabel metal2 s 10782 0 10838 800 6 wbs_dat_o[0]
port 348 nsew signal output
rlabel metal2 s 54482 0 54538 800 6 wbs_dat_o[10]
port 349 nsew signal output
rlabel metal2 s 58346 0 58402 800 6 wbs_dat_o[11]
port 350 nsew signal output
rlabel metal2 s 62210 0 62266 800 6 wbs_dat_o[12]
port 351 nsew signal output
rlabel metal2 s 66074 0 66130 800 6 wbs_dat_o[13]
port 352 nsew signal output
rlabel metal2 s 69938 0 69994 800 6 wbs_dat_o[14]
port 353 nsew signal output
rlabel metal2 s 73802 0 73858 800 6 wbs_dat_o[15]
port 354 nsew signal output
rlabel metal2 s 77666 0 77722 800 6 wbs_dat_o[16]
port 355 nsew signal output
rlabel metal2 s 81530 0 81586 800 6 wbs_dat_o[17]
port 356 nsew signal output
rlabel metal2 s 85394 0 85450 800 6 wbs_dat_o[18]
port 357 nsew signal output
rlabel metal2 s 89258 0 89314 800 6 wbs_dat_o[19]
port 358 nsew signal output
rlabel metal2 s 15934 0 15990 800 6 wbs_dat_o[1]
port 359 nsew signal output
rlabel metal2 s 93030 0 93086 800 6 wbs_dat_o[20]
port 360 nsew signal output
rlabel metal2 s 96894 0 96950 800 6 wbs_dat_o[21]
port 361 nsew signal output
rlabel metal2 s 100758 0 100814 800 6 wbs_dat_o[22]
port 362 nsew signal output
rlabel metal2 s 104622 0 104678 800 6 wbs_dat_o[23]
port 363 nsew signal output
rlabel metal2 s 108486 0 108542 800 6 wbs_dat_o[24]
port 364 nsew signal output
rlabel metal2 s 112350 0 112406 800 6 wbs_dat_o[25]
port 365 nsew signal output
rlabel metal2 s 116214 0 116270 800 6 wbs_dat_o[26]
port 366 nsew signal output
rlabel metal2 s 120078 0 120134 800 6 wbs_dat_o[27]
port 367 nsew signal output
rlabel metal2 s 123942 0 123998 800 6 wbs_dat_o[28]
port 368 nsew signal output
rlabel metal2 s 127806 0 127862 800 6 wbs_dat_o[29]
port 369 nsew signal output
rlabel metal2 s 21086 0 21142 800 6 wbs_dat_o[2]
port 370 nsew signal output
rlabel metal2 s 131670 0 131726 800 6 wbs_dat_o[30]
port 371 nsew signal output
rlabel metal2 s 135442 0 135498 800 6 wbs_dat_o[31]
port 372 nsew signal output
rlabel metal2 s 26238 0 26294 800 6 wbs_dat_o[3]
port 373 nsew signal output
rlabel metal2 s 31390 0 31446 800 6 wbs_dat_o[4]
port 374 nsew signal output
rlabel metal2 s 35254 0 35310 800 6 wbs_dat_o[5]
port 375 nsew signal output
rlabel metal2 s 39118 0 39174 800 6 wbs_dat_o[6]
port 376 nsew signal output
rlabel metal2 s 42982 0 43038 800 6 wbs_dat_o[7]
port 377 nsew signal output
rlabel metal2 s 46754 0 46810 800 6 wbs_dat_o[8]
port 378 nsew signal output
rlabel metal2 s 50618 0 50674 800 6 wbs_dat_o[9]
port 379 nsew signal output
rlabel metal2 s 12070 0 12126 800 6 wbs_sel_i[0]
port 380 nsew signal input
rlabel metal2 s 17222 0 17278 800 6 wbs_sel_i[1]
port 381 nsew signal input
rlabel metal2 s 22374 0 22430 800 6 wbs_sel_i[2]
port 382 nsew signal input
rlabel metal2 s 27526 0 27582 800 6 wbs_sel_i[3]
port 383 nsew signal input
rlabel metal2 s 5630 0 5686 800 6 wbs_stb_i
port 384 nsew signal input
rlabel metal2 s 6918 0 6974 800 6 wbs_we_i
port 385 nsew signal input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 178659 180803
string LEFview TRUE
string GDS_FILE /project/openlane/user_proj/runs/user_proj/results/magic/user_proj.gds
string GDS_END 81877708
string GDS_START 1439632
<< end >>

