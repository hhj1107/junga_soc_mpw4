* NGSPICE file created from user_proj.ext - technology: sky130A

.subckt user_proj clk_i i_dout0[0] i_dout0[10] i_dout0[11] i_dout0[12] i_dout0[13]
+ i_dout0[14] i_dout0[15] i_dout0[16] i_dout0[17] i_dout0[18] i_dout0[19] i_dout0[1]
+ i_dout0[20] i_dout0[21] i_dout0[22] i_dout0[23] i_dout0[24] i_dout0[25] i_dout0[26]
+ i_dout0[27] i_dout0[28] i_dout0[29] i_dout0[2] i_dout0[30] i_dout0[31] i_dout0[3]
+ i_dout0[4] i_dout0[5] i_dout0[6] i_dout0[7] i_dout0[8] i_dout0[9] i_dout0_1[0] i_dout0_1[10]
+ i_dout0_1[11] i_dout0_1[12] i_dout0_1[13] i_dout0_1[14] i_dout0_1[15] i_dout0_1[16]
+ i_dout0_1[17] i_dout0_1[18] i_dout0_1[19] i_dout0_1[1] i_dout0_1[20] i_dout0_1[21]
+ i_dout0_1[22] i_dout0_1[23] i_dout0_1[24] i_dout0_1[25] i_dout0_1[26] i_dout0_1[27]
+ i_dout0_1[28] i_dout0_1[29] i_dout0_1[2] i_dout0_1[30] i_dout0_1[31] i_dout0_1[3]
+ i_dout0_1[4] i_dout0_1[5] i_dout0_1[6] i_dout0_1[7] i_dout0_1[8] i_dout0_1[9] io_in[0]
+ io_in[10] io_in[11] io_in[12] io_in[13] io_in[14] io_in[15] io_in[16] io_in[17]
+ io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22] io_in[23] io_in[24] io_in[25]
+ io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30] io_in[31] io_in[32] io_in[33]
+ io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7]
+ io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14]
+ io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21]
+ io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27] io_oeb[28] io_oeb[29]
+ io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34] io_oeb[35] io_oeb[36]
+ io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9]
+ io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15] io_out[16]
+ io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22] io_out[23]
+ io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29] io_out[2] io_out[30]
+ io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36] io_out[37] io_out[3]
+ io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9] irq[0] irq[1] irq[2]
+ o_csb0 o_csb0_1 o_din0[0] o_din0[10] o_din0[11] o_din0[12] o_din0[13] o_din0[14]
+ o_din0[15] o_din0[16] o_din0[17] o_din0[18] o_din0[19] o_din0[1] o_din0[20] o_din0[21]
+ o_din0[22] o_din0[23] o_din0[24] o_din0[25] o_din0[26] o_din0[27] o_din0[28] o_din0[29]
+ o_din0[2] o_din0[30] o_din0[31] o_din0[3] o_din0[4] o_din0[5] o_din0[6] o_din0[7]
+ o_din0[8] o_din0[9] o_din0_1[0] o_din0_1[10] o_din0_1[11] o_din0_1[12] o_din0_1[13]
+ o_din0_1[14] o_din0_1[15] o_din0_1[16] o_din0_1[17] o_din0_1[18] o_din0_1[19] o_din0_1[1]
+ o_din0_1[20] o_din0_1[21] o_din0_1[22] o_din0_1[23] o_din0_1[24] o_din0_1[25] o_din0_1[26]
+ o_din0_1[27] o_din0_1[28] o_din0_1[29] o_din0_1[2] o_din0_1[30] o_din0_1[31] o_din0_1[3]
+ o_din0_1[4] o_din0_1[5] o_din0_1[6] o_din0_1[7] o_din0_1[8] o_din0_1[9] o_waddr0[0]
+ o_waddr0[1] o_waddr0[2] o_waddr0[3] o_waddr0[4] o_waddr0[5] o_waddr0[6] o_waddr0[7]
+ o_waddr0[8] o_waddr0_1[0] o_waddr0_1[1] o_waddr0_1[2] o_waddr0_1[3] o_waddr0_1[4]
+ o_waddr0_1[5] o_waddr0_1[6] o_waddr0_1[7] o_waddr0_1[8] o_web0 o_web0_1 o_wmask0[0]
+ o_wmask0[1] o_wmask0[2] o_wmask0[3] o_wmask0_1[0] o_wmask0_1[1] o_wmask0_1[2] o_wmask0_1[3]
+ rst_i vccd1 vssd1 wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11]
+ wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17]
+ wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22]
+ wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28]
+ wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4]
+ wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0]
+ wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15]
+ wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20]
+ wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26]
+ wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31]
+ wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9]
+ wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14]
+ wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1]
+ wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25]
+ wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30]
+ wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8]
+ wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
.ends

