magic
tech sky130A
magscale 1 2
timestamp 1639355506
<< obsli1 >>
rect 1104 2159 558808 697425
<< obsm1 >>
rect 566 1640 559438 697456
<< metal2 >>
rect 2410 699200 2466 700000
rect 7286 699200 7342 700000
rect 12162 699200 12218 700000
rect 17130 699200 17186 700000
rect 22006 699200 22062 700000
rect 26882 699200 26938 700000
rect 31850 699200 31906 700000
rect 36726 699200 36782 700000
rect 41694 699200 41750 700000
rect 46570 699200 46626 700000
rect 51446 699200 51502 700000
rect 56414 699200 56470 700000
rect 61290 699200 61346 700000
rect 66258 699200 66314 700000
rect 71134 699200 71190 700000
rect 76010 699200 76066 700000
rect 80978 699200 81034 700000
rect 85854 699200 85910 700000
rect 90822 699200 90878 700000
rect 95698 699200 95754 700000
rect 100574 699200 100630 700000
rect 105542 699200 105598 700000
rect 110418 699200 110474 700000
rect 115386 699200 115442 700000
rect 120262 699200 120318 700000
rect 125138 699200 125194 700000
rect 130106 699200 130162 700000
rect 134982 699200 135038 700000
rect 139950 699200 140006 700000
rect 144826 699200 144882 700000
rect 149702 699200 149758 700000
rect 154670 699200 154726 700000
rect 159546 699200 159602 700000
rect 164514 699200 164570 700000
rect 169390 699200 169446 700000
rect 174266 699200 174322 700000
rect 179234 699200 179290 700000
rect 184110 699200 184166 700000
rect 189078 699200 189134 700000
rect 193954 699200 194010 700000
rect 198830 699200 198886 700000
rect 203798 699200 203854 700000
rect 208674 699200 208730 700000
rect 213550 699200 213606 700000
rect 218518 699200 218574 700000
rect 223394 699200 223450 700000
rect 228362 699200 228418 700000
rect 233238 699200 233294 700000
rect 238114 699200 238170 700000
rect 243082 699200 243138 700000
rect 247958 699200 248014 700000
rect 252926 699200 252982 700000
rect 257802 699200 257858 700000
rect 262678 699200 262734 700000
rect 267646 699200 267702 700000
rect 272522 699200 272578 700000
rect 277490 699200 277546 700000
rect 282366 699200 282422 700000
rect 287242 699200 287298 700000
rect 292210 699200 292266 700000
rect 297086 699200 297142 700000
rect 302054 699200 302110 700000
rect 306930 699200 306986 700000
rect 311806 699200 311862 700000
rect 316774 699200 316830 700000
rect 321650 699200 321706 700000
rect 326618 699200 326674 700000
rect 331494 699200 331550 700000
rect 336370 699200 336426 700000
rect 341338 699200 341394 700000
rect 346214 699200 346270 700000
rect 351182 699200 351238 700000
rect 356058 699200 356114 700000
rect 360934 699200 360990 700000
rect 365902 699200 365958 700000
rect 370778 699200 370834 700000
rect 375746 699200 375802 700000
rect 380622 699200 380678 700000
rect 385498 699200 385554 700000
rect 390466 699200 390522 700000
rect 395342 699200 395398 700000
rect 400218 699200 400274 700000
rect 405186 699200 405242 700000
rect 410062 699200 410118 700000
rect 415030 699200 415086 700000
rect 419906 699200 419962 700000
rect 424782 699200 424838 700000
rect 429750 699200 429806 700000
rect 434626 699200 434682 700000
rect 439594 699200 439650 700000
rect 444470 699200 444526 700000
rect 449346 699200 449402 700000
rect 454314 699200 454370 700000
rect 459190 699200 459246 700000
rect 464158 699200 464214 700000
rect 469034 699200 469090 700000
rect 473910 699200 473966 700000
rect 478878 699200 478934 700000
rect 483754 699200 483810 700000
rect 488722 699200 488778 700000
rect 493598 699200 493654 700000
rect 498474 699200 498530 700000
rect 503442 699200 503498 700000
rect 508318 699200 508374 700000
rect 513286 699200 513342 700000
rect 518162 699200 518218 700000
rect 523038 699200 523094 700000
rect 528006 699200 528062 700000
rect 532882 699200 532938 700000
rect 537850 699200 537906 700000
rect 542726 699200 542782 700000
rect 547602 699200 547658 700000
rect 552570 699200 552626 700000
rect 557446 699200 557502 700000
rect 570 0 626 800
rect 1674 0 1730 800
rect 2778 0 2834 800
rect 3974 0 4030 800
rect 5078 0 5134 800
rect 6182 0 6238 800
rect 7378 0 7434 800
rect 8482 0 8538 800
rect 9586 0 9642 800
rect 10782 0 10838 800
rect 11886 0 11942 800
rect 12990 0 13046 800
rect 14186 0 14242 800
rect 15290 0 15346 800
rect 16394 0 16450 800
rect 17590 0 17646 800
rect 18694 0 18750 800
rect 19798 0 19854 800
rect 20994 0 21050 800
rect 22098 0 22154 800
rect 23202 0 23258 800
rect 24398 0 24454 800
rect 25502 0 25558 800
rect 26606 0 26662 800
rect 27802 0 27858 800
rect 28906 0 28962 800
rect 30102 0 30158 800
rect 31206 0 31262 800
rect 32310 0 32366 800
rect 33506 0 33562 800
rect 34610 0 34666 800
rect 35714 0 35770 800
rect 36910 0 36966 800
rect 38014 0 38070 800
rect 39118 0 39174 800
rect 40314 0 40370 800
rect 41418 0 41474 800
rect 42522 0 42578 800
rect 43718 0 43774 800
rect 44822 0 44878 800
rect 45926 0 45982 800
rect 47122 0 47178 800
rect 48226 0 48282 800
rect 49330 0 49386 800
rect 50526 0 50582 800
rect 51630 0 51686 800
rect 52734 0 52790 800
rect 53930 0 53986 800
rect 55034 0 55090 800
rect 56138 0 56194 800
rect 57334 0 57390 800
rect 58438 0 58494 800
rect 59634 0 59690 800
rect 60738 0 60794 800
rect 61842 0 61898 800
rect 63038 0 63094 800
rect 64142 0 64198 800
rect 65246 0 65302 800
rect 66442 0 66498 800
rect 67546 0 67602 800
rect 68650 0 68706 800
rect 69846 0 69902 800
rect 70950 0 71006 800
rect 72054 0 72110 800
rect 73250 0 73306 800
rect 74354 0 74410 800
rect 75458 0 75514 800
rect 76654 0 76710 800
rect 77758 0 77814 800
rect 78862 0 78918 800
rect 80058 0 80114 800
rect 81162 0 81218 800
rect 82266 0 82322 800
rect 83462 0 83518 800
rect 84566 0 84622 800
rect 85762 0 85818 800
rect 86866 0 86922 800
rect 87970 0 88026 800
rect 89166 0 89222 800
rect 90270 0 90326 800
rect 91374 0 91430 800
rect 92570 0 92626 800
rect 93674 0 93730 800
rect 94778 0 94834 800
rect 95974 0 96030 800
rect 97078 0 97134 800
rect 98182 0 98238 800
rect 99378 0 99434 800
rect 100482 0 100538 800
rect 101586 0 101642 800
rect 102782 0 102838 800
rect 103886 0 103942 800
rect 104990 0 105046 800
rect 106186 0 106242 800
rect 107290 0 107346 800
rect 108394 0 108450 800
rect 109590 0 109646 800
rect 110694 0 110750 800
rect 111798 0 111854 800
rect 112994 0 113050 800
rect 114098 0 114154 800
rect 115294 0 115350 800
rect 116398 0 116454 800
rect 117502 0 117558 800
rect 118698 0 118754 800
rect 119802 0 119858 800
rect 120906 0 120962 800
rect 122102 0 122158 800
rect 123206 0 123262 800
rect 124310 0 124366 800
rect 125506 0 125562 800
rect 126610 0 126666 800
rect 127714 0 127770 800
rect 128910 0 128966 800
rect 130014 0 130070 800
rect 131118 0 131174 800
rect 132314 0 132370 800
rect 133418 0 133474 800
rect 134522 0 134578 800
rect 135718 0 135774 800
rect 136822 0 136878 800
rect 137926 0 137982 800
rect 139122 0 139178 800
rect 140226 0 140282 800
rect 141422 0 141478 800
rect 142526 0 142582 800
rect 143630 0 143686 800
rect 144826 0 144882 800
rect 145930 0 145986 800
rect 147034 0 147090 800
rect 148230 0 148286 800
rect 149334 0 149390 800
rect 150438 0 150494 800
rect 151634 0 151690 800
rect 152738 0 152794 800
rect 153842 0 153898 800
rect 155038 0 155094 800
rect 156142 0 156198 800
rect 157246 0 157302 800
rect 158442 0 158498 800
rect 159546 0 159602 800
rect 160650 0 160706 800
rect 161846 0 161902 800
rect 162950 0 163006 800
rect 164054 0 164110 800
rect 165250 0 165306 800
rect 166354 0 166410 800
rect 167458 0 167514 800
rect 168654 0 168710 800
rect 169758 0 169814 800
rect 170954 0 171010 800
rect 172058 0 172114 800
rect 173162 0 173218 800
rect 174358 0 174414 800
rect 175462 0 175518 800
rect 176566 0 176622 800
rect 177762 0 177818 800
rect 178866 0 178922 800
rect 179970 0 180026 800
rect 181166 0 181222 800
rect 182270 0 182326 800
rect 183374 0 183430 800
rect 184570 0 184626 800
rect 185674 0 185730 800
rect 186778 0 186834 800
rect 187974 0 188030 800
rect 189078 0 189134 800
rect 190182 0 190238 800
rect 191378 0 191434 800
rect 192482 0 192538 800
rect 193586 0 193642 800
rect 194782 0 194838 800
rect 195886 0 195942 800
rect 197082 0 197138 800
rect 198186 0 198242 800
rect 199290 0 199346 800
rect 200486 0 200542 800
rect 201590 0 201646 800
rect 202694 0 202750 800
rect 203890 0 203946 800
rect 204994 0 205050 800
rect 206098 0 206154 800
rect 207294 0 207350 800
rect 208398 0 208454 800
rect 209502 0 209558 800
rect 210698 0 210754 800
rect 211802 0 211858 800
rect 212906 0 212962 800
rect 214102 0 214158 800
rect 215206 0 215262 800
rect 216310 0 216366 800
rect 217506 0 217562 800
rect 218610 0 218666 800
rect 219714 0 219770 800
rect 220910 0 220966 800
rect 222014 0 222070 800
rect 223118 0 223174 800
rect 224314 0 224370 800
rect 225418 0 225474 800
rect 226614 0 226670 800
rect 227718 0 227774 800
rect 228822 0 228878 800
rect 230018 0 230074 800
rect 231122 0 231178 800
rect 232226 0 232282 800
rect 233422 0 233478 800
rect 234526 0 234582 800
rect 235630 0 235686 800
rect 236826 0 236882 800
rect 237930 0 237986 800
rect 239034 0 239090 800
rect 240230 0 240286 800
rect 241334 0 241390 800
rect 242438 0 242494 800
rect 243634 0 243690 800
rect 244738 0 244794 800
rect 245842 0 245898 800
rect 247038 0 247094 800
rect 248142 0 248198 800
rect 249246 0 249302 800
rect 250442 0 250498 800
rect 251546 0 251602 800
rect 252742 0 252798 800
rect 253846 0 253902 800
rect 254950 0 255006 800
rect 256146 0 256202 800
rect 257250 0 257306 800
rect 258354 0 258410 800
rect 259550 0 259606 800
rect 260654 0 260710 800
rect 261758 0 261814 800
rect 262954 0 263010 800
rect 264058 0 264114 800
rect 265162 0 265218 800
rect 266358 0 266414 800
rect 267462 0 267518 800
rect 268566 0 268622 800
rect 269762 0 269818 800
rect 270866 0 270922 800
rect 271970 0 272026 800
rect 273166 0 273222 800
rect 274270 0 274326 800
rect 275374 0 275430 800
rect 276570 0 276626 800
rect 277674 0 277730 800
rect 278778 0 278834 800
rect 279974 0 280030 800
rect 281078 0 281134 800
rect 282274 0 282330 800
rect 283378 0 283434 800
rect 284482 0 284538 800
rect 285678 0 285734 800
rect 286782 0 286838 800
rect 287886 0 287942 800
rect 289082 0 289138 800
rect 290186 0 290242 800
rect 291290 0 291346 800
rect 292486 0 292542 800
rect 293590 0 293646 800
rect 294694 0 294750 800
rect 295890 0 295946 800
rect 296994 0 297050 800
rect 298098 0 298154 800
rect 299294 0 299350 800
rect 300398 0 300454 800
rect 301502 0 301558 800
rect 302698 0 302754 800
rect 303802 0 303858 800
rect 304906 0 304962 800
rect 306102 0 306158 800
rect 307206 0 307262 800
rect 308310 0 308366 800
rect 309506 0 309562 800
rect 310610 0 310666 800
rect 311806 0 311862 800
rect 312910 0 312966 800
rect 314014 0 314070 800
rect 315210 0 315266 800
rect 316314 0 316370 800
rect 317418 0 317474 800
rect 318614 0 318670 800
rect 319718 0 319774 800
rect 320822 0 320878 800
rect 322018 0 322074 800
rect 323122 0 323178 800
rect 324226 0 324282 800
rect 325422 0 325478 800
rect 326526 0 326582 800
rect 327630 0 327686 800
rect 328826 0 328882 800
rect 329930 0 329986 800
rect 331034 0 331090 800
rect 332230 0 332286 800
rect 333334 0 333390 800
rect 334438 0 334494 800
rect 335634 0 335690 800
rect 336738 0 336794 800
rect 337934 0 337990 800
rect 339038 0 339094 800
rect 340142 0 340198 800
rect 341338 0 341394 800
rect 342442 0 342498 800
rect 343546 0 343602 800
rect 344742 0 344798 800
rect 345846 0 345902 800
rect 346950 0 347006 800
rect 348146 0 348202 800
rect 349250 0 349306 800
rect 350354 0 350410 800
rect 351550 0 351606 800
rect 352654 0 352710 800
rect 353758 0 353814 800
rect 354954 0 355010 800
rect 356058 0 356114 800
rect 357162 0 357218 800
rect 358358 0 358414 800
rect 359462 0 359518 800
rect 360566 0 360622 800
rect 361762 0 361818 800
rect 362866 0 362922 800
rect 363970 0 364026 800
rect 365166 0 365222 800
rect 366270 0 366326 800
rect 367466 0 367522 800
rect 368570 0 368626 800
rect 369674 0 369730 800
rect 370870 0 370926 800
rect 371974 0 372030 800
rect 373078 0 373134 800
rect 374274 0 374330 800
rect 375378 0 375434 800
rect 376482 0 376538 800
rect 377678 0 377734 800
rect 378782 0 378838 800
rect 379886 0 379942 800
rect 381082 0 381138 800
rect 382186 0 382242 800
rect 383290 0 383346 800
rect 384486 0 384542 800
rect 385590 0 385646 800
rect 386694 0 386750 800
rect 387890 0 387946 800
rect 388994 0 389050 800
rect 390098 0 390154 800
rect 391294 0 391350 800
rect 392398 0 392454 800
rect 393594 0 393650 800
rect 394698 0 394754 800
rect 395802 0 395858 800
rect 396998 0 397054 800
rect 398102 0 398158 800
rect 399206 0 399262 800
rect 400402 0 400458 800
rect 401506 0 401562 800
rect 402610 0 402666 800
rect 403806 0 403862 800
rect 404910 0 404966 800
rect 406014 0 406070 800
rect 407210 0 407266 800
rect 408314 0 408370 800
rect 409418 0 409474 800
rect 410614 0 410670 800
rect 411718 0 411774 800
rect 412822 0 412878 800
rect 414018 0 414074 800
rect 415122 0 415178 800
rect 416226 0 416282 800
rect 417422 0 417478 800
rect 418526 0 418582 800
rect 419630 0 419686 800
rect 420826 0 420882 800
rect 421930 0 421986 800
rect 423126 0 423182 800
rect 424230 0 424286 800
rect 425334 0 425390 800
rect 426530 0 426586 800
rect 427634 0 427690 800
rect 428738 0 428794 800
rect 429934 0 429990 800
rect 431038 0 431094 800
rect 432142 0 432198 800
rect 433338 0 433394 800
rect 434442 0 434498 800
rect 435546 0 435602 800
rect 436742 0 436798 800
rect 437846 0 437902 800
rect 438950 0 439006 800
rect 440146 0 440202 800
rect 441250 0 441306 800
rect 442354 0 442410 800
rect 443550 0 443606 800
rect 444654 0 444710 800
rect 445758 0 445814 800
rect 446954 0 447010 800
rect 448058 0 448114 800
rect 449254 0 449310 800
rect 450358 0 450414 800
rect 451462 0 451518 800
rect 452658 0 452714 800
rect 453762 0 453818 800
rect 454866 0 454922 800
rect 456062 0 456118 800
rect 457166 0 457222 800
rect 458270 0 458326 800
rect 459466 0 459522 800
rect 460570 0 460626 800
rect 461674 0 461730 800
rect 462870 0 462926 800
rect 463974 0 464030 800
rect 465078 0 465134 800
rect 466274 0 466330 800
rect 467378 0 467434 800
rect 468482 0 468538 800
rect 469678 0 469734 800
rect 470782 0 470838 800
rect 471886 0 471942 800
rect 473082 0 473138 800
rect 474186 0 474242 800
rect 475290 0 475346 800
rect 476486 0 476542 800
rect 477590 0 477646 800
rect 478786 0 478842 800
rect 479890 0 479946 800
rect 480994 0 481050 800
rect 482190 0 482246 800
rect 483294 0 483350 800
rect 484398 0 484454 800
rect 485594 0 485650 800
rect 486698 0 486754 800
rect 487802 0 487858 800
rect 488998 0 489054 800
rect 490102 0 490158 800
rect 491206 0 491262 800
rect 492402 0 492458 800
rect 493506 0 493562 800
rect 494610 0 494666 800
rect 495806 0 495862 800
rect 496910 0 496966 800
rect 498014 0 498070 800
rect 499210 0 499266 800
rect 500314 0 500370 800
rect 501418 0 501474 800
rect 502614 0 502670 800
rect 503718 0 503774 800
rect 504914 0 504970 800
rect 506018 0 506074 800
rect 507122 0 507178 800
rect 508318 0 508374 800
rect 509422 0 509478 800
rect 510526 0 510582 800
rect 511722 0 511778 800
rect 512826 0 512882 800
rect 513930 0 513986 800
rect 515126 0 515182 800
rect 516230 0 516286 800
rect 517334 0 517390 800
rect 518530 0 518586 800
rect 519634 0 519690 800
rect 520738 0 520794 800
rect 521934 0 521990 800
rect 523038 0 523094 800
rect 524142 0 524198 800
rect 525338 0 525394 800
rect 526442 0 526498 800
rect 527546 0 527602 800
rect 528742 0 528798 800
rect 529846 0 529902 800
rect 530950 0 531006 800
rect 532146 0 532202 800
rect 533250 0 533306 800
rect 534446 0 534502 800
rect 535550 0 535606 800
rect 536654 0 536710 800
rect 537850 0 537906 800
rect 538954 0 539010 800
rect 540058 0 540114 800
rect 541254 0 541310 800
rect 542358 0 542414 800
rect 543462 0 543518 800
rect 544658 0 544714 800
rect 545762 0 545818 800
rect 546866 0 546922 800
rect 548062 0 548118 800
rect 549166 0 549222 800
rect 550270 0 550326 800
rect 551466 0 551522 800
rect 552570 0 552626 800
rect 553674 0 553730 800
rect 554870 0 554926 800
rect 555974 0 556030 800
rect 557078 0 557134 800
rect 558274 0 558330 800
rect 559378 0 559434 800
<< obsm2 >>
rect 572 699144 2354 699258
rect 2522 699144 7230 699258
rect 7398 699144 12106 699258
rect 12274 699144 17074 699258
rect 17242 699144 21950 699258
rect 22118 699144 26826 699258
rect 26994 699144 31794 699258
rect 31962 699144 36670 699258
rect 36838 699144 41638 699258
rect 41806 699144 46514 699258
rect 46682 699144 51390 699258
rect 51558 699144 56358 699258
rect 56526 699144 61234 699258
rect 61402 699144 66202 699258
rect 66370 699144 71078 699258
rect 71246 699144 75954 699258
rect 76122 699144 80922 699258
rect 81090 699144 85798 699258
rect 85966 699144 90766 699258
rect 90934 699144 95642 699258
rect 95810 699144 100518 699258
rect 100686 699144 105486 699258
rect 105654 699144 110362 699258
rect 110530 699144 115330 699258
rect 115498 699144 120206 699258
rect 120374 699144 125082 699258
rect 125250 699144 130050 699258
rect 130218 699144 134926 699258
rect 135094 699144 139894 699258
rect 140062 699144 144770 699258
rect 144938 699144 149646 699258
rect 149814 699144 154614 699258
rect 154782 699144 159490 699258
rect 159658 699144 164458 699258
rect 164626 699144 169334 699258
rect 169502 699144 174210 699258
rect 174378 699144 179178 699258
rect 179346 699144 184054 699258
rect 184222 699144 189022 699258
rect 189190 699144 193898 699258
rect 194066 699144 198774 699258
rect 198942 699144 203742 699258
rect 203910 699144 208618 699258
rect 208786 699144 213494 699258
rect 213662 699144 218462 699258
rect 218630 699144 223338 699258
rect 223506 699144 228306 699258
rect 228474 699144 233182 699258
rect 233350 699144 238058 699258
rect 238226 699144 243026 699258
rect 243194 699144 247902 699258
rect 248070 699144 252870 699258
rect 253038 699144 257746 699258
rect 257914 699144 262622 699258
rect 262790 699144 267590 699258
rect 267758 699144 272466 699258
rect 272634 699144 277434 699258
rect 277602 699144 282310 699258
rect 282478 699144 287186 699258
rect 287354 699144 292154 699258
rect 292322 699144 297030 699258
rect 297198 699144 301998 699258
rect 302166 699144 306874 699258
rect 307042 699144 311750 699258
rect 311918 699144 316718 699258
rect 316886 699144 321594 699258
rect 321762 699144 326562 699258
rect 326730 699144 331438 699258
rect 331606 699144 336314 699258
rect 336482 699144 341282 699258
rect 341450 699144 346158 699258
rect 346326 699144 351126 699258
rect 351294 699144 356002 699258
rect 356170 699144 360878 699258
rect 361046 699144 365846 699258
rect 366014 699144 370722 699258
rect 370890 699144 375690 699258
rect 375858 699144 380566 699258
rect 380734 699144 385442 699258
rect 385610 699144 390410 699258
rect 390578 699144 395286 699258
rect 395454 699144 400162 699258
rect 400330 699144 405130 699258
rect 405298 699144 410006 699258
rect 410174 699144 414974 699258
rect 415142 699144 419850 699258
rect 420018 699144 424726 699258
rect 424894 699144 429694 699258
rect 429862 699144 434570 699258
rect 434738 699144 439538 699258
rect 439706 699144 444414 699258
rect 444582 699144 449290 699258
rect 449458 699144 454258 699258
rect 454426 699144 459134 699258
rect 459302 699144 464102 699258
rect 464270 699144 468978 699258
rect 469146 699144 473854 699258
rect 474022 699144 478822 699258
rect 478990 699144 483698 699258
rect 483866 699144 488666 699258
rect 488834 699144 493542 699258
rect 493710 699144 498418 699258
rect 498586 699144 503386 699258
rect 503554 699144 508262 699258
rect 508430 699144 513230 699258
rect 513398 699144 518106 699258
rect 518274 699144 522982 699258
rect 523150 699144 527950 699258
rect 528118 699144 532826 699258
rect 532994 699144 537794 699258
rect 537962 699144 542670 699258
rect 542838 699144 547546 699258
rect 547714 699144 552514 699258
rect 552682 699144 557390 699258
rect 557558 699144 559432 699258
rect 572 856 559432 699144
rect 682 734 1618 856
rect 1786 734 2722 856
rect 2890 734 3918 856
rect 4086 734 5022 856
rect 5190 734 6126 856
rect 6294 734 7322 856
rect 7490 734 8426 856
rect 8594 734 9530 856
rect 9698 734 10726 856
rect 10894 734 11830 856
rect 11998 734 12934 856
rect 13102 734 14130 856
rect 14298 734 15234 856
rect 15402 734 16338 856
rect 16506 734 17534 856
rect 17702 734 18638 856
rect 18806 734 19742 856
rect 19910 734 20938 856
rect 21106 734 22042 856
rect 22210 734 23146 856
rect 23314 734 24342 856
rect 24510 734 25446 856
rect 25614 734 26550 856
rect 26718 734 27746 856
rect 27914 734 28850 856
rect 29018 734 30046 856
rect 30214 734 31150 856
rect 31318 734 32254 856
rect 32422 734 33450 856
rect 33618 734 34554 856
rect 34722 734 35658 856
rect 35826 734 36854 856
rect 37022 734 37958 856
rect 38126 734 39062 856
rect 39230 734 40258 856
rect 40426 734 41362 856
rect 41530 734 42466 856
rect 42634 734 43662 856
rect 43830 734 44766 856
rect 44934 734 45870 856
rect 46038 734 47066 856
rect 47234 734 48170 856
rect 48338 734 49274 856
rect 49442 734 50470 856
rect 50638 734 51574 856
rect 51742 734 52678 856
rect 52846 734 53874 856
rect 54042 734 54978 856
rect 55146 734 56082 856
rect 56250 734 57278 856
rect 57446 734 58382 856
rect 58550 734 59578 856
rect 59746 734 60682 856
rect 60850 734 61786 856
rect 61954 734 62982 856
rect 63150 734 64086 856
rect 64254 734 65190 856
rect 65358 734 66386 856
rect 66554 734 67490 856
rect 67658 734 68594 856
rect 68762 734 69790 856
rect 69958 734 70894 856
rect 71062 734 71998 856
rect 72166 734 73194 856
rect 73362 734 74298 856
rect 74466 734 75402 856
rect 75570 734 76598 856
rect 76766 734 77702 856
rect 77870 734 78806 856
rect 78974 734 80002 856
rect 80170 734 81106 856
rect 81274 734 82210 856
rect 82378 734 83406 856
rect 83574 734 84510 856
rect 84678 734 85706 856
rect 85874 734 86810 856
rect 86978 734 87914 856
rect 88082 734 89110 856
rect 89278 734 90214 856
rect 90382 734 91318 856
rect 91486 734 92514 856
rect 92682 734 93618 856
rect 93786 734 94722 856
rect 94890 734 95918 856
rect 96086 734 97022 856
rect 97190 734 98126 856
rect 98294 734 99322 856
rect 99490 734 100426 856
rect 100594 734 101530 856
rect 101698 734 102726 856
rect 102894 734 103830 856
rect 103998 734 104934 856
rect 105102 734 106130 856
rect 106298 734 107234 856
rect 107402 734 108338 856
rect 108506 734 109534 856
rect 109702 734 110638 856
rect 110806 734 111742 856
rect 111910 734 112938 856
rect 113106 734 114042 856
rect 114210 734 115238 856
rect 115406 734 116342 856
rect 116510 734 117446 856
rect 117614 734 118642 856
rect 118810 734 119746 856
rect 119914 734 120850 856
rect 121018 734 122046 856
rect 122214 734 123150 856
rect 123318 734 124254 856
rect 124422 734 125450 856
rect 125618 734 126554 856
rect 126722 734 127658 856
rect 127826 734 128854 856
rect 129022 734 129958 856
rect 130126 734 131062 856
rect 131230 734 132258 856
rect 132426 734 133362 856
rect 133530 734 134466 856
rect 134634 734 135662 856
rect 135830 734 136766 856
rect 136934 734 137870 856
rect 138038 734 139066 856
rect 139234 734 140170 856
rect 140338 734 141366 856
rect 141534 734 142470 856
rect 142638 734 143574 856
rect 143742 734 144770 856
rect 144938 734 145874 856
rect 146042 734 146978 856
rect 147146 734 148174 856
rect 148342 734 149278 856
rect 149446 734 150382 856
rect 150550 734 151578 856
rect 151746 734 152682 856
rect 152850 734 153786 856
rect 153954 734 154982 856
rect 155150 734 156086 856
rect 156254 734 157190 856
rect 157358 734 158386 856
rect 158554 734 159490 856
rect 159658 734 160594 856
rect 160762 734 161790 856
rect 161958 734 162894 856
rect 163062 734 163998 856
rect 164166 734 165194 856
rect 165362 734 166298 856
rect 166466 734 167402 856
rect 167570 734 168598 856
rect 168766 734 169702 856
rect 169870 734 170898 856
rect 171066 734 172002 856
rect 172170 734 173106 856
rect 173274 734 174302 856
rect 174470 734 175406 856
rect 175574 734 176510 856
rect 176678 734 177706 856
rect 177874 734 178810 856
rect 178978 734 179914 856
rect 180082 734 181110 856
rect 181278 734 182214 856
rect 182382 734 183318 856
rect 183486 734 184514 856
rect 184682 734 185618 856
rect 185786 734 186722 856
rect 186890 734 187918 856
rect 188086 734 189022 856
rect 189190 734 190126 856
rect 190294 734 191322 856
rect 191490 734 192426 856
rect 192594 734 193530 856
rect 193698 734 194726 856
rect 194894 734 195830 856
rect 195998 734 197026 856
rect 197194 734 198130 856
rect 198298 734 199234 856
rect 199402 734 200430 856
rect 200598 734 201534 856
rect 201702 734 202638 856
rect 202806 734 203834 856
rect 204002 734 204938 856
rect 205106 734 206042 856
rect 206210 734 207238 856
rect 207406 734 208342 856
rect 208510 734 209446 856
rect 209614 734 210642 856
rect 210810 734 211746 856
rect 211914 734 212850 856
rect 213018 734 214046 856
rect 214214 734 215150 856
rect 215318 734 216254 856
rect 216422 734 217450 856
rect 217618 734 218554 856
rect 218722 734 219658 856
rect 219826 734 220854 856
rect 221022 734 221958 856
rect 222126 734 223062 856
rect 223230 734 224258 856
rect 224426 734 225362 856
rect 225530 734 226558 856
rect 226726 734 227662 856
rect 227830 734 228766 856
rect 228934 734 229962 856
rect 230130 734 231066 856
rect 231234 734 232170 856
rect 232338 734 233366 856
rect 233534 734 234470 856
rect 234638 734 235574 856
rect 235742 734 236770 856
rect 236938 734 237874 856
rect 238042 734 238978 856
rect 239146 734 240174 856
rect 240342 734 241278 856
rect 241446 734 242382 856
rect 242550 734 243578 856
rect 243746 734 244682 856
rect 244850 734 245786 856
rect 245954 734 246982 856
rect 247150 734 248086 856
rect 248254 734 249190 856
rect 249358 734 250386 856
rect 250554 734 251490 856
rect 251658 734 252686 856
rect 252854 734 253790 856
rect 253958 734 254894 856
rect 255062 734 256090 856
rect 256258 734 257194 856
rect 257362 734 258298 856
rect 258466 734 259494 856
rect 259662 734 260598 856
rect 260766 734 261702 856
rect 261870 734 262898 856
rect 263066 734 264002 856
rect 264170 734 265106 856
rect 265274 734 266302 856
rect 266470 734 267406 856
rect 267574 734 268510 856
rect 268678 734 269706 856
rect 269874 734 270810 856
rect 270978 734 271914 856
rect 272082 734 273110 856
rect 273278 734 274214 856
rect 274382 734 275318 856
rect 275486 734 276514 856
rect 276682 734 277618 856
rect 277786 734 278722 856
rect 278890 734 279918 856
rect 280086 734 281022 856
rect 281190 734 282218 856
rect 282386 734 283322 856
rect 283490 734 284426 856
rect 284594 734 285622 856
rect 285790 734 286726 856
rect 286894 734 287830 856
rect 287998 734 289026 856
rect 289194 734 290130 856
rect 290298 734 291234 856
rect 291402 734 292430 856
rect 292598 734 293534 856
rect 293702 734 294638 856
rect 294806 734 295834 856
rect 296002 734 296938 856
rect 297106 734 298042 856
rect 298210 734 299238 856
rect 299406 734 300342 856
rect 300510 734 301446 856
rect 301614 734 302642 856
rect 302810 734 303746 856
rect 303914 734 304850 856
rect 305018 734 306046 856
rect 306214 734 307150 856
rect 307318 734 308254 856
rect 308422 734 309450 856
rect 309618 734 310554 856
rect 310722 734 311750 856
rect 311918 734 312854 856
rect 313022 734 313958 856
rect 314126 734 315154 856
rect 315322 734 316258 856
rect 316426 734 317362 856
rect 317530 734 318558 856
rect 318726 734 319662 856
rect 319830 734 320766 856
rect 320934 734 321962 856
rect 322130 734 323066 856
rect 323234 734 324170 856
rect 324338 734 325366 856
rect 325534 734 326470 856
rect 326638 734 327574 856
rect 327742 734 328770 856
rect 328938 734 329874 856
rect 330042 734 330978 856
rect 331146 734 332174 856
rect 332342 734 333278 856
rect 333446 734 334382 856
rect 334550 734 335578 856
rect 335746 734 336682 856
rect 336850 734 337878 856
rect 338046 734 338982 856
rect 339150 734 340086 856
rect 340254 734 341282 856
rect 341450 734 342386 856
rect 342554 734 343490 856
rect 343658 734 344686 856
rect 344854 734 345790 856
rect 345958 734 346894 856
rect 347062 734 348090 856
rect 348258 734 349194 856
rect 349362 734 350298 856
rect 350466 734 351494 856
rect 351662 734 352598 856
rect 352766 734 353702 856
rect 353870 734 354898 856
rect 355066 734 356002 856
rect 356170 734 357106 856
rect 357274 734 358302 856
rect 358470 734 359406 856
rect 359574 734 360510 856
rect 360678 734 361706 856
rect 361874 734 362810 856
rect 362978 734 363914 856
rect 364082 734 365110 856
rect 365278 734 366214 856
rect 366382 734 367410 856
rect 367578 734 368514 856
rect 368682 734 369618 856
rect 369786 734 370814 856
rect 370982 734 371918 856
rect 372086 734 373022 856
rect 373190 734 374218 856
rect 374386 734 375322 856
rect 375490 734 376426 856
rect 376594 734 377622 856
rect 377790 734 378726 856
rect 378894 734 379830 856
rect 379998 734 381026 856
rect 381194 734 382130 856
rect 382298 734 383234 856
rect 383402 734 384430 856
rect 384598 734 385534 856
rect 385702 734 386638 856
rect 386806 734 387834 856
rect 388002 734 388938 856
rect 389106 734 390042 856
rect 390210 734 391238 856
rect 391406 734 392342 856
rect 392510 734 393538 856
rect 393706 734 394642 856
rect 394810 734 395746 856
rect 395914 734 396942 856
rect 397110 734 398046 856
rect 398214 734 399150 856
rect 399318 734 400346 856
rect 400514 734 401450 856
rect 401618 734 402554 856
rect 402722 734 403750 856
rect 403918 734 404854 856
rect 405022 734 405958 856
rect 406126 734 407154 856
rect 407322 734 408258 856
rect 408426 734 409362 856
rect 409530 734 410558 856
rect 410726 734 411662 856
rect 411830 734 412766 856
rect 412934 734 413962 856
rect 414130 734 415066 856
rect 415234 734 416170 856
rect 416338 734 417366 856
rect 417534 734 418470 856
rect 418638 734 419574 856
rect 419742 734 420770 856
rect 420938 734 421874 856
rect 422042 734 423070 856
rect 423238 734 424174 856
rect 424342 734 425278 856
rect 425446 734 426474 856
rect 426642 734 427578 856
rect 427746 734 428682 856
rect 428850 734 429878 856
rect 430046 734 430982 856
rect 431150 734 432086 856
rect 432254 734 433282 856
rect 433450 734 434386 856
rect 434554 734 435490 856
rect 435658 734 436686 856
rect 436854 734 437790 856
rect 437958 734 438894 856
rect 439062 734 440090 856
rect 440258 734 441194 856
rect 441362 734 442298 856
rect 442466 734 443494 856
rect 443662 734 444598 856
rect 444766 734 445702 856
rect 445870 734 446898 856
rect 447066 734 448002 856
rect 448170 734 449198 856
rect 449366 734 450302 856
rect 450470 734 451406 856
rect 451574 734 452602 856
rect 452770 734 453706 856
rect 453874 734 454810 856
rect 454978 734 456006 856
rect 456174 734 457110 856
rect 457278 734 458214 856
rect 458382 734 459410 856
rect 459578 734 460514 856
rect 460682 734 461618 856
rect 461786 734 462814 856
rect 462982 734 463918 856
rect 464086 734 465022 856
rect 465190 734 466218 856
rect 466386 734 467322 856
rect 467490 734 468426 856
rect 468594 734 469622 856
rect 469790 734 470726 856
rect 470894 734 471830 856
rect 471998 734 473026 856
rect 473194 734 474130 856
rect 474298 734 475234 856
rect 475402 734 476430 856
rect 476598 734 477534 856
rect 477702 734 478730 856
rect 478898 734 479834 856
rect 480002 734 480938 856
rect 481106 734 482134 856
rect 482302 734 483238 856
rect 483406 734 484342 856
rect 484510 734 485538 856
rect 485706 734 486642 856
rect 486810 734 487746 856
rect 487914 734 488942 856
rect 489110 734 490046 856
rect 490214 734 491150 856
rect 491318 734 492346 856
rect 492514 734 493450 856
rect 493618 734 494554 856
rect 494722 734 495750 856
rect 495918 734 496854 856
rect 497022 734 497958 856
rect 498126 734 499154 856
rect 499322 734 500258 856
rect 500426 734 501362 856
rect 501530 734 502558 856
rect 502726 734 503662 856
rect 503830 734 504858 856
rect 505026 734 505962 856
rect 506130 734 507066 856
rect 507234 734 508262 856
rect 508430 734 509366 856
rect 509534 734 510470 856
rect 510638 734 511666 856
rect 511834 734 512770 856
rect 512938 734 513874 856
rect 514042 734 515070 856
rect 515238 734 516174 856
rect 516342 734 517278 856
rect 517446 734 518474 856
rect 518642 734 519578 856
rect 519746 734 520682 856
rect 520850 734 521878 856
rect 522046 734 522982 856
rect 523150 734 524086 856
rect 524254 734 525282 856
rect 525450 734 526386 856
rect 526554 734 527490 856
rect 527658 734 528686 856
rect 528854 734 529790 856
rect 529958 734 530894 856
rect 531062 734 532090 856
rect 532258 734 533194 856
rect 533362 734 534390 856
rect 534558 734 535494 856
rect 535662 734 536598 856
rect 536766 734 537794 856
rect 537962 734 538898 856
rect 539066 734 540002 856
rect 540170 734 541198 856
rect 541366 734 542302 856
rect 542470 734 543406 856
rect 543574 734 544602 856
rect 544770 734 545706 856
rect 545874 734 546810 856
rect 546978 734 548006 856
rect 548174 734 549110 856
rect 549278 734 550214 856
rect 550382 734 551410 856
rect 551578 734 552514 856
rect 552682 734 553618 856
rect 553786 734 554814 856
rect 554982 734 555918 856
rect 556086 734 557022 856
rect 557190 734 558218 856
rect 558386 734 559322 856
<< obsm3 >>
rect 3417 2143 557488 697441
<< metal4 >>
rect 4208 2128 4528 697456
rect 19568 2128 19888 697456
rect 34928 2128 35248 697456
rect 50288 2128 50608 697456
rect 65648 2128 65968 697456
rect 81008 2128 81328 697456
rect 96368 2128 96688 697456
rect 111728 2128 112048 697456
rect 127088 2128 127408 697456
rect 142448 2128 142768 697456
rect 157808 2128 158128 697456
rect 173168 2128 173488 697456
rect 188528 2128 188848 697456
rect 203888 2128 204208 697456
rect 219248 2128 219568 697456
rect 234608 2128 234928 697456
rect 249968 2128 250288 697456
rect 265328 2128 265648 697456
rect 280688 2128 281008 697456
rect 296048 2128 296368 697456
rect 311408 2128 311728 697456
rect 326768 2128 327088 697456
rect 342128 2128 342448 697456
rect 357488 2128 357808 697456
rect 372848 2128 373168 697456
rect 388208 2128 388528 697456
rect 403568 2128 403888 697456
rect 418928 2128 419248 697456
rect 434288 2128 434608 697456
rect 449648 2128 449968 697456
rect 465008 2128 465328 697456
rect 480368 2128 480688 697456
rect 495728 2128 496048 697456
rect 511088 2128 511408 697456
rect 526448 2128 526768 697456
rect 541808 2128 542128 697456
rect 557168 2128 557488 697456
<< obsm4 >>
rect 28395 29275 34848 238781
rect 35328 29275 50208 238781
rect 50688 29275 65568 238781
rect 66048 29275 80928 238781
rect 81408 29275 96288 238781
rect 96768 29275 111648 238781
rect 112128 29275 127008 238781
rect 127488 29275 142368 238781
rect 142848 29275 157728 238781
rect 158208 29275 173088 238781
rect 173568 29275 188448 238781
rect 188928 29275 193141 238781
<< labels >>
rlabel metal2 s 2410 699200 2466 700000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 149702 699200 149758 700000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 164514 699200 164570 700000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 179234 699200 179290 700000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 193954 699200 194010 700000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 208674 699200 208730 700000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 223394 699200 223450 700000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 238114 699200 238170 700000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 252926 699200 252982 700000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 267646 699200 267702 700000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 282366 699200 282422 700000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 17130 699200 17186 700000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 297086 699200 297142 700000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 311806 699200 311862 700000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 326618 699200 326674 700000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 341338 699200 341394 700000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 356058 699200 356114 700000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 370778 699200 370834 700000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 385498 699200 385554 700000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 400218 699200 400274 700000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 415030 699200 415086 700000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 429750 699200 429806 700000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 31850 699200 31906 700000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 444470 699200 444526 700000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 459190 699200 459246 700000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 473910 699200 473966 700000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 488722 699200 488778 700000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 503442 699200 503498 700000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 518162 699200 518218 700000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 532882 699200 532938 700000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 547602 699200 547658 700000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 46570 699200 46626 700000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 61290 699200 61346 700000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 76010 699200 76066 700000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 90822 699200 90878 700000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 105542 699200 105598 700000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 120262 699200 120318 700000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 134982 699200 135038 700000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 7286 699200 7342 700000 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 154670 699200 154726 700000 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 169390 699200 169446 700000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 184110 699200 184166 700000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 198830 699200 198886 700000 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 213550 699200 213606 700000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 228362 699200 228418 700000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 243082 699200 243138 700000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 257802 699200 257858 700000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 272522 699200 272578 700000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 287242 699200 287298 700000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 22006 699200 22062 700000 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 302054 699200 302110 700000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 316774 699200 316830 700000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 331494 699200 331550 700000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 346214 699200 346270 700000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 360934 699200 360990 700000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 375746 699200 375802 700000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 390466 699200 390522 700000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 405186 699200 405242 700000 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 419906 699200 419962 700000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 434626 699200 434682 700000 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 36726 699200 36782 700000 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 449346 699200 449402 700000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 464158 699200 464214 700000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 478878 699200 478934 700000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 493598 699200 493654 700000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 508318 699200 508374 700000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 523038 699200 523094 700000 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 537850 699200 537906 700000 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 552570 699200 552626 700000 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 51446 699200 51502 700000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 66258 699200 66314 700000 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 80978 699200 81034 700000 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 95698 699200 95754 700000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 110418 699200 110474 700000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 125138 699200 125194 700000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 139950 699200 140006 700000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 12162 699200 12218 700000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 159546 699200 159602 700000 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 174266 699200 174322 700000 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 189078 699200 189134 700000 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 203798 699200 203854 700000 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 218518 699200 218574 700000 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 233238 699200 233294 700000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 247958 699200 248014 700000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 262678 699200 262734 700000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 277490 699200 277546 700000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 292210 699200 292266 700000 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 26882 699200 26938 700000 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 306930 699200 306986 700000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 321650 699200 321706 700000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 336370 699200 336426 700000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 351182 699200 351238 700000 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 365902 699200 365958 700000 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 380622 699200 380678 700000 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 395342 699200 395398 700000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 410062 699200 410118 700000 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 424782 699200 424838 700000 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 439594 699200 439650 700000 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 41694 699200 41750 700000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 454314 699200 454370 700000 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 469034 699200 469090 700000 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 483754 699200 483810 700000 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 498474 699200 498530 700000 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 513286 699200 513342 700000 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 528006 699200 528062 700000 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 542726 699200 542782 700000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 557446 699200 557502 700000 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 56414 699200 56470 700000 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 71134 699200 71190 700000 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 85854 699200 85910 700000 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 100574 699200 100630 700000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 115386 699200 115442 700000 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 130106 699200 130162 700000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 144826 699200 144882 700000 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 557078 0 557134 800 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 558274 0 558330 800 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 559378 0 559434 800 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 120906 0 120962 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 461674 0 461730 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 465078 0 465134 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 468482 0 468538 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 471886 0 471942 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 475290 0 475346 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 478786 0 478842 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 482190 0 482246 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 485594 0 485650 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 488998 0 489054 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 492402 0 492458 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 155038 0 155094 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 495806 0 495862 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 499210 0 499266 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 502614 0 502670 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 506018 0 506074 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 509422 0 509478 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 512826 0 512882 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 516230 0 516286 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 519634 0 519690 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 523038 0 523094 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 526442 0 526498 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 158442 0 158498 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 529846 0 529902 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 533250 0 533306 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 536654 0 536710 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 540058 0 540114 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 543462 0 543518 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 546866 0 546922 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 550270 0 550326 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 553674 0 553730 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 161846 0 161902 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 165250 0 165306 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 168654 0 168710 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 172058 0 172114 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 175462 0 175518 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 178866 0 178922 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 182270 0 182326 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 185674 0 185730 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 124310 0 124366 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 189078 0 189134 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 192482 0 192538 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 195886 0 195942 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 199290 0 199346 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 202694 0 202750 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 206098 0 206154 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 209502 0 209558 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 212906 0 212962 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 216310 0 216366 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 219714 0 219770 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 127714 0 127770 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 223118 0 223174 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 226614 0 226670 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 230018 0 230074 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 233422 0 233478 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 236826 0 236882 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 240230 0 240286 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 243634 0 243690 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 247038 0 247094 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 250442 0 250498 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 253846 0 253902 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 131118 0 131174 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 257250 0 257306 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 260654 0 260710 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 264058 0 264114 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 267462 0 267518 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 270866 0 270922 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 274270 0 274326 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 277674 0 277730 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 281078 0 281134 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 284482 0 284538 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 287886 0 287942 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 134522 0 134578 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 291290 0 291346 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 294694 0 294750 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 298098 0 298154 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 301502 0 301558 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 304906 0 304962 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 308310 0 308366 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 311806 0 311862 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 315210 0 315266 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 318614 0 318670 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 322018 0 322074 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 137926 0 137982 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 325422 0 325478 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 328826 0 328882 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 332230 0 332286 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 335634 0 335690 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 339038 0 339094 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 342442 0 342498 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 345846 0 345902 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 349250 0 349306 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 352654 0 352710 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 356058 0 356114 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 141422 0 141478 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 359462 0 359518 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 362866 0 362922 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 366270 0 366326 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 369674 0 369730 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 373078 0 373134 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 376482 0 376538 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 379886 0 379942 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 383290 0 383346 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 386694 0 386750 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 390098 0 390154 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 144826 0 144882 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 393594 0 393650 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 396998 0 397054 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 400402 0 400458 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 403806 0 403862 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 407210 0 407266 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 410614 0 410670 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 414018 0 414074 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 417422 0 417478 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 420826 0 420882 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 424230 0 424286 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 148230 0 148286 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 427634 0 427690 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 431038 0 431094 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 434442 0 434498 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 437846 0 437902 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 441250 0 441306 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 444654 0 444710 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 448058 0 448114 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 451462 0 451518 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 454866 0 454922 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 458270 0 458326 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 151634 0 151690 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 122102 0 122158 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 462870 0 462926 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 466274 0 466330 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 469678 0 469734 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 473082 0 473138 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 476486 0 476542 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 479890 0 479946 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 483294 0 483350 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 486698 0 486754 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 490102 0 490158 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 493506 0 493562 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 156142 0 156198 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 496910 0 496966 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 500314 0 500370 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 503718 0 503774 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 507122 0 507178 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 510526 0 510582 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 513930 0 513986 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 517334 0 517390 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 520738 0 520794 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 524142 0 524198 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 527546 0 527602 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 159546 0 159602 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 530950 0 531006 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 534446 0 534502 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 537850 0 537906 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 541254 0 541310 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 544658 0 544714 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 548062 0 548118 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 551466 0 551522 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 554870 0 554926 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 162950 0 163006 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 166354 0 166410 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 169758 0 169814 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 173162 0 173218 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 176566 0 176622 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 179970 0 180026 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 183374 0 183430 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 186778 0 186834 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 125506 0 125562 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 190182 0 190238 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 193586 0 193642 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 197082 0 197138 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 200486 0 200542 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 203890 0 203946 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 207294 0 207350 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 210698 0 210754 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 214102 0 214158 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 217506 0 217562 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 220910 0 220966 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 128910 0 128966 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 224314 0 224370 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 227718 0 227774 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 231122 0 231178 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 234526 0 234582 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 237930 0 237986 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 241334 0 241390 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 244738 0 244794 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 248142 0 248198 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 251546 0 251602 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 254950 0 255006 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 132314 0 132370 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 258354 0 258410 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 261758 0 261814 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 265162 0 265218 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 268566 0 268622 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 271970 0 272026 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 275374 0 275430 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 278778 0 278834 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 282274 0 282330 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 285678 0 285734 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 289082 0 289138 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 135718 0 135774 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 292486 0 292542 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 295890 0 295946 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 299294 0 299350 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 302698 0 302754 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 306102 0 306158 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 309506 0 309562 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 312910 0 312966 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 316314 0 316370 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 319718 0 319774 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 323122 0 323178 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 139122 0 139178 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 326526 0 326582 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 329930 0 329986 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 333334 0 333390 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 336738 0 336794 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 340142 0 340198 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 343546 0 343602 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 346950 0 347006 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 350354 0 350410 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 353758 0 353814 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 357162 0 357218 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 142526 0 142582 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 360566 0 360622 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 363970 0 364026 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 367466 0 367522 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 370870 0 370926 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 374274 0 374330 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 377678 0 377734 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 381082 0 381138 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 384486 0 384542 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 387890 0 387946 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 391294 0 391350 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 145930 0 145986 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 394698 0 394754 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 398102 0 398158 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 401506 0 401562 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 404910 0 404966 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 408314 0 408370 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 411718 0 411774 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 415122 0 415178 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 418526 0 418582 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 421930 0 421986 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 425334 0 425390 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 149334 0 149390 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 428738 0 428794 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 432142 0 432198 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 435546 0 435602 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 438950 0 439006 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 442354 0 442410 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 445758 0 445814 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 449254 0 449310 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 452658 0 452714 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 456062 0 456118 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 459466 0 459522 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 152738 0 152794 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 123206 0 123262 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 463974 0 464030 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 467378 0 467434 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 470782 0 470838 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 474186 0 474242 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 477590 0 477646 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 480994 0 481050 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 484398 0 484454 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 487802 0 487858 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 491206 0 491262 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 494610 0 494666 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 157246 0 157302 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 498014 0 498070 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 501418 0 501474 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 504914 0 504970 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 508318 0 508374 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 511722 0 511778 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 515126 0 515182 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 518530 0 518586 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 521934 0 521990 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 525338 0 525394 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 528742 0 528798 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 160650 0 160706 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 532146 0 532202 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 535550 0 535606 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 538954 0 539010 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 542358 0 542414 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 545762 0 545818 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 549166 0 549222 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 552570 0 552626 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 555974 0 556030 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 164054 0 164110 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 167458 0 167514 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 170954 0 171010 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 174358 0 174414 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 177762 0 177818 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 181166 0 181222 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 184570 0 184626 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 187974 0 188030 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 126610 0 126666 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 191378 0 191434 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 194782 0 194838 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 198186 0 198242 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 201590 0 201646 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 204994 0 205050 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 208398 0 208454 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 211802 0 211858 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 215206 0 215262 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 218610 0 218666 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 222014 0 222070 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 130014 0 130070 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 225418 0 225474 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 228822 0 228878 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 232226 0 232282 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 235630 0 235686 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 239034 0 239090 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 242438 0 242494 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 245842 0 245898 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 249246 0 249302 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 252742 0 252798 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 256146 0 256202 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 133418 0 133474 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 259550 0 259606 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 262954 0 263010 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 266358 0 266414 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 269762 0 269818 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 273166 0 273222 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 276570 0 276626 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 279974 0 280030 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 283378 0 283434 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 286782 0 286838 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 290186 0 290242 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 136822 0 136878 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 293590 0 293646 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 296994 0 297050 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 300398 0 300454 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 303802 0 303858 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 307206 0 307262 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 310610 0 310666 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 314014 0 314070 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 317418 0 317474 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 320822 0 320878 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 324226 0 324282 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 140226 0 140282 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 327630 0 327686 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 331034 0 331090 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 334438 0 334494 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 337934 0 337990 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 341338 0 341394 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 344742 0 344798 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 348146 0 348202 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 351550 0 351606 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 354954 0 355010 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 358358 0 358414 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 143630 0 143686 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 361762 0 361818 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 365166 0 365222 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 368570 0 368626 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 371974 0 372030 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 375378 0 375434 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 378782 0 378838 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 382186 0 382242 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 385590 0 385646 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 388994 0 389050 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 392398 0 392454 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 147034 0 147090 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 395802 0 395858 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 399206 0 399262 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 402610 0 402666 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 406014 0 406070 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 409418 0 409474 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 412822 0 412878 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 416226 0 416282 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 419630 0 419686 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 423126 0 423182 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 426530 0 426586 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 150438 0 150494 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 429934 0 429990 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 433338 0 433394 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 436742 0 436798 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 440146 0 440202 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 443550 0 443606 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 446954 0 447010 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 450358 0 450414 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 453762 0 453818 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 457166 0 457222 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 460570 0 460626 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 153842 0 153898 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal4 s 4208 2128 4528 697456 6 vccd1
port 502 nsew power input
rlabel metal4 s 34928 2128 35248 697456 6 vccd1
port 502 nsew power input
rlabel metal4 s 65648 2128 65968 697456 6 vccd1
port 502 nsew power input
rlabel metal4 s 96368 2128 96688 697456 6 vccd1
port 502 nsew power input
rlabel metal4 s 127088 2128 127408 697456 6 vccd1
port 502 nsew power input
rlabel metal4 s 157808 2128 158128 697456 6 vccd1
port 502 nsew power input
rlabel metal4 s 188528 2128 188848 697456 6 vccd1
port 502 nsew power input
rlabel metal4 s 219248 2128 219568 697456 6 vccd1
port 502 nsew power input
rlabel metal4 s 249968 2128 250288 697456 6 vccd1
port 502 nsew power input
rlabel metal4 s 280688 2128 281008 697456 6 vccd1
port 502 nsew power input
rlabel metal4 s 311408 2128 311728 697456 6 vccd1
port 502 nsew power input
rlabel metal4 s 342128 2128 342448 697456 6 vccd1
port 502 nsew power input
rlabel metal4 s 372848 2128 373168 697456 6 vccd1
port 502 nsew power input
rlabel metal4 s 403568 2128 403888 697456 6 vccd1
port 502 nsew power input
rlabel metal4 s 434288 2128 434608 697456 6 vccd1
port 502 nsew power input
rlabel metal4 s 465008 2128 465328 697456 6 vccd1
port 502 nsew power input
rlabel metal4 s 495728 2128 496048 697456 6 vccd1
port 502 nsew power input
rlabel metal4 s 526448 2128 526768 697456 6 vccd1
port 502 nsew power input
rlabel metal4 s 557168 2128 557488 697456 6 vccd1
port 502 nsew power input
rlabel metal4 s 19568 2128 19888 697456 6 vssd1
port 503 nsew ground input
rlabel metal4 s 50288 2128 50608 697456 6 vssd1
port 503 nsew ground input
rlabel metal4 s 81008 2128 81328 697456 6 vssd1
port 503 nsew ground input
rlabel metal4 s 111728 2128 112048 697456 6 vssd1
port 503 nsew ground input
rlabel metal4 s 142448 2128 142768 697456 6 vssd1
port 503 nsew ground input
rlabel metal4 s 173168 2128 173488 697456 6 vssd1
port 503 nsew ground input
rlabel metal4 s 203888 2128 204208 697456 6 vssd1
port 503 nsew ground input
rlabel metal4 s 234608 2128 234928 697456 6 vssd1
port 503 nsew ground input
rlabel metal4 s 265328 2128 265648 697456 6 vssd1
port 503 nsew ground input
rlabel metal4 s 296048 2128 296368 697456 6 vssd1
port 503 nsew ground input
rlabel metal4 s 326768 2128 327088 697456 6 vssd1
port 503 nsew ground input
rlabel metal4 s 357488 2128 357808 697456 6 vssd1
port 503 nsew ground input
rlabel metal4 s 388208 2128 388528 697456 6 vssd1
port 503 nsew ground input
rlabel metal4 s 418928 2128 419248 697456 6 vssd1
port 503 nsew ground input
rlabel metal4 s 449648 2128 449968 697456 6 vssd1
port 503 nsew ground input
rlabel metal4 s 480368 2128 480688 697456 6 vssd1
port 503 nsew ground input
rlabel metal4 s 511088 2128 511408 697456 6 vssd1
port 503 nsew ground input
rlabel metal4 s 541808 2128 542128 697456 6 vssd1
port 503 nsew ground input
rlabel metal2 s 570 0 626 800 6 wb_clk_i
port 504 nsew signal input
rlabel metal2 s 1674 0 1730 800 6 wb_rst_i
port 505 nsew signal input
rlabel metal2 s 2778 0 2834 800 6 wbs_ack_o
port 506 nsew signal output
rlabel metal2 s 7378 0 7434 800 6 wbs_adr_i[0]
port 507 nsew signal input
rlabel metal2 s 45926 0 45982 800 6 wbs_adr_i[10]
port 508 nsew signal input
rlabel metal2 s 49330 0 49386 800 6 wbs_adr_i[11]
port 509 nsew signal input
rlabel metal2 s 52734 0 52790 800 6 wbs_adr_i[12]
port 510 nsew signal input
rlabel metal2 s 56138 0 56194 800 6 wbs_adr_i[13]
port 511 nsew signal input
rlabel metal2 s 59634 0 59690 800 6 wbs_adr_i[14]
port 512 nsew signal input
rlabel metal2 s 63038 0 63094 800 6 wbs_adr_i[15]
port 513 nsew signal input
rlabel metal2 s 66442 0 66498 800 6 wbs_adr_i[16]
port 514 nsew signal input
rlabel metal2 s 69846 0 69902 800 6 wbs_adr_i[17]
port 515 nsew signal input
rlabel metal2 s 73250 0 73306 800 6 wbs_adr_i[18]
port 516 nsew signal input
rlabel metal2 s 76654 0 76710 800 6 wbs_adr_i[19]
port 517 nsew signal input
rlabel metal2 s 11886 0 11942 800 6 wbs_adr_i[1]
port 518 nsew signal input
rlabel metal2 s 80058 0 80114 800 6 wbs_adr_i[20]
port 519 nsew signal input
rlabel metal2 s 83462 0 83518 800 6 wbs_adr_i[21]
port 520 nsew signal input
rlabel metal2 s 86866 0 86922 800 6 wbs_adr_i[22]
port 521 nsew signal input
rlabel metal2 s 90270 0 90326 800 6 wbs_adr_i[23]
port 522 nsew signal input
rlabel metal2 s 93674 0 93730 800 6 wbs_adr_i[24]
port 523 nsew signal input
rlabel metal2 s 97078 0 97134 800 6 wbs_adr_i[25]
port 524 nsew signal input
rlabel metal2 s 100482 0 100538 800 6 wbs_adr_i[26]
port 525 nsew signal input
rlabel metal2 s 103886 0 103942 800 6 wbs_adr_i[27]
port 526 nsew signal input
rlabel metal2 s 107290 0 107346 800 6 wbs_adr_i[28]
port 527 nsew signal input
rlabel metal2 s 110694 0 110750 800 6 wbs_adr_i[29]
port 528 nsew signal input
rlabel metal2 s 16394 0 16450 800 6 wbs_adr_i[2]
port 529 nsew signal input
rlabel metal2 s 114098 0 114154 800 6 wbs_adr_i[30]
port 530 nsew signal input
rlabel metal2 s 117502 0 117558 800 6 wbs_adr_i[31]
port 531 nsew signal input
rlabel metal2 s 20994 0 21050 800 6 wbs_adr_i[3]
port 532 nsew signal input
rlabel metal2 s 25502 0 25558 800 6 wbs_adr_i[4]
port 533 nsew signal input
rlabel metal2 s 28906 0 28962 800 6 wbs_adr_i[5]
port 534 nsew signal input
rlabel metal2 s 32310 0 32366 800 6 wbs_adr_i[6]
port 535 nsew signal input
rlabel metal2 s 35714 0 35770 800 6 wbs_adr_i[7]
port 536 nsew signal input
rlabel metal2 s 39118 0 39174 800 6 wbs_adr_i[8]
port 537 nsew signal input
rlabel metal2 s 42522 0 42578 800 6 wbs_adr_i[9]
port 538 nsew signal input
rlabel metal2 s 3974 0 4030 800 6 wbs_cyc_i
port 539 nsew signal input
rlabel metal2 s 8482 0 8538 800 6 wbs_dat_i[0]
port 540 nsew signal input
rlabel metal2 s 47122 0 47178 800 6 wbs_dat_i[10]
port 541 nsew signal input
rlabel metal2 s 50526 0 50582 800 6 wbs_dat_i[11]
port 542 nsew signal input
rlabel metal2 s 53930 0 53986 800 6 wbs_dat_i[12]
port 543 nsew signal input
rlabel metal2 s 57334 0 57390 800 6 wbs_dat_i[13]
port 544 nsew signal input
rlabel metal2 s 60738 0 60794 800 6 wbs_dat_i[14]
port 545 nsew signal input
rlabel metal2 s 64142 0 64198 800 6 wbs_dat_i[15]
port 546 nsew signal input
rlabel metal2 s 67546 0 67602 800 6 wbs_dat_i[16]
port 547 nsew signal input
rlabel metal2 s 70950 0 71006 800 6 wbs_dat_i[17]
port 548 nsew signal input
rlabel metal2 s 74354 0 74410 800 6 wbs_dat_i[18]
port 549 nsew signal input
rlabel metal2 s 77758 0 77814 800 6 wbs_dat_i[19]
port 550 nsew signal input
rlabel metal2 s 12990 0 13046 800 6 wbs_dat_i[1]
port 551 nsew signal input
rlabel metal2 s 81162 0 81218 800 6 wbs_dat_i[20]
port 552 nsew signal input
rlabel metal2 s 84566 0 84622 800 6 wbs_dat_i[21]
port 553 nsew signal input
rlabel metal2 s 87970 0 88026 800 6 wbs_dat_i[22]
port 554 nsew signal input
rlabel metal2 s 91374 0 91430 800 6 wbs_dat_i[23]
port 555 nsew signal input
rlabel metal2 s 94778 0 94834 800 6 wbs_dat_i[24]
port 556 nsew signal input
rlabel metal2 s 98182 0 98238 800 6 wbs_dat_i[25]
port 557 nsew signal input
rlabel metal2 s 101586 0 101642 800 6 wbs_dat_i[26]
port 558 nsew signal input
rlabel metal2 s 104990 0 105046 800 6 wbs_dat_i[27]
port 559 nsew signal input
rlabel metal2 s 108394 0 108450 800 6 wbs_dat_i[28]
port 560 nsew signal input
rlabel metal2 s 111798 0 111854 800 6 wbs_dat_i[29]
port 561 nsew signal input
rlabel metal2 s 17590 0 17646 800 6 wbs_dat_i[2]
port 562 nsew signal input
rlabel metal2 s 115294 0 115350 800 6 wbs_dat_i[30]
port 563 nsew signal input
rlabel metal2 s 118698 0 118754 800 6 wbs_dat_i[31]
port 564 nsew signal input
rlabel metal2 s 22098 0 22154 800 6 wbs_dat_i[3]
port 565 nsew signal input
rlabel metal2 s 26606 0 26662 800 6 wbs_dat_i[4]
port 566 nsew signal input
rlabel metal2 s 30102 0 30158 800 6 wbs_dat_i[5]
port 567 nsew signal input
rlabel metal2 s 33506 0 33562 800 6 wbs_dat_i[6]
port 568 nsew signal input
rlabel metal2 s 36910 0 36966 800 6 wbs_dat_i[7]
port 569 nsew signal input
rlabel metal2 s 40314 0 40370 800 6 wbs_dat_i[8]
port 570 nsew signal input
rlabel metal2 s 43718 0 43774 800 6 wbs_dat_i[9]
port 571 nsew signal input
rlabel metal2 s 9586 0 9642 800 6 wbs_dat_o[0]
port 572 nsew signal output
rlabel metal2 s 48226 0 48282 800 6 wbs_dat_o[10]
port 573 nsew signal output
rlabel metal2 s 51630 0 51686 800 6 wbs_dat_o[11]
port 574 nsew signal output
rlabel metal2 s 55034 0 55090 800 6 wbs_dat_o[12]
port 575 nsew signal output
rlabel metal2 s 58438 0 58494 800 6 wbs_dat_o[13]
port 576 nsew signal output
rlabel metal2 s 61842 0 61898 800 6 wbs_dat_o[14]
port 577 nsew signal output
rlabel metal2 s 65246 0 65302 800 6 wbs_dat_o[15]
port 578 nsew signal output
rlabel metal2 s 68650 0 68706 800 6 wbs_dat_o[16]
port 579 nsew signal output
rlabel metal2 s 72054 0 72110 800 6 wbs_dat_o[17]
port 580 nsew signal output
rlabel metal2 s 75458 0 75514 800 6 wbs_dat_o[18]
port 581 nsew signal output
rlabel metal2 s 78862 0 78918 800 6 wbs_dat_o[19]
port 582 nsew signal output
rlabel metal2 s 14186 0 14242 800 6 wbs_dat_o[1]
port 583 nsew signal output
rlabel metal2 s 82266 0 82322 800 6 wbs_dat_o[20]
port 584 nsew signal output
rlabel metal2 s 85762 0 85818 800 6 wbs_dat_o[21]
port 585 nsew signal output
rlabel metal2 s 89166 0 89222 800 6 wbs_dat_o[22]
port 586 nsew signal output
rlabel metal2 s 92570 0 92626 800 6 wbs_dat_o[23]
port 587 nsew signal output
rlabel metal2 s 95974 0 96030 800 6 wbs_dat_o[24]
port 588 nsew signal output
rlabel metal2 s 99378 0 99434 800 6 wbs_dat_o[25]
port 589 nsew signal output
rlabel metal2 s 102782 0 102838 800 6 wbs_dat_o[26]
port 590 nsew signal output
rlabel metal2 s 106186 0 106242 800 6 wbs_dat_o[27]
port 591 nsew signal output
rlabel metal2 s 109590 0 109646 800 6 wbs_dat_o[28]
port 592 nsew signal output
rlabel metal2 s 112994 0 113050 800 6 wbs_dat_o[29]
port 593 nsew signal output
rlabel metal2 s 18694 0 18750 800 6 wbs_dat_o[2]
port 594 nsew signal output
rlabel metal2 s 116398 0 116454 800 6 wbs_dat_o[30]
port 595 nsew signal output
rlabel metal2 s 119802 0 119858 800 6 wbs_dat_o[31]
port 596 nsew signal output
rlabel metal2 s 23202 0 23258 800 6 wbs_dat_o[3]
port 597 nsew signal output
rlabel metal2 s 27802 0 27858 800 6 wbs_dat_o[4]
port 598 nsew signal output
rlabel metal2 s 31206 0 31262 800 6 wbs_dat_o[5]
port 599 nsew signal output
rlabel metal2 s 34610 0 34666 800 6 wbs_dat_o[6]
port 600 nsew signal output
rlabel metal2 s 38014 0 38070 800 6 wbs_dat_o[7]
port 601 nsew signal output
rlabel metal2 s 41418 0 41474 800 6 wbs_dat_o[8]
port 602 nsew signal output
rlabel metal2 s 44822 0 44878 800 6 wbs_dat_o[9]
port 603 nsew signal output
rlabel metal2 s 10782 0 10838 800 6 wbs_sel_i[0]
port 604 nsew signal input
rlabel metal2 s 15290 0 15346 800 6 wbs_sel_i[1]
port 605 nsew signal input
rlabel metal2 s 19798 0 19854 800 6 wbs_sel_i[2]
port 606 nsew signal input
rlabel metal2 s 24398 0 24454 800 6 wbs_sel_i[3]
port 607 nsew signal input
rlabel metal2 s 5078 0 5134 800 6 wbs_stb_i
port 608 nsew signal input
rlabel metal2 s 6182 0 6238 800 6 wbs_we_i
port 609 nsew signal input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 560000 700000
string LEFview TRUE
string GDS_FILE /project/openlane/user_proj/runs/user_proj/results/magic/user_proj.gds
string GDS_END 170973788
string GDS_START 1441646
<< end >>

