magic
tech sky130A
magscale 1 2
timestamp 1640797500
<< obsli1 >>
rect 1409 1921 165387 165291
<< obsm1 >>
rect 658 756 165494 167408
<< metal2 >>
rect 478 166914 534 167714
rect 1490 166914 1546 167714
rect 2594 166914 2650 167714
rect 3606 166914 3662 167714
rect 4710 166914 4766 167714
rect 5814 166914 5870 167714
rect 6826 166914 6882 167714
rect 7930 166914 7986 167714
rect 8942 166914 8998 167714
rect 10046 166914 10102 167714
rect 11150 166914 11206 167714
rect 12162 166914 12218 167714
rect 13266 166914 13322 167714
rect 14278 166914 14334 167714
rect 15382 166914 15438 167714
rect 16486 166914 16542 167714
rect 17498 166914 17554 167714
rect 18602 166914 18658 167714
rect 19706 166914 19762 167714
rect 20718 166914 20774 167714
rect 21822 166914 21878 167714
rect 22834 166914 22890 167714
rect 23938 166914 23994 167714
rect 25042 166914 25098 167714
rect 26054 166914 26110 167714
rect 27158 166914 27214 167714
rect 28170 166914 28226 167714
rect 29274 166914 29330 167714
rect 30378 166914 30434 167714
rect 31390 166914 31446 167714
rect 32494 166914 32550 167714
rect 33598 166914 33654 167714
rect 34610 166914 34666 167714
rect 35714 166914 35770 167714
rect 36726 166914 36782 167714
rect 37830 166914 37886 167714
rect 38934 166914 38990 167714
rect 39946 166914 40002 167714
rect 41050 166914 41106 167714
rect 42062 166914 42118 167714
rect 43166 166914 43222 167714
rect 44270 166914 44326 167714
rect 45282 166914 45338 167714
rect 46386 166914 46442 167714
rect 47398 166914 47454 167714
rect 48502 166914 48558 167714
rect 49606 166914 49662 167714
rect 50618 166914 50674 167714
rect 51722 166914 51778 167714
rect 52826 166914 52882 167714
rect 53838 166914 53894 167714
rect 54942 166914 54998 167714
rect 55954 166914 56010 167714
rect 57058 166914 57114 167714
rect 58162 166914 58218 167714
rect 59174 166914 59230 167714
rect 60278 166914 60334 167714
rect 61290 166914 61346 167714
rect 62394 166914 62450 167714
rect 63498 166914 63554 167714
rect 64510 166914 64566 167714
rect 65614 166914 65670 167714
rect 66718 166914 66774 167714
rect 67730 166914 67786 167714
rect 68834 166914 68890 167714
rect 69846 166914 69902 167714
rect 70950 166914 71006 167714
rect 72054 166914 72110 167714
rect 73066 166914 73122 167714
rect 74170 166914 74226 167714
rect 75182 166914 75238 167714
rect 76286 166914 76342 167714
rect 77390 166914 77446 167714
rect 78402 166914 78458 167714
rect 79506 166914 79562 167714
rect 80518 166914 80574 167714
rect 81622 166914 81678 167714
rect 82726 166914 82782 167714
rect 83738 166914 83794 167714
rect 84842 166914 84898 167714
rect 85946 166914 86002 167714
rect 86958 166914 87014 167714
rect 88062 166914 88118 167714
rect 89074 166914 89130 167714
rect 90178 166914 90234 167714
rect 91282 166914 91338 167714
rect 92294 166914 92350 167714
rect 93398 166914 93454 167714
rect 94410 166914 94466 167714
rect 95514 166914 95570 167714
rect 96618 166914 96674 167714
rect 97630 166914 97686 167714
rect 98734 166914 98790 167714
rect 99838 166914 99894 167714
rect 100850 166914 100906 167714
rect 101954 166914 102010 167714
rect 102966 166914 103022 167714
rect 104070 166914 104126 167714
rect 105174 166914 105230 167714
rect 106186 166914 106242 167714
rect 107290 166914 107346 167714
rect 108302 166914 108358 167714
rect 109406 166914 109462 167714
rect 110510 166914 110566 167714
rect 111522 166914 111578 167714
rect 112626 166914 112682 167714
rect 113638 166914 113694 167714
rect 114742 166914 114798 167714
rect 115846 166914 115902 167714
rect 116858 166914 116914 167714
rect 117962 166914 118018 167714
rect 119066 166914 119122 167714
rect 120078 166914 120134 167714
rect 121182 166914 121238 167714
rect 122194 166914 122250 167714
rect 123298 166914 123354 167714
rect 124402 166914 124458 167714
rect 125414 166914 125470 167714
rect 126518 166914 126574 167714
rect 127530 166914 127586 167714
rect 128634 166914 128690 167714
rect 129738 166914 129794 167714
rect 130750 166914 130806 167714
rect 131854 166914 131910 167714
rect 132958 166914 133014 167714
rect 133970 166914 134026 167714
rect 135074 166914 135130 167714
rect 136086 166914 136142 167714
rect 137190 166914 137246 167714
rect 138294 166914 138350 167714
rect 139306 166914 139362 167714
rect 140410 166914 140466 167714
rect 141422 166914 141478 167714
rect 142526 166914 142582 167714
rect 143630 166914 143686 167714
rect 144642 166914 144698 167714
rect 145746 166914 145802 167714
rect 146758 166914 146814 167714
rect 147862 166914 147918 167714
rect 148966 166914 149022 167714
rect 149978 166914 150034 167714
rect 151082 166914 151138 167714
rect 152186 166914 152242 167714
rect 153198 166914 153254 167714
rect 154302 166914 154358 167714
rect 155314 166914 155370 167714
rect 156418 166914 156474 167714
rect 157522 166914 157578 167714
rect 158534 166914 158590 167714
rect 159638 166914 159694 167714
rect 160650 166914 160706 167714
rect 161754 166914 161810 167714
rect 162858 166914 162914 167714
rect 163870 166914 163926 167714
rect 164974 166914 165030 167714
rect 570 0 626 800
rect 1674 0 1730 800
rect 2870 0 2926 800
rect 4066 0 4122 800
rect 5262 0 5318 800
rect 6366 0 6422 800
rect 7562 0 7618 800
rect 8758 0 8814 800
rect 9954 0 10010 800
rect 11058 0 11114 800
rect 12254 0 12310 800
rect 13450 0 13506 800
rect 14646 0 14702 800
rect 15750 0 15806 800
rect 16946 0 17002 800
rect 18142 0 18198 800
rect 19338 0 19394 800
rect 20534 0 20590 800
rect 21638 0 21694 800
rect 22834 0 22890 800
rect 24030 0 24086 800
rect 25226 0 25282 800
rect 26330 0 26386 800
rect 27526 0 27582 800
rect 28722 0 28778 800
rect 29918 0 29974 800
rect 31022 0 31078 800
rect 32218 0 32274 800
rect 33414 0 33470 800
rect 34610 0 34666 800
rect 35714 0 35770 800
rect 36910 0 36966 800
rect 38106 0 38162 800
rect 39302 0 39358 800
rect 40498 0 40554 800
rect 41602 0 41658 800
rect 42798 0 42854 800
rect 43994 0 44050 800
rect 45190 0 45246 800
rect 46294 0 46350 800
rect 47490 0 47546 800
rect 48686 0 48742 800
rect 49882 0 49938 800
rect 50986 0 51042 800
rect 52182 0 52238 800
rect 53378 0 53434 800
rect 54574 0 54630 800
rect 55770 0 55826 800
rect 56874 0 56930 800
rect 58070 0 58126 800
rect 59266 0 59322 800
rect 60462 0 60518 800
rect 61566 0 61622 800
rect 62762 0 62818 800
rect 63958 0 64014 800
rect 65154 0 65210 800
rect 66258 0 66314 800
rect 67454 0 67510 800
rect 68650 0 68706 800
rect 69846 0 69902 800
rect 70950 0 71006 800
rect 72146 0 72202 800
rect 73342 0 73398 800
rect 74538 0 74594 800
rect 75734 0 75790 800
rect 76838 0 76894 800
rect 78034 0 78090 800
rect 79230 0 79286 800
rect 80426 0 80482 800
rect 81530 0 81586 800
rect 82726 0 82782 800
rect 83922 0 83978 800
rect 85118 0 85174 800
rect 86222 0 86278 800
rect 87418 0 87474 800
rect 88614 0 88670 800
rect 89810 0 89866 800
rect 90914 0 90970 800
rect 92110 0 92166 800
rect 93306 0 93362 800
rect 94502 0 94558 800
rect 95698 0 95754 800
rect 96802 0 96858 800
rect 97998 0 98054 800
rect 99194 0 99250 800
rect 100390 0 100446 800
rect 101494 0 101550 800
rect 102690 0 102746 800
rect 103886 0 103942 800
rect 105082 0 105138 800
rect 106186 0 106242 800
rect 107382 0 107438 800
rect 108578 0 108634 800
rect 109774 0 109830 800
rect 110970 0 111026 800
rect 112074 0 112130 800
rect 113270 0 113326 800
rect 114466 0 114522 800
rect 115662 0 115718 800
rect 116766 0 116822 800
rect 117962 0 118018 800
rect 119158 0 119214 800
rect 120354 0 120410 800
rect 121458 0 121514 800
rect 122654 0 122710 800
rect 123850 0 123906 800
rect 125046 0 125102 800
rect 126150 0 126206 800
rect 127346 0 127402 800
rect 128542 0 128598 800
rect 129738 0 129794 800
rect 130934 0 130990 800
rect 132038 0 132094 800
rect 133234 0 133290 800
rect 134430 0 134486 800
rect 135626 0 135682 800
rect 136730 0 136786 800
rect 137926 0 137982 800
rect 139122 0 139178 800
rect 140318 0 140374 800
rect 141422 0 141478 800
rect 142618 0 142674 800
rect 143814 0 143870 800
rect 145010 0 145066 800
rect 146114 0 146170 800
rect 147310 0 147366 800
rect 148506 0 148562 800
rect 149702 0 149758 800
rect 150898 0 150954 800
rect 152002 0 152058 800
rect 153198 0 153254 800
rect 154394 0 154450 800
rect 155590 0 155646 800
rect 156694 0 156750 800
rect 157890 0 157946 800
rect 159086 0 159142 800
rect 160282 0 160338 800
rect 161386 0 161442 800
rect 162582 0 162638 800
rect 163778 0 163834 800
rect 164974 0 165030 800
<< obsm2 >>
rect 18 166858 422 167657
rect 590 166858 1434 167657
rect 1602 166858 2538 167657
rect 2706 166858 3550 167657
rect 3718 166858 4654 167657
rect 4822 166858 5758 167657
rect 5926 166858 6770 167657
rect 6938 166858 7874 167657
rect 8042 166858 8886 167657
rect 9054 166858 9990 167657
rect 10158 166858 11094 167657
rect 11262 166858 12106 167657
rect 12274 166858 13210 167657
rect 13378 166858 14222 167657
rect 14390 166858 15326 167657
rect 15494 166858 16430 167657
rect 16598 166858 17442 167657
rect 17610 166858 18546 167657
rect 18714 166858 19650 167657
rect 19818 166858 20662 167657
rect 20830 166858 21766 167657
rect 21934 166858 22778 167657
rect 22946 166858 23882 167657
rect 24050 166858 24986 167657
rect 25154 166858 25998 167657
rect 26166 166858 27102 167657
rect 27270 166858 28114 167657
rect 28282 166858 29218 167657
rect 29386 166858 30322 167657
rect 30490 166858 31334 167657
rect 31502 166858 32438 167657
rect 32606 166858 33542 167657
rect 33710 166858 34554 167657
rect 34722 166858 35658 167657
rect 35826 166858 36670 167657
rect 36838 166858 37774 167657
rect 37942 166858 38878 167657
rect 39046 166858 39890 167657
rect 40058 166858 40994 167657
rect 41162 166858 42006 167657
rect 42174 166858 43110 167657
rect 43278 166858 44214 167657
rect 44382 166858 45226 167657
rect 45394 166858 46330 167657
rect 46498 166858 47342 167657
rect 47510 166858 48446 167657
rect 48614 166858 49550 167657
rect 49718 166858 50562 167657
rect 50730 166858 51666 167657
rect 51834 166858 52770 167657
rect 52938 166858 53782 167657
rect 53950 166858 54886 167657
rect 55054 166858 55898 167657
rect 56066 166858 57002 167657
rect 57170 166858 58106 167657
rect 58274 166858 59118 167657
rect 59286 166858 60222 167657
rect 60390 166858 61234 167657
rect 61402 166858 62338 167657
rect 62506 166858 63442 167657
rect 63610 166858 64454 167657
rect 64622 166858 65558 167657
rect 65726 166858 66662 167657
rect 66830 166858 67674 167657
rect 67842 166858 68778 167657
rect 68946 166858 69790 167657
rect 69958 166858 70894 167657
rect 71062 166858 71998 167657
rect 72166 166858 73010 167657
rect 73178 166858 74114 167657
rect 74282 166858 75126 167657
rect 75294 166858 76230 167657
rect 76398 166858 77334 167657
rect 77502 166858 78346 167657
rect 78514 166858 79450 167657
rect 79618 166858 80462 167657
rect 80630 166858 81566 167657
rect 81734 166858 82670 167657
rect 82838 166858 83682 167657
rect 83850 166858 84786 167657
rect 84954 166858 85890 167657
rect 86058 166858 86902 167657
rect 87070 166858 88006 167657
rect 88174 166858 89018 167657
rect 89186 166858 90122 167657
rect 90290 166858 91226 167657
rect 91394 166858 92238 167657
rect 92406 166858 93342 167657
rect 93510 166858 94354 167657
rect 94522 166858 95458 167657
rect 95626 166858 96562 167657
rect 96730 166858 97574 167657
rect 97742 166858 98678 167657
rect 98846 166858 99782 167657
rect 99950 166858 100794 167657
rect 100962 166858 101898 167657
rect 102066 166858 102910 167657
rect 103078 166858 104014 167657
rect 104182 166858 105118 167657
rect 105286 166858 106130 167657
rect 106298 166858 107234 167657
rect 107402 166858 108246 167657
rect 108414 166858 109350 167657
rect 109518 166858 110454 167657
rect 110622 166858 111466 167657
rect 111634 166858 112570 167657
rect 112738 166858 113582 167657
rect 113750 166858 114686 167657
rect 114854 166858 115790 167657
rect 115958 166858 116802 167657
rect 116970 166858 117906 167657
rect 118074 166858 119010 167657
rect 119178 166858 120022 167657
rect 120190 166858 121126 167657
rect 121294 166858 122138 167657
rect 122306 166858 123242 167657
rect 123410 166858 124346 167657
rect 124514 166858 125358 167657
rect 125526 166858 126462 167657
rect 126630 166858 127474 167657
rect 127642 166858 128578 167657
rect 128746 166858 129682 167657
rect 129850 166858 130694 167657
rect 130862 166858 131798 167657
rect 131966 166858 132902 167657
rect 133070 166858 133914 167657
rect 134082 166858 135018 167657
rect 135186 166858 136030 167657
rect 136198 166858 137134 167657
rect 137302 166858 138238 167657
rect 138406 166858 139250 167657
rect 139418 166858 140354 167657
rect 140522 166858 141366 167657
rect 141534 166858 142470 167657
rect 142638 166858 143574 167657
rect 143742 166858 144586 167657
rect 144754 166858 145690 167657
rect 145858 166858 146702 167657
rect 146870 166858 147806 167657
rect 147974 166858 148910 167657
rect 149078 166858 149922 167657
rect 150090 166858 151026 167657
rect 151194 166858 152130 167657
rect 152298 166858 153142 167657
rect 153310 166858 154246 167657
rect 154414 166858 155258 167657
rect 155426 166858 156362 167657
rect 156530 166858 157466 167657
rect 157634 166858 158478 167657
rect 158646 166858 159582 167657
rect 159750 166858 160594 167657
rect 160762 166858 161698 167657
rect 161866 166858 162802 167657
rect 162970 166858 163814 167657
rect 163982 166858 164918 167657
rect 165086 166858 165568 167657
rect 18 856 165568 166858
rect 18 734 514 856
rect 682 734 1618 856
rect 1786 734 2814 856
rect 2982 734 4010 856
rect 4178 734 5206 856
rect 5374 734 6310 856
rect 6478 734 7506 856
rect 7674 734 8702 856
rect 8870 734 9898 856
rect 10066 734 11002 856
rect 11170 734 12198 856
rect 12366 734 13394 856
rect 13562 734 14590 856
rect 14758 734 15694 856
rect 15862 734 16890 856
rect 17058 734 18086 856
rect 18254 734 19282 856
rect 19450 734 20478 856
rect 20646 734 21582 856
rect 21750 734 22778 856
rect 22946 734 23974 856
rect 24142 734 25170 856
rect 25338 734 26274 856
rect 26442 734 27470 856
rect 27638 734 28666 856
rect 28834 734 29862 856
rect 30030 734 30966 856
rect 31134 734 32162 856
rect 32330 734 33358 856
rect 33526 734 34554 856
rect 34722 734 35658 856
rect 35826 734 36854 856
rect 37022 734 38050 856
rect 38218 734 39246 856
rect 39414 734 40442 856
rect 40610 734 41546 856
rect 41714 734 42742 856
rect 42910 734 43938 856
rect 44106 734 45134 856
rect 45302 734 46238 856
rect 46406 734 47434 856
rect 47602 734 48630 856
rect 48798 734 49826 856
rect 49994 734 50930 856
rect 51098 734 52126 856
rect 52294 734 53322 856
rect 53490 734 54518 856
rect 54686 734 55714 856
rect 55882 734 56818 856
rect 56986 734 58014 856
rect 58182 734 59210 856
rect 59378 734 60406 856
rect 60574 734 61510 856
rect 61678 734 62706 856
rect 62874 734 63902 856
rect 64070 734 65098 856
rect 65266 734 66202 856
rect 66370 734 67398 856
rect 67566 734 68594 856
rect 68762 734 69790 856
rect 69958 734 70894 856
rect 71062 734 72090 856
rect 72258 734 73286 856
rect 73454 734 74482 856
rect 74650 734 75678 856
rect 75846 734 76782 856
rect 76950 734 77978 856
rect 78146 734 79174 856
rect 79342 734 80370 856
rect 80538 734 81474 856
rect 81642 734 82670 856
rect 82838 734 83866 856
rect 84034 734 85062 856
rect 85230 734 86166 856
rect 86334 734 87362 856
rect 87530 734 88558 856
rect 88726 734 89754 856
rect 89922 734 90858 856
rect 91026 734 92054 856
rect 92222 734 93250 856
rect 93418 734 94446 856
rect 94614 734 95642 856
rect 95810 734 96746 856
rect 96914 734 97942 856
rect 98110 734 99138 856
rect 99306 734 100334 856
rect 100502 734 101438 856
rect 101606 734 102634 856
rect 102802 734 103830 856
rect 103998 734 105026 856
rect 105194 734 106130 856
rect 106298 734 107326 856
rect 107494 734 108522 856
rect 108690 734 109718 856
rect 109886 734 110914 856
rect 111082 734 112018 856
rect 112186 734 113214 856
rect 113382 734 114410 856
rect 114578 734 115606 856
rect 115774 734 116710 856
rect 116878 734 117906 856
rect 118074 734 119102 856
rect 119270 734 120298 856
rect 120466 734 121402 856
rect 121570 734 122598 856
rect 122766 734 123794 856
rect 123962 734 124990 856
rect 125158 734 126094 856
rect 126262 734 127290 856
rect 127458 734 128486 856
rect 128654 734 129682 856
rect 129850 734 130878 856
rect 131046 734 131982 856
rect 132150 734 133178 856
rect 133346 734 134374 856
rect 134542 734 135570 856
rect 135738 734 136674 856
rect 136842 734 137870 856
rect 138038 734 139066 856
rect 139234 734 140262 856
rect 140430 734 141366 856
rect 141534 734 142562 856
rect 142730 734 143758 856
rect 143926 734 144954 856
rect 145122 734 146058 856
rect 146226 734 147254 856
rect 147422 734 148450 856
rect 148618 734 149646 856
rect 149814 734 150842 856
rect 151010 734 151946 856
rect 152114 734 153142 856
rect 153310 734 154338 856
rect 154506 734 155534 856
rect 155702 734 156638 856
rect 156806 734 157834 856
rect 158002 734 159030 856
rect 159198 734 160226 856
rect 160394 734 161330 856
rect 161498 734 162526 856
rect 162694 734 163722 856
rect 163890 734 164918 856
rect 165086 734 165568 856
<< metal3 >>
rect 0 165792 800 165912
rect 164770 165520 165570 165640
rect 0 162256 800 162376
rect 164770 161304 165570 161424
rect 0 158720 800 158840
rect 164770 157088 165570 157208
rect 0 155184 800 155304
rect 164770 152872 165570 152992
rect 0 151512 800 151632
rect 164770 148656 165570 148776
rect 0 147976 800 148096
rect 0 144440 800 144560
rect 164770 144576 165570 144696
rect 0 140904 800 141024
rect 164770 140360 165570 140480
rect 0 137232 800 137352
rect 164770 136144 165570 136264
rect 0 133696 800 133816
rect 164770 131928 165570 132048
rect 0 130160 800 130280
rect 164770 127712 165570 127832
rect 0 126624 800 126744
rect 164770 123496 165570 123616
rect 0 122952 800 123072
rect 0 119416 800 119536
rect 164770 119416 165570 119536
rect 0 115880 800 116000
rect 164770 115200 165570 115320
rect 0 112344 800 112464
rect 164770 110984 165570 111104
rect 0 108808 800 108928
rect 164770 106768 165570 106888
rect 0 105136 800 105256
rect 164770 102552 165570 102672
rect 0 101600 800 101720
rect 164770 98336 165570 98456
rect 0 98064 800 98184
rect 0 94528 800 94648
rect 164770 94256 165570 94376
rect 0 90856 800 90976
rect 164770 90040 165570 90160
rect 0 87320 800 87440
rect 164770 85824 165570 85944
rect 0 83784 800 83904
rect 164770 81608 165570 81728
rect 0 80248 800 80368
rect 164770 77392 165570 77512
rect 0 76576 800 76696
rect 164770 73312 165570 73432
rect 0 73040 800 73160
rect 0 69504 800 69624
rect 164770 69096 165570 69216
rect 0 65968 800 66088
rect 164770 64880 165570 65000
rect 0 62296 800 62416
rect 164770 60664 165570 60784
rect 0 58760 800 58880
rect 164770 56448 165570 56568
rect 0 55224 800 55344
rect 164770 52232 165570 52352
rect 0 51688 800 51808
rect 0 48152 800 48272
rect 164770 48152 165570 48272
rect 0 44480 800 44600
rect 164770 43936 165570 44056
rect 0 40944 800 41064
rect 164770 39720 165570 39840
rect 0 37408 800 37528
rect 164770 35504 165570 35624
rect 0 33872 800 33992
rect 164770 31288 165570 31408
rect 0 30200 800 30320
rect 164770 27072 165570 27192
rect 0 26664 800 26784
rect 0 23128 800 23248
rect 164770 22992 165570 23112
rect 0 19592 800 19712
rect 164770 18776 165570 18896
rect 0 15920 800 16040
rect 164770 14560 165570 14680
rect 0 12384 800 12504
rect 164770 10344 165570 10464
rect 0 8848 800 8968
rect 164770 6128 165570 6248
rect 0 5312 800 5432
rect 164770 2048 165570 2168
rect 0 1776 800 1896
<< obsm3 >>
rect 13 165992 165403 167653
rect 880 165720 165403 165992
rect 880 165712 164690 165720
rect 13 165440 164690 165712
rect 13 162456 165403 165440
rect 880 162176 165403 162456
rect 13 161504 165403 162176
rect 13 161224 164690 161504
rect 13 158920 165403 161224
rect 880 158640 165403 158920
rect 13 157288 165403 158640
rect 13 157008 164690 157288
rect 13 155384 165403 157008
rect 880 155104 165403 155384
rect 13 153072 165403 155104
rect 13 152792 164690 153072
rect 13 151712 165403 152792
rect 880 151432 165403 151712
rect 13 148856 165403 151432
rect 13 148576 164690 148856
rect 13 148176 165403 148576
rect 880 147896 165403 148176
rect 13 144776 165403 147896
rect 13 144640 164690 144776
rect 880 144496 164690 144640
rect 880 144360 165403 144496
rect 13 141104 165403 144360
rect 880 140824 165403 141104
rect 13 140560 165403 140824
rect 13 140280 164690 140560
rect 13 137432 165403 140280
rect 880 137152 165403 137432
rect 13 136344 165403 137152
rect 13 136064 164690 136344
rect 13 133896 165403 136064
rect 880 133616 165403 133896
rect 13 132128 165403 133616
rect 13 131848 164690 132128
rect 13 130360 165403 131848
rect 880 130080 165403 130360
rect 13 127912 165403 130080
rect 13 127632 164690 127912
rect 13 126824 165403 127632
rect 880 126544 165403 126824
rect 13 123696 165403 126544
rect 13 123416 164690 123696
rect 13 123152 165403 123416
rect 880 122872 165403 123152
rect 13 119616 165403 122872
rect 880 119336 164690 119616
rect 13 116080 165403 119336
rect 880 115800 165403 116080
rect 13 115400 165403 115800
rect 13 115120 164690 115400
rect 13 112544 165403 115120
rect 880 112264 165403 112544
rect 13 111184 165403 112264
rect 13 110904 164690 111184
rect 13 109008 165403 110904
rect 880 108728 165403 109008
rect 13 106968 165403 108728
rect 13 106688 164690 106968
rect 13 105336 165403 106688
rect 880 105056 165403 105336
rect 13 102752 165403 105056
rect 13 102472 164690 102752
rect 13 101800 165403 102472
rect 880 101520 165403 101800
rect 13 98536 165403 101520
rect 13 98264 164690 98536
rect 880 98256 164690 98264
rect 880 97984 165403 98256
rect 13 94728 165403 97984
rect 880 94456 165403 94728
rect 880 94448 164690 94456
rect 13 94176 164690 94448
rect 13 91056 165403 94176
rect 880 90776 165403 91056
rect 13 90240 165403 90776
rect 13 89960 164690 90240
rect 13 87520 165403 89960
rect 880 87240 165403 87520
rect 13 86024 165403 87240
rect 13 85744 164690 86024
rect 13 83984 165403 85744
rect 880 83704 165403 83984
rect 13 81808 165403 83704
rect 13 81528 164690 81808
rect 13 80448 165403 81528
rect 880 80168 165403 80448
rect 13 77592 165403 80168
rect 13 77312 164690 77592
rect 13 76776 165403 77312
rect 880 76496 165403 76776
rect 13 73512 165403 76496
rect 13 73240 164690 73512
rect 880 73232 164690 73240
rect 880 72960 165403 73232
rect 13 69704 165403 72960
rect 880 69424 165403 69704
rect 13 69296 165403 69424
rect 13 69016 164690 69296
rect 13 66168 165403 69016
rect 880 65888 165403 66168
rect 13 65080 165403 65888
rect 13 64800 164690 65080
rect 13 62496 165403 64800
rect 880 62216 165403 62496
rect 13 60864 165403 62216
rect 13 60584 164690 60864
rect 13 58960 165403 60584
rect 880 58680 165403 58960
rect 13 56648 165403 58680
rect 13 56368 164690 56648
rect 13 55424 165403 56368
rect 880 55144 165403 55424
rect 13 52432 165403 55144
rect 13 52152 164690 52432
rect 13 51888 165403 52152
rect 880 51608 165403 51888
rect 13 48352 165403 51608
rect 880 48072 164690 48352
rect 13 44680 165403 48072
rect 880 44400 165403 44680
rect 13 44136 165403 44400
rect 13 43856 164690 44136
rect 13 41144 165403 43856
rect 880 40864 165403 41144
rect 13 39920 165403 40864
rect 13 39640 164690 39920
rect 13 37608 165403 39640
rect 880 37328 165403 37608
rect 13 35704 165403 37328
rect 13 35424 164690 35704
rect 13 34072 165403 35424
rect 880 33792 165403 34072
rect 13 31488 165403 33792
rect 13 31208 164690 31488
rect 13 30400 165403 31208
rect 880 30120 165403 30400
rect 13 27272 165403 30120
rect 13 26992 164690 27272
rect 13 26864 165403 26992
rect 880 26584 165403 26864
rect 13 23328 165403 26584
rect 880 23192 165403 23328
rect 880 23048 164690 23192
rect 13 22912 164690 23048
rect 13 19792 165403 22912
rect 880 19512 165403 19792
rect 13 18976 165403 19512
rect 13 18696 164690 18976
rect 13 16120 165403 18696
rect 880 15840 165403 16120
rect 13 14760 165403 15840
rect 13 14480 164690 14760
rect 13 12584 165403 14480
rect 880 12304 165403 12584
rect 13 10544 165403 12304
rect 13 10264 164690 10544
rect 13 9048 165403 10264
rect 880 8768 165403 9048
rect 13 6328 165403 8768
rect 13 6048 164690 6328
rect 13 5512 165403 6048
rect 880 5232 165403 5512
rect 13 2248 165403 5232
rect 13 1976 164690 2248
rect 880 1968 164690 1976
rect 880 1803 165403 1968
<< metal4 >>
rect 4208 2128 4528 165424
rect 19568 2128 19888 165424
rect 34928 2128 35248 165424
rect 50288 2128 50608 165424
rect 65648 2128 65968 165424
rect 81008 2128 81328 165424
rect 96368 2128 96688 165424
rect 111728 2128 112048 165424
rect 127088 2128 127408 165424
rect 142448 2128 142768 165424
rect 157808 2128 158128 165424
<< obsm4 >>
rect 14227 165504 162781 167653
rect 14227 3027 19488 165504
rect 19968 3027 34848 165504
rect 35328 3027 50208 165504
rect 50688 3027 65568 165504
rect 66048 3027 80928 165504
rect 81408 3027 96288 165504
rect 96768 3027 111648 165504
rect 112128 3027 127008 165504
rect 127488 3027 142368 165504
rect 142848 3027 157728 165504
rect 158208 3027 162781 165504
<< labels >>
rlabel metal3 s 0 1776 800 1896 6 clk_i
port 1 nsew signal input
rlabel metal2 s 129738 0 129794 800 6 i_dout0[0]
port 2 nsew signal input
rlabel metal2 s 152002 0 152058 800 6 i_dout0[10]
port 3 nsew signal input
rlabel metal2 s 153198 0 153254 800 6 i_dout0[11]
port 4 nsew signal input
rlabel metal2 s 154394 0 154450 800 6 i_dout0[12]
port 5 nsew signal input
rlabel metal3 s 0 80248 800 80368 6 i_dout0[13]
port 6 nsew signal input
rlabel metal3 s 164770 77392 165570 77512 6 i_dout0[14]
port 7 nsew signal input
rlabel metal2 s 156694 0 156750 800 6 i_dout0[15]
port 8 nsew signal input
rlabel metal2 s 148966 166914 149022 167714 6 i_dout0[16]
port 9 nsew signal input
rlabel metal3 s 0 98064 800 98184 6 i_dout0[17]
port 10 nsew signal input
rlabel metal2 s 152186 166914 152242 167714 6 i_dout0[18]
port 11 nsew signal input
rlabel metal3 s 0 108808 800 108928 6 i_dout0[19]
port 12 nsew signal input
rlabel metal3 s 0 23128 800 23248 6 i_dout0[1]
port 13 nsew signal input
rlabel metal3 s 164770 106768 165570 106888 6 i_dout0[20]
port 14 nsew signal input
rlabel metal2 s 154302 166914 154358 167714 6 i_dout0[21]
port 15 nsew signal input
rlabel metal2 s 155314 166914 155370 167714 6 i_dout0[22]
port 16 nsew signal input
rlabel metal2 s 156418 166914 156474 167714 6 i_dout0[23]
port 17 nsew signal input
rlabel metal2 s 157522 166914 157578 167714 6 i_dout0[24]
port 18 nsew signal input
rlabel metal3 s 164770 127712 165570 127832 6 i_dout0[25]
port 19 nsew signal input
rlabel metal3 s 164770 131928 165570 132048 6 i_dout0[26]
port 20 nsew signal input
rlabel metal3 s 0 151512 800 151632 6 i_dout0[27]
port 21 nsew signal input
rlabel metal3 s 0 155184 800 155304 6 i_dout0[28]
port 22 nsew signal input
rlabel metal2 s 163778 0 163834 800 6 i_dout0[29]
port 23 nsew signal input
rlabel metal2 s 136730 0 136786 800 6 i_dout0[2]
port 24 nsew signal input
rlabel metal3 s 0 162256 800 162376 6 i_dout0[30]
port 25 nsew signal input
rlabel metal2 s 164974 0 165030 800 6 i_dout0[31]
port 26 nsew signal input
rlabel metal2 s 127530 166914 127586 167714 6 i_dout0[3]
port 27 nsew signal input
rlabel metal3 s 0 37408 800 37528 6 i_dout0[4]
port 28 nsew signal input
rlabel metal3 s 0 48152 800 48272 6 i_dout0[5]
port 29 nsew signal input
rlabel metal2 s 145010 0 145066 800 6 i_dout0[6]
port 30 nsew signal input
rlabel metal2 s 135074 166914 135130 167714 6 i_dout0[7]
port 31 nsew signal input
rlabel metal2 s 138294 166914 138350 167714 6 i_dout0[8]
port 32 nsew signal input
rlabel metal2 s 149702 0 149758 800 6 i_dout0[9]
port 33 nsew signal input
rlabel metal3 s 164770 6128 165570 6248 6 i_dout0_1[0]
port 34 nsew signal input
rlabel metal2 s 150898 0 150954 800 6 i_dout0_1[10]
port 35 nsew signal input
rlabel metal2 s 143630 166914 143686 167714 6 i_dout0_1[11]
port 36 nsew signal input
rlabel metal2 s 144642 166914 144698 167714 6 i_dout0_1[12]
port 37 nsew signal input
rlabel metal2 s 145746 166914 145802 167714 6 i_dout0_1[13]
port 38 nsew signal input
rlabel metal2 s 147862 166914 147918 167714 6 i_dout0_1[14]
port 39 nsew signal input
rlabel metal2 s 155590 0 155646 800 6 i_dout0_1[15]
port 40 nsew signal input
rlabel metal3 s 0 90856 800 90976 6 i_dout0_1[16]
port 41 nsew signal input
rlabel metal3 s 0 94528 800 94648 6 i_dout0_1[17]
port 42 nsew signal input
rlabel metal3 s 0 105136 800 105256 6 i_dout0_1[18]
port 43 nsew signal input
rlabel metal3 s 164770 94256 165570 94376 6 i_dout0_1[19]
port 44 nsew signal input
rlabel metal3 s 0 19592 800 19712 6 i_dout0_1[1]
port 45 nsew signal input
rlabel metal3 s 164770 102552 165570 102672 6 i_dout0_1[20]
port 46 nsew signal input
rlabel metal2 s 161386 0 161442 800 6 i_dout0_1[21]
port 47 nsew signal input
rlabel metal3 s 0 119416 800 119536 6 i_dout0_1[22]
port 48 nsew signal input
rlabel metal3 s 0 122952 800 123072 6 i_dout0_1[23]
port 49 nsew signal input
rlabel metal3 s 0 130160 800 130280 6 i_dout0_1[24]
port 50 nsew signal input
rlabel metal3 s 164770 123496 165570 123616 6 i_dout0_1[25]
port 51 nsew signal input
rlabel metal2 s 160650 166914 160706 167714 6 i_dout0_1[26]
port 52 nsew signal input
rlabel metal3 s 0 147976 800 148096 6 i_dout0_1[27]
port 53 nsew signal input
rlabel metal3 s 164770 136144 165570 136264 6 i_dout0_1[28]
port 54 nsew signal input
rlabel metal2 s 164974 166914 165030 167714 6 i_dout0_1[29]
port 55 nsew signal input
rlabel metal3 s 164770 22992 165570 23112 6 i_dout0_1[2]
port 56 nsew signal input
rlabel metal3 s 164770 148656 165570 148776 6 i_dout0_1[30]
port 57 nsew signal input
rlabel metal3 s 164770 161304 165570 161424 6 i_dout0_1[31]
port 58 nsew signal input
rlabel metal3 s 0 30200 800 30320 6 i_dout0_1[3]
port 59 nsew signal input
rlabel metal3 s 164770 35504 165570 35624 6 i_dout0_1[4]
port 60 nsew signal input
rlabel metal3 s 0 44480 800 44600 6 i_dout0_1[5]
port 61 nsew signal input
rlabel metal3 s 164770 48152 165570 48272 6 i_dout0_1[6]
port 62 nsew signal input
rlabel metal2 s 133970 166914 134026 167714 6 i_dout0_1[7]
port 63 nsew signal input
rlabel metal2 s 148506 0 148562 800 6 i_dout0_1[8]
port 64 nsew signal input
rlabel metal2 s 140410 166914 140466 167714 6 i_dout0_1[9]
port 65 nsew signal input
rlabel metal2 s 478 166914 534 167714 6 io_in[0]
port 66 nsew signal input
rlabel metal2 s 32494 166914 32550 167714 6 io_in[10]
port 67 nsew signal input
rlabel metal2 s 35714 166914 35770 167714 6 io_in[11]
port 68 nsew signal input
rlabel metal2 s 38934 166914 38990 167714 6 io_in[12]
port 69 nsew signal input
rlabel metal2 s 42062 166914 42118 167714 6 io_in[13]
port 70 nsew signal input
rlabel metal2 s 45282 166914 45338 167714 6 io_in[14]
port 71 nsew signal input
rlabel metal2 s 48502 166914 48558 167714 6 io_in[15]
port 72 nsew signal input
rlabel metal2 s 51722 166914 51778 167714 6 io_in[16]
port 73 nsew signal input
rlabel metal2 s 54942 166914 54998 167714 6 io_in[17]
port 74 nsew signal input
rlabel metal2 s 58162 166914 58218 167714 6 io_in[18]
port 75 nsew signal input
rlabel metal2 s 61290 166914 61346 167714 6 io_in[19]
port 76 nsew signal input
rlabel metal2 s 3606 166914 3662 167714 6 io_in[1]
port 77 nsew signal input
rlabel metal2 s 64510 166914 64566 167714 6 io_in[20]
port 78 nsew signal input
rlabel metal2 s 67730 166914 67786 167714 6 io_in[21]
port 79 nsew signal input
rlabel metal2 s 70950 166914 71006 167714 6 io_in[22]
port 80 nsew signal input
rlabel metal2 s 74170 166914 74226 167714 6 io_in[23]
port 81 nsew signal input
rlabel metal2 s 77390 166914 77446 167714 6 io_in[24]
port 82 nsew signal input
rlabel metal2 s 80518 166914 80574 167714 6 io_in[25]
port 83 nsew signal input
rlabel metal2 s 83738 166914 83794 167714 6 io_in[26]
port 84 nsew signal input
rlabel metal2 s 86958 166914 87014 167714 6 io_in[27]
port 85 nsew signal input
rlabel metal2 s 90178 166914 90234 167714 6 io_in[28]
port 86 nsew signal input
rlabel metal2 s 93398 166914 93454 167714 6 io_in[29]
port 87 nsew signal input
rlabel metal2 s 6826 166914 6882 167714 6 io_in[2]
port 88 nsew signal input
rlabel metal2 s 96618 166914 96674 167714 6 io_in[30]
port 89 nsew signal input
rlabel metal2 s 99838 166914 99894 167714 6 io_in[31]
port 90 nsew signal input
rlabel metal2 s 102966 166914 103022 167714 6 io_in[32]
port 91 nsew signal input
rlabel metal2 s 106186 166914 106242 167714 6 io_in[33]
port 92 nsew signal input
rlabel metal2 s 109406 166914 109462 167714 6 io_in[34]
port 93 nsew signal input
rlabel metal2 s 112626 166914 112682 167714 6 io_in[35]
port 94 nsew signal input
rlabel metal2 s 115846 166914 115902 167714 6 io_in[36]
port 95 nsew signal input
rlabel metal2 s 119066 166914 119122 167714 6 io_in[37]
port 96 nsew signal input
rlabel metal2 s 10046 166914 10102 167714 6 io_in[3]
port 97 nsew signal input
rlabel metal2 s 13266 166914 13322 167714 6 io_in[4]
port 98 nsew signal input
rlabel metal2 s 16486 166914 16542 167714 6 io_in[5]
port 99 nsew signal input
rlabel metal2 s 19706 166914 19762 167714 6 io_in[6]
port 100 nsew signal input
rlabel metal2 s 22834 166914 22890 167714 6 io_in[7]
port 101 nsew signal input
rlabel metal2 s 26054 166914 26110 167714 6 io_in[8]
port 102 nsew signal input
rlabel metal2 s 29274 166914 29330 167714 6 io_in[9]
port 103 nsew signal input
rlabel metal2 s 1490 166914 1546 167714 6 io_oeb[0]
port 104 nsew signal output
rlabel metal2 s 33598 166914 33654 167714 6 io_oeb[10]
port 105 nsew signal output
rlabel metal2 s 36726 166914 36782 167714 6 io_oeb[11]
port 106 nsew signal output
rlabel metal2 s 39946 166914 40002 167714 6 io_oeb[12]
port 107 nsew signal output
rlabel metal2 s 43166 166914 43222 167714 6 io_oeb[13]
port 108 nsew signal output
rlabel metal2 s 46386 166914 46442 167714 6 io_oeb[14]
port 109 nsew signal output
rlabel metal2 s 49606 166914 49662 167714 6 io_oeb[15]
port 110 nsew signal output
rlabel metal2 s 52826 166914 52882 167714 6 io_oeb[16]
port 111 nsew signal output
rlabel metal2 s 55954 166914 56010 167714 6 io_oeb[17]
port 112 nsew signal output
rlabel metal2 s 59174 166914 59230 167714 6 io_oeb[18]
port 113 nsew signal output
rlabel metal2 s 62394 166914 62450 167714 6 io_oeb[19]
port 114 nsew signal output
rlabel metal2 s 4710 166914 4766 167714 6 io_oeb[1]
port 115 nsew signal output
rlabel metal2 s 65614 166914 65670 167714 6 io_oeb[20]
port 116 nsew signal output
rlabel metal2 s 68834 166914 68890 167714 6 io_oeb[21]
port 117 nsew signal output
rlabel metal2 s 72054 166914 72110 167714 6 io_oeb[22]
port 118 nsew signal output
rlabel metal2 s 75182 166914 75238 167714 6 io_oeb[23]
port 119 nsew signal output
rlabel metal2 s 78402 166914 78458 167714 6 io_oeb[24]
port 120 nsew signal output
rlabel metal2 s 81622 166914 81678 167714 6 io_oeb[25]
port 121 nsew signal output
rlabel metal2 s 84842 166914 84898 167714 6 io_oeb[26]
port 122 nsew signal output
rlabel metal2 s 88062 166914 88118 167714 6 io_oeb[27]
port 123 nsew signal output
rlabel metal2 s 91282 166914 91338 167714 6 io_oeb[28]
port 124 nsew signal output
rlabel metal2 s 94410 166914 94466 167714 6 io_oeb[29]
port 125 nsew signal output
rlabel metal2 s 7930 166914 7986 167714 6 io_oeb[2]
port 126 nsew signal output
rlabel metal2 s 97630 166914 97686 167714 6 io_oeb[30]
port 127 nsew signal output
rlabel metal2 s 100850 166914 100906 167714 6 io_oeb[31]
port 128 nsew signal output
rlabel metal2 s 104070 166914 104126 167714 6 io_oeb[32]
port 129 nsew signal output
rlabel metal2 s 107290 166914 107346 167714 6 io_oeb[33]
port 130 nsew signal output
rlabel metal2 s 110510 166914 110566 167714 6 io_oeb[34]
port 131 nsew signal output
rlabel metal2 s 113638 166914 113694 167714 6 io_oeb[35]
port 132 nsew signal output
rlabel metal2 s 116858 166914 116914 167714 6 io_oeb[36]
port 133 nsew signal output
rlabel metal2 s 120078 166914 120134 167714 6 io_oeb[37]
port 134 nsew signal output
rlabel metal2 s 11150 166914 11206 167714 6 io_oeb[3]
port 135 nsew signal output
rlabel metal2 s 14278 166914 14334 167714 6 io_oeb[4]
port 136 nsew signal output
rlabel metal2 s 17498 166914 17554 167714 6 io_oeb[5]
port 137 nsew signal output
rlabel metal2 s 20718 166914 20774 167714 6 io_oeb[6]
port 138 nsew signal output
rlabel metal2 s 23938 166914 23994 167714 6 io_oeb[7]
port 139 nsew signal output
rlabel metal2 s 27158 166914 27214 167714 6 io_oeb[8]
port 140 nsew signal output
rlabel metal2 s 30378 166914 30434 167714 6 io_oeb[9]
port 141 nsew signal output
rlabel metal2 s 2594 166914 2650 167714 6 io_out[0]
port 142 nsew signal output
rlabel metal2 s 34610 166914 34666 167714 6 io_out[10]
port 143 nsew signal output
rlabel metal2 s 37830 166914 37886 167714 6 io_out[11]
port 144 nsew signal output
rlabel metal2 s 41050 166914 41106 167714 6 io_out[12]
port 145 nsew signal output
rlabel metal2 s 44270 166914 44326 167714 6 io_out[13]
port 146 nsew signal output
rlabel metal2 s 47398 166914 47454 167714 6 io_out[14]
port 147 nsew signal output
rlabel metal2 s 50618 166914 50674 167714 6 io_out[15]
port 148 nsew signal output
rlabel metal2 s 53838 166914 53894 167714 6 io_out[16]
port 149 nsew signal output
rlabel metal2 s 57058 166914 57114 167714 6 io_out[17]
port 150 nsew signal output
rlabel metal2 s 60278 166914 60334 167714 6 io_out[18]
port 151 nsew signal output
rlabel metal2 s 63498 166914 63554 167714 6 io_out[19]
port 152 nsew signal output
rlabel metal2 s 5814 166914 5870 167714 6 io_out[1]
port 153 nsew signal output
rlabel metal2 s 66718 166914 66774 167714 6 io_out[20]
port 154 nsew signal output
rlabel metal2 s 69846 166914 69902 167714 6 io_out[21]
port 155 nsew signal output
rlabel metal2 s 73066 166914 73122 167714 6 io_out[22]
port 156 nsew signal output
rlabel metal2 s 76286 166914 76342 167714 6 io_out[23]
port 157 nsew signal output
rlabel metal2 s 79506 166914 79562 167714 6 io_out[24]
port 158 nsew signal output
rlabel metal2 s 82726 166914 82782 167714 6 io_out[25]
port 159 nsew signal output
rlabel metal2 s 85946 166914 86002 167714 6 io_out[26]
port 160 nsew signal output
rlabel metal2 s 89074 166914 89130 167714 6 io_out[27]
port 161 nsew signal output
rlabel metal2 s 92294 166914 92350 167714 6 io_out[28]
port 162 nsew signal output
rlabel metal2 s 95514 166914 95570 167714 6 io_out[29]
port 163 nsew signal output
rlabel metal2 s 8942 166914 8998 167714 6 io_out[2]
port 164 nsew signal output
rlabel metal2 s 98734 166914 98790 167714 6 io_out[30]
port 165 nsew signal output
rlabel metal2 s 101954 166914 102010 167714 6 io_out[31]
port 166 nsew signal output
rlabel metal2 s 105174 166914 105230 167714 6 io_out[32]
port 167 nsew signal output
rlabel metal2 s 108302 166914 108358 167714 6 io_out[33]
port 168 nsew signal output
rlabel metal2 s 111522 166914 111578 167714 6 io_out[34]
port 169 nsew signal output
rlabel metal2 s 114742 166914 114798 167714 6 io_out[35]
port 170 nsew signal output
rlabel metal2 s 117962 166914 118018 167714 6 io_out[36]
port 171 nsew signal output
rlabel metal2 s 121182 166914 121238 167714 6 io_out[37]
port 172 nsew signal output
rlabel metal2 s 12162 166914 12218 167714 6 io_out[3]
port 173 nsew signal output
rlabel metal2 s 15382 166914 15438 167714 6 io_out[4]
port 174 nsew signal output
rlabel metal2 s 18602 166914 18658 167714 6 io_out[5]
port 175 nsew signal output
rlabel metal2 s 21822 166914 21878 167714 6 io_out[6]
port 176 nsew signal output
rlabel metal2 s 25042 166914 25098 167714 6 io_out[7]
port 177 nsew signal output
rlabel metal2 s 28170 166914 28226 167714 6 io_out[8]
port 178 nsew signal output
rlabel metal2 s 31390 166914 31446 167714 6 io_out[9]
port 179 nsew signal output
rlabel metal2 s 125046 0 125102 800 6 irq[0]
port 180 nsew signal output
rlabel metal2 s 126150 0 126206 800 6 irq[1]
port 181 nsew signal output
rlabel metal2 s 127346 0 127402 800 6 irq[2]
port 182 nsew signal output
rlabel metal3 s 0 5312 800 5432 6 o_csb0
port 183 nsew signal output
rlabel metal2 s 128542 0 128598 800 6 o_csb0_1
port 184 nsew signal output
rlabel metal2 s 123298 166914 123354 167714 6 o_din0[0]
port 185 nsew signal output
rlabel metal3 s 164770 60664 165570 60784 6 o_din0[10]
port 186 nsew signal output
rlabel metal3 s 0 73040 800 73160 6 o_din0[11]
port 187 nsew signal output
rlabel metal3 s 0 76576 800 76696 6 o_din0[12]
port 188 nsew signal output
rlabel metal3 s 164770 73312 165570 73432 6 o_din0[13]
port 189 nsew signal output
rlabel metal3 s 164770 81608 165570 81728 6 o_din0[14]
port 190 nsew signal output
rlabel metal3 s 0 87320 800 87440 6 o_din0[15]
port 191 nsew signal output
rlabel metal2 s 151082 166914 151138 167714 6 o_din0[16]
port 192 nsew signal output
rlabel metal2 s 157890 0 157946 800 6 o_din0[17]
port 193 nsew signal output
rlabel metal3 s 164770 90040 165570 90160 6 o_din0[18]
port 194 nsew signal output
rlabel metal3 s 164770 98336 165570 98456 6 o_din0[19]
port 195 nsew signal output
rlabel metal3 s 164770 14560 165570 14680 6 o_din0[1]
port 196 nsew signal output
rlabel metal3 s 164770 110984 165570 111104 6 o_din0[20]
port 197 nsew signal output
rlabel metal3 s 0 115880 800 116000 6 o_din0[21]
port 198 nsew signal output
rlabel metal2 s 162582 0 162638 800 6 o_din0[22]
port 199 nsew signal output
rlabel metal3 s 0 126624 800 126744 6 o_din0[23]
port 200 nsew signal output
rlabel metal2 s 158534 166914 158590 167714 6 o_din0[24]
port 201 nsew signal output
rlabel metal2 s 159638 166914 159694 167714 6 o_din0[25]
port 202 nsew signal output
rlabel metal3 s 0 144440 800 144560 6 o_din0[26]
port 203 nsew signal output
rlabel metal2 s 162858 166914 162914 167714 6 o_din0[27]
port 204 nsew signal output
rlabel metal3 s 164770 140360 165570 140480 6 o_din0[28]
port 205 nsew signal output
rlabel metal3 s 164770 144576 165570 144696 6 o_din0[29]
port 206 nsew signal output
rlabel metal2 s 137926 0 137982 800 6 o_din0[2]
port 207 nsew signal output
rlabel metal3 s 164770 157088 165570 157208 6 o_din0[30]
port 208 nsew signal output
rlabel metal3 s 0 165792 800 165912 6 o_din0[31]
port 209 nsew signal output
rlabel metal2 s 141422 0 141478 800 6 o_din0[3]
port 210 nsew signal output
rlabel metal3 s 0 40944 800 41064 6 o_din0[4]
port 211 nsew signal output
rlabel metal3 s 0 51688 800 51808 6 o_din0[5]
port 212 nsew signal output
rlabel metal2 s 131854 166914 131910 167714 6 o_din0[6]
port 213 nsew signal output
rlabel metal2 s 136086 166914 136142 167714 6 o_din0[7]
port 214 nsew signal output
rlabel metal3 s 0 65968 800 66088 6 o_din0[8]
port 215 nsew signal output
rlabel metal2 s 141422 166914 141478 167714 6 o_din0[9]
port 216 nsew signal output
rlabel metal3 s 164770 10344 165570 10464 6 o_din0_1[0]
port 217 nsew signal output
rlabel metal2 s 142526 166914 142582 167714 6 o_din0_1[10]
port 218 nsew signal output
rlabel metal3 s 164770 64880 165570 65000 6 o_din0_1[11]
port 219 nsew signal output
rlabel metal3 s 164770 69096 165570 69216 6 o_din0_1[12]
port 220 nsew signal output
rlabel metal2 s 146758 166914 146814 167714 6 o_din0_1[13]
port 221 nsew signal output
rlabel metal3 s 0 83784 800 83904 6 o_din0_1[14]
port 222 nsew signal output
rlabel metal3 s 164770 85824 165570 85944 6 o_din0_1[15]
port 223 nsew signal output
rlabel metal2 s 149978 166914 150034 167714 6 o_din0_1[16]
port 224 nsew signal output
rlabel metal3 s 0 101600 800 101720 6 o_din0_1[17]
port 225 nsew signal output
rlabel metal2 s 159086 0 159142 800 6 o_din0_1[18]
port 226 nsew signal output
rlabel metal2 s 160282 0 160338 800 6 o_din0_1[19]
port 227 nsew signal output
rlabel metal3 s 0 26664 800 26784 6 o_din0_1[1]
port 228 nsew signal output
rlabel metal2 s 153198 166914 153254 167714 6 o_din0_1[20]
port 229 nsew signal output
rlabel metal3 s 0 112344 800 112464 6 o_din0_1[21]
port 230 nsew signal output
rlabel metal3 s 164770 115200 165570 115320 6 o_din0_1[22]
port 231 nsew signal output
rlabel metal3 s 164770 119416 165570 119536 6 o_din0_1[23]
port 232 nsew signal output
rlabel metal3 s 0 133696 800 133816 6 o_din0_1[24]
port 233 nsew signal output
rlabel metal3 s 0 137232 800 137352 6 o_din0_1[25]
port 234 nsew signal output
rlabel metal3 s 0 140904 800 141024 6 o_din0_1[26]
port 235 nsew signal output
rlabel metal2 s 161754 166914 161810 167714 6 o_din0_1[27]
port 236 nsew signal output
rlabel metal2 s 163870 166914 163926 167714 6 o_din0_1[28]
port 237 nsew signal output
rlabel metal3 s 0 158720 800 158840 6 o_din0_1[29]
port 238 nsew signal output
rlabel metal2 s 124402 166914 124458 167714 6 o_din0_1[2]
port 239 nsew signal output
rlabel metal3 s 164770 152872 165570 152992 6 o_din0_1[30]
port 240 nsew signal output
rlabel metal3 s 164770 165520 165570 165640 6 o_din0_1[31]
port 241 nsew signal output
rlabel metal3 s 164770 27072 165570 27192 6 o_din0_1[3]
port 242 nsew signal output
rlabel metal2 s 143814 0 143870 800 6 o_din0_1[4]
port 243 nsew signal output
rlabel metal2 s 129738 166914 129794 167714 6 o_din0_1[5]
port 244 nsew signal output
rlabel metal2 s 130750 166914 130806 167714 6 o_din0_1[6]
port 245 nsew signal output
rlabel metal2 s 146114 0 146170 800 6 o_din0_1[7]
port 246 nsew signal output
rlabel metal3 s 0 62296 800 62416 6 o_din0_1[8]
port 247 nsew signal output
rlabel metal3 s 164770 56448 165570 56568 6 o_din0_1[9]
port 248 nsew signal output
rlabel metal3 s 0 12384 800 12504 6 o_waddr0[0]
port 249 nsew signal output
rlabel metal2 s 133234 0 133290 800 6 o_waddr0[1]
port 250 nsew signal output
rlabel metal2 s 139122 0 139178 800 6 o_waddr0[2]
port 251 nsew signal output
rlabel metal2 s 142618 0 142674 800 6 o_waddr0[3]
port 252 nsew signal output
rlabel metal3 s 164770 43936 165570 44056 6 o_waddr0[4]
port 253 nsew signal output
rlabel metal3 s 0 58760 800 58880 6 o_waddr0[5]
port 254 nsew signal output
rlabel metal2 s 132958 166914 133014 167714 6 o_waddr0[6]
port 255 nsew signal output
rlabel metal2 s 137190 166914 137246 167714 6 o_waddr0[7]
port 256 nsew signal output
rlabel metal3 s 0 69504 800 69624 6 o_waddr0[8]
port 257 nsew signal output
rlabel metal3 s 0 15920 800 16040 6 o_waddr0_1[0]
port 258 nsew signal output
rlabel metal3 s 164770 18776 165570 18896 6 o_waddr0_1[1]
port 259 nsew signal output
rlabel metal2 s 125414 166914 125470 167714 6 o_waddr0_1[2]
port 260 nsew signal output
rlabel metal3 s 164770 31288 165570 31408 6 o_waddr0_1[3]
port 261 nsew signal output
rlabel metal3 s 164770 39720 165570 39840 6 o_waddr0_1[4]
port 262 nsew signal output
rlabel metal3 s 0 55224 800 55344 6 o_waddr0_1[5]
port 263 nsew signal output
rlabel metal3 s 164770 52232 165570 52352 6 o_waddr0_1[6]
port 264 nsew signal output
rlabel metal2 s 147310 0 147366 800 6 o_waddr0_1[7]
port 265 nsew signal output
rlabel metal2 s 139306 166914 139362 167714 6 o_waddr0_1[8]
port 266 nsew signal output
rlabel metal2 s 122194 166914 122250 167714 6 o_web0
port 267 nsew signal output
rlabel metal3 s 0 8848 800 8968 6 o_web0_1
port 268 nsew signal output
rlabel metal2 s 130934 0 130990 800 6 o_wmask0[0]
port 269 nsew signal output
rlabel metal2 s 135626 0 135682 800 6 o_wmask0[1]
port 270 nsew signal output
rlabel metal2 s 126518 166914 126574 167714 6 o_wmask0[2]
port 271 nsew signal output
rlabel metal3 s 0 33872 800 33992 6 o_wmask0[3]
port 272 nsew signal output
rlabel metal2 s 132038 0 132094 800 6 o_wmask0_1[0]
port 273 nsew signal output
rlabel metal2 s 134430 0 134486 800 6 o_wmask0_1[1]
port 274 nsew signal output
rlabel metal2 s 140318 0 140374 800 6 o_wmask0_1[2]
port 275 nsew signal output
rlabel metal2 s 128634 166914 128690 167714 6 o_wmask0_1[3]
port 276 nsew signal output
rlabel metal3 s 164770 2048 165570 2168 6 rst_i
port 277 nsew signal input
rlabel metal4 s 4208 2128 4528 165424 6 vccd1
port 278 nsew power input
rlabel metal4 s 34928 2128 35248 165424 6 vccd1
port 278 nsew power input
rlabel metal4 s 65648 2128 65968 165424 6 vccd1
port 278 nsew power input
rlabel metal4 s 96368 2128 96688 165424 6 vccd1
port 278 nsew power input
rlabel metal4 s 127088 2128 127408 165424 6 vccd1
port 278 nsew power input
rlabel metal4 s 157808 2128 158128 165424 6 vccd1
port 278 nsew power input
rlabel metal4 s 19568 2128 19888 165424 6 vssd1
port 279 nsew ground input
rlabel metal4 s 50288 2128 50608 165424 6 vssd1
port 279 nsew ground input
rlabel metal4 s 81008 2128 81328 165424 6 vssd1
port 279 nsew ground input
rlabel metal4 s 111728 2128 112048 165424 6 vssd1
port 279 nsew ground input
rlabel metal4 s 142448 2128 142768 165424 6 vssd1
port 279 nsew ground input
rlabel metal2 s 570 0 626 800 6 wb_clk_i
port 280 nsew signal input
rlabel metal2 s 1674 0 1730 800 6 wb_rst_i
port 281 nsew signal input
rlabel metal2 s 2870 0 2926 800 6 wbs_ack_o
port 282 nsew signal output
rlabel metal2 s 7562 0 7618 800 6 wbs_adr_i[0]
port 283 nsew signal input
rlabel metal2 s 47490 0 47546 800 6 wbs_adr_i[10]
port 284 nsew signal input
rlabel metal2 s 50986 0 51042 800 6 wbs_adr_i[11]
port 285 nsew signal input
rlabel metal2 s 54574 0 54630 800 6 wbs_adr_i[12]
port 286 nsew signal input
rlabel metal2 s 58070 0 58126 800 6 wbs_adr_i[13]
port 287 nsew signal input
rlabel metal2 s 61566 0 61622 800 6 wbs_adr_i[14]
port 288 nsew signal input
rlabel metal2 s 65154 0 65210 800 6 wbs_adr_i[15]
port 289 nsew signal input
rlabel metal2 s 68650 0 68706 800 6 wbs_adr_i[16]
port 290 nsew signal input
rlabel metal2 s 72146 0 72202 800 6 wbs_adr_i[17]
port 291 nsew signal input
rlabel metal2 s 75734 0 75790 800 6 wbs_adr_i[18]
port 292 nsew signal input
rlabel metal2 s 79230 0 79286 800 6 wbs_adr_i[19]
port 293 nsew signal input
rlabel metal2 s 12254 0 12310 800 6 wbs_adr_i[1]
port 294 nsew signal input
rlabel metal2 s 82726 0 82782 800 6 wbs_adr_i[20]
port 295 nsew signal input
rlabel metal2 s 86222 0 86278 800 6 wbs_adr_i[21]
port 296 nsew signal input
rlabel metal2 s 89810 0 89866 800 6 wbs_adr_i[22]
port 297 nsew signal input
rlabel metal2 s 93306 0 93362 800 6 wbs_adr_i[23]
port 298 nsew signal input
rlabel metal2 s 96802 0 96858 800 6 wbs_adr_i[24]
port 299 nsew signal input
rlabel metal2 s 100390 0 100446 800 6 wbs_adr_i[25]
port 300 nsew signal input
rlabel metal2 s 103886 0 103942 800 6 wbs_adr_i[26]
port 301 nsew signal input
rlabel metal2 s 107382 0 107438 800 6 wbs_adr_i[27]
port 302 nsew signal input
rlabel metal2 s 110970 0 111026 800 6 wbs_adr_i[28]
port 303 nsew signal input
rlabel metal2 s 114466 0 114522 800 6 wbs_adr_i[29]
port 304 nsew signal input
rlabel metal2 s 16946 0 17002 800 6 wbs_adr_i[2]
port 305 nsew signal input
rlabel metal2 s 117962 0 118018 800 6 wbs_adr_i[30]
port 306 nsew signal input
rlabel metal2 s 121458 0 121514 800 6 wbs_adr_i[31]
port 307 nsew signal input
rlabel metal2 s 21638 0 21694 800 6 wbs_adr_i[3]
port 308 nsew signal input
rlabel metal2 s 26330 0 26386 800 6 wbs_adr_i[4]
port 309 nsew signal input
rlabel metal2 s 29918 0 29974 800 6 wbs_adr_i[5]
port 310 nsew signal input
rlabel metal2 s 33414 0 33470 800 6 wbs_adr_i[6]
port 311 nsew signal input
rlabel metal2 s 36910 0 36966 800 6 wbs_adr_i[7]
port 312 nsew signal input
rlabel metal2 s 40498 0 40554 800 6 wbs_adr_i[8]
port 313 nsew signal input
rlabel metal2 s 43994 0 44050 800 6 wbs_adr_i[9]
port 314 nsew signal input
rlabel metal2 s 4066 0 4122 800 6 wbs_cyc_i
port 315 nsew signal input
rlabel metal2 s 8758 0 8814 800 6 wbs_dat_i[0]
port 316 nsew signal input
rlabel metal2 s 48686 0 48742 800 6 wbs_dat_i[10]
port 317 nsew signal input
rlabel metal2 s 52182 0 52238 800 6 wbs_dat_i[11]
port 318 nsew signal input
rlabel metal2 s 55770 0 55826 800 6 wbs_dat_i[12]
port 319 nsew signal input
rlabel metal2 s 59266 0 59322 800 6 wbs_dat_i[13]
port 320 nsew signal input
rlabel metal2 s 62762 0 62818 800 6 wbs_dat_i[14]
port 321 nsew signal input
rlabel metal2 s 66258 0 66314 800 6 wbs_dat_i[15]
port 322 nsew signal input
rlabel metal2 s 69846 0 69902 800 6 wbs_dat_i[16]
port 323 nsew signal input
rlabel metal2 s 73342 0 73398 800 6 wbs_dat_i[17]
port 324 nsew signal input
rlabel metal2 s 76838 0 76894 800 6 wbs_dat_i[18]
port 325 nsew signal input
rlabel metal2 s 80426 0 80482 800 6 wbs_dat_i[19]
port 326 nsew signal input
rlabel metal2 s 13450 0 13506 800 6 wbs_dat_i[1]
port 327 nsew signal input
rlabel metal2 s 83922 0 83978 800 6 wbs_dat_i[20]
port 328 nsew signal input
rlabel metal2 s 87418 0 87474 800 6 wbs_dat_i[21]
port 329 nsew signal input
rlabel metal2 s 90914 0 90970 800 6 wbs_dat_i[22]
port 330 nsew signal input
rlabel metal2 s 94502 0 94558 800 6 wbs_dat_i[23]
port 331 nsew signal input
rlabel metal2 s 97998 0 98054 800 6 wbs_dat_i[24]
port 332 nsew signal input
rlabel metal2 s 101494 0 101550 800 6 wbs_dat_i[25]
port 333 nsew signal input
rlabel metal2 s 105082 0 105138 800 6 wbs_dat_i[26]
port 334 nsew signal input
rlabel metal2 s 108578 0 108634 800 6 wbs_dat_i[27]
port 335 nsew signal input
rlabel metal2 s 112074 0 112130 800 6 wbs_dat_i[28]
port 336 nsew signal input
rlabel metal2 s 115662 0 115718 800 6 wbs_dat_i[29]
port 337 nsew signal input
rlabel metal2 s 18142 0 18198 800 6 wbs_dat_i[2]
port 338 nsew signal input
rlabel metal2 s 119158 0 119214 800 6 wbs_dat_i[30]
port 339 nsew signal input
rlabel metal2 s 122654 0 122710 800 6 wbs_dat_i[31]
port 340 nsew signal input
rlabel metal2 s 22834 0 22890 800 6 wbs_dat_i[3]
port 341 nsew signal input
rlabel metal2 s 27526 0 27582 800 6 wbs_dat_i[4]
port 342 nsew signal input
rlabel metal2 s 31022 0 31078 800 6 wbs_dat_i[5]
port 343 nsew signal input
rlabel metal2 s 34610 0 34666 800 6 wbs_dat_i[6]
port 344 nsew signal input
rlabel metal2 s 38106 0 38162 800 6 wbs_dat_i[7]
port 345 nsew signal input
rlabel metal2 s 41602 0 41658 800 6 wbs_dat_i[8]
port 346 nsew signal input
rlabel metal2 s 45190 0 45246 800 6 wbs_dat_i[9]
port 347 nsew signal input
rlabel metal2 s 9954 0 10010 800 6 wbs_dat_o[0]
port 348 nsew signal output
rlabel metal2 s 49882 0 49938 800 6 wbs_dat_o[10]
port 349 nsew signal output
rlabel metal2 s 53378 0 53434 800 6 wbs_dat_o[11]
port 350 nsew signal output
rlabel metal2 s 56874 0 56930 800 6 wbs_dat_o[12]
port 351 nsew signal output
rlabel metal2 s 60462 0 60518 800 6 wbs_dat_o[13]
port 352 nsew signal output
rlabel metal2 s 63958 0 64014 800 6 wbs_dat_o[14]
port 353 nsew signal output
rlabel metal2 s 67454 0 67510 800 6 wbs_dat_o[15]
port 354 nsew signal output
rlabel metal2 s 70950 0 71006 800 6 wbs_dat_o[16]
port 355 nsew signal output
rlabel metal2 s 74538 0 74594 800 6 wbs_dat_o[17]
port 356 nsew signal output
rlabel metal2 s 78034 0 78090 800 6 wbs_dat_o[18]
port 357 nsew signal output
rlabel metal2 s 81530 0 81586 800 6 wbs_dat_o[19]
port 358 nsew signal output
rlabel metal2 s 14646 0 14702 800 6 wbs_dat_o[1]
port 359 nsew signal output
rlabel metal2 s 85118 0 85174 800 6 wbs_dat_o[20]
port 360 nsew signal output
rlabel metal2 s 88614 0 88670 800 6 wbs_dat_o[21]
port 361 nsew signal output
rlabel metal2 s 92110 0 92166 800 6 wbs_dat_o[22]
port 362 nsew signal output
rlabel metal2 s 95698 0 95754 800 6 wbs_dat_o[23]
port 363 nsew signal output
rlabel metal2 s 99194 0 99250 800 6 wbs_dat_o[24]
port 364 nsew signal output
rlabel metal2 s 102690 0 102746 800 6 wbs_dat_o[25]
port 365 nsew signal output
rlabel metal2 s 106186 0 106242 800 6 wbs_dat_o[26]
port 366 nsew signal output
rlabel metal2 s 109774 0 109830 800 6 wbs_dat_o[27]
port 367 nsew signal output
rlabel metal2 s 113270 0 113326 800 6 wbs_dat_o[28]
port 368 nsew signal output
rlabel metal2 s 116766 0 116822 800 6 wbs_dat_o[29]
port 369 nsew signal output
rlabel metal2 s 19338 0 19394 800 6 wbs_dat_o[2]
port 370 nsew signal output
rlabel metal2 s 120354 0 120410 800 6 wbs_dat_o[30]
port 371 nsew signal output
rlabel metal2 s 123850 0 123906 800 6 wbs_dat_o[31]
port 372 nsew signal output
rlabel metal2 s 24030 0 24086 800 6 wbs_dat_o[3]
port 373 nsew signal output
rlabel metal2 s 28722 0 28778 800 6 wbs_dat_o[4]
port 374 nsew signal output
rlabel metal2 s 32218 0 32274 800 6 wbs_dat_o[5]
port 375 nsew signal output
rlabel metal2 s 35714 0 35770 800 6 wbs_dat_o[6]
port 376 nsew signal output
rlabel metal2 s 39302 0 39358 800 6 wbs_dat_o[7]
port 377 nsew signal output
rlabel metal2 s 42798 0 42854 800 6 wbs_dat_o[8]
port 378 nsew signal output
rlabel metal2 s 46294 0 46350 800 6 wbs_dat_o[9]
port 379 nsew signal output
rlabel metal2 s 11058 0 11114 800 6 wbs_sel_i[0]
port 380 nsew signal input
rlabel metal2 s 15750 0 15806 800 6 wbs_sel_i[1]
port 381 nsew signal input
rlabel metal2 s 20534 0 20590 800 6 wbs_sel_i[2]
port 382 nsew signal input
rlabel metal2 s 25226 0 25282 800 6 wbs_sel_i[3]
port 383 nsew signal input
rlabel metal2 s 5262 0 5318 800 6 wbs_stb_i
port 384 nsew signal input
rlabel metal2 s 6366 0 6422 800 6 wbs_we_i
port 385 nsew signal input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 165570 167714
string LEFview TRUE
string GDS_FILE /project/openlane/user_proj/runs/user_proj/results/magic/user_proj.gds
string GDS_END 71126858
string GDS_START 110
<< end >>

