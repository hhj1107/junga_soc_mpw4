magic
tech sky130A
magscale 1 2
timestamp 1640496040
<< obsli1 >>
rect 1104 2159 164559 164305
<< obsm1 >>
rect 14 688 164574 164336
<< metal2 >>
rect 478 165957 534 166757
rect 1398 165957 1454 166757
rect 2318 165957 2374 166757
rect 3238 165957 3294 166757
rect 4250 165957 4306 166757
rect 5170 165957 5226 166757
rect 6090 165957 6146 166757
rect 7010 165957 7066 166757
rect 8022 165957 8078 166757
rect 8942 165957 8998 166757
rect 9862 165957 9918 166757
rect 10874 165957 10930 166757
rect 11794 165957 11850 166757
rect 12714 165957 12770 166757
rect 13634 165957 13690 166757
rect 14646 165957 14702 166757
rect 15566 165957 15622 166757
rect 16486 165957 16542 166757
rect 17498 165957 17554 166757
rect 18418 165957 18474 166757
rect 19338 165957 19394 166757
rect 20258 165957 20314 166757
rect 21270 165957 21326 166757
rect 22190 165957 22246 166757
rect 23110 165957 23166 166757
rect 24122 165957 24178 166757
rect 25042 165957 25098 166757
rect 25962 165957 26018 166757
rect 26882 165957 26938 166757
rect 27894 165957 27950 166757
rect 28814 165957 28870 166757
rect 29734 165957 29790 166757
rect 30746 165957 30802 166757
rect 31666 165957 31722 166757
rect 32586 165957 32642 166757
rect 33506 165957 33562 166757
rect 34518 165957 34574 166757
rect 35438 165957 35494 166757
rect 36358 165957 36414 166757
rect 37278 165957 37334 166757
rect 38290 165957 38346 166757
rect 39210 165957 39266 166757
rect 40130 165957 40186 166757
rect 41142 165957 41198 166757
rect 42062 165957 42118 166757
rect 42982 165957 43038 166757
rect 43902 165957 43958 166757
rect 44914 165957 44970 166757
rect 45834 165957 45890 166757
rect 46754 165957 46810 166757
rect 47766 165957 47822 166757
rect 48686 165957 48742 166757
rect 49606 165957 49662 166757
rect 50526 165957 50582 166757
rect 51538 165957 51594 166757
rect 52458 165957 52514 166757
rect 53378 165957 53434 166757
rect 54390 165957 54446 166757
rect 55310 165957 55366 166757
rect 56230 165957 56286 166757
rect 57150 165957 57206 166757
rect 58162 165957 58218 166757
rect 59082 165957 59138 166757
rect 60002 165957 60058 166757
rect 61014 165957 61070 166757
rect 61934 165957 61990 166757
rect 62854 165957 62910 166757
rect 63774 165957 63830 166757
rect 64786 165957 64842 166757
rect 65706 165957 65762 166757
rect 66626 165957 66682 166757
rect 67546 165957 67602 166757
rect 68558 165957 68614 166757
rect 69478 165957 69534 166757
rect 70398 165957 70454 166757
rect 71410 165957 71466 166757
rect 72330 165957 72386 166757
rect 73250 165957 73306 166757
rect 74170 165957 74226 166757
rect 75182 165957 75238 166757
rect 76102 165957 76158 166757
rect 77022 165957 77078 166757
rect 78034 165957 78090 166757
rect 78954 165957 79010 166757
rect 79874 165957 79930 166757
rect 80794 165957 80850 166757
rect 81806 165957 81862 166757
rect 82726 165957 82782 166757
rect 83646 165957 83702 166757
rect 84658 165957 84714 166757
rect 85578 165957 85634 166757
rect 86498 165957 86554 166757
rect 87418 165957 87474 166757
rect 88430 165957 88486 166757
rect 89350 165957 89406 166757
rect 90270 165957 90326 166757
rect 91282 165957 91338 166757
rect 92202 165957 92258 166757
rect 93122 165957 93178 166757
rect 94042 165957 94098 166757
rect 95054 165957 95110 166757
rect 95974 165957 96030 166757
rect 96894 165957 96950 166757
rect 97906 165957 97962 166757
rect 98826 165957 98882 166757
rect 99746 165957 99802 166757
rect 100666 165957 100722 166757
rect 101678 165957 101734 166757
rect 102598 165957 102654 166757
rect 103518 165957 103574 166757
rect 104438 165957 104494 166757
rect 105450 165957 105506 166757
rect 106370 165957 106426 166757
rect 107290 165957 107346 166757
rect 108302 165957 108358 166757
rect 109222 165957 109278 166757
rect 110142 165957 110198 166757
rect 111062 165957 111118 166757
rect 112074 165957 112130 166757
rect 112994 165957 113050 166757
rect 113914 165957 113970 166757
rect 114926 165957 114982 166757
rect 115846 165957 115902 166757
rect 116766 165957 116822 166757
rect 117686 165957 117742 166757
rect 118698 165957 118754 166757
rect 119618 165957 119674 166757
rect 120538 165957 120594 166757
rect 121550 165957 121606 166757
rect 122470 165957 122526 166757
rect 123390 165957 123446 166757
rect 124310 165957 124366 166757
rect 125322 165957 125378 166757
rect 126242 165957 126298 166757
rect 127162 165957 127218 166757
rect 128174 165957 128230 166757
rect 129094 165957 129150 166757
rect 130014 165957 130070 166757
rect 130934 165957 130990 166757
rect 131946 165957 132002 166757
rect 132866 165957 132922 166757
rect 133786 165957 133842 166757
rect 134706 165957 134762 166757
rect 135718 165957 135774 166757
rect 136638 165957 136694 166757
rect 137558 165957 137614 166757
rect 138570 165957 138626 166757
rect 139490 165957 139546 166757
rect 140410 165957 140466 166757
rect 141330 165957 141386 166757
rect 142342 165957 142398 166757
rect 143262 165957 143318 166757
rect 144182 165957 144238 166757
rect 145194 165957 145250 166757
rect 146114 165957 146170 166757
rect 147034 165957 147090 166757
rect 147954 165957 148010 166757
rect 148966 165957 149022 166757
rect 149886 165957 149942 166757
rect 150806 165957 150862 166757
rect 151818 165957 151874 166757
rect 152738 165957 152794 166757
rect 153658 165957 153714 166757
rect 154578 165957 154634 166757
rect 155590 165957 155646 166757
rect 156510 165957 156566 166757
rect 157430 165957 157486 166757
rect 158442 165957 158498 166757
rect 159362 165957 159418 166757
rect 160282 165957 160338 166757
rect 161202 165957 161258 166757
rect 162214 165957 162270 166757
rect 163134 165957 163190 166757
rect 164054 165957 164110 166757
rect 478 0 534 800
rect 1398 0 1454 800
rect 2318 0 2374 800
rect 3330 0 3386 800
rect 4250 0 4306 800
rect 5262 0 5318 800
rect 6182 0 6238 800
rect 7102 0 7158 800
rect 8114 0 8170 800
rect 9034 0 9090 800
rect 10046 0 10102 800
rect 10966 0 11022 800
rect 11886 0 11942 800
rect 12898 0 12954 800
rect 13818 0 13874 800
rect 14830 0 14886 800
rect 15750 0 15806 800
rect 16670 0 16726 800
rect 17682 0 17738 800
rect 18602 0 18658 800
rect 19614 0 19670 800
rect 20534 0 20590 800
rect 21454 0 21510 800
rect 22466 0 22522 800
rect 23386 0 23442 800
rect 24398 0 24454 800
rect 25318 0 25374 800
rect 26238 0 26294 800
rect 27250 0 27306 800
rect 28170 0 28226 800
rect 29182 0 29238 800
rect 30102 0 30158 800
rect 31022 0 31078 800
rect 32034 0 32090 800
rect 32954 0 33010 800
rect 33966 0 34022 800
rect 34886 0 34942 800
rect 35806 0 35862 800
rect 36818 0 36874 800
rect 37738 0 37794 800
rect 38750 0 38806 800
rect 39670 0 39726 800
rect 40590 0 40646 800
rect 41602 0 41658 800
rect 42522 0 42578 800
rect 43534 0 43590 800
rect 44454 0 44510 800
rect 45374 0 45430 800
rect 46386 0 46442 800
rect 47306 0 47362 800
rect 48318 0 48374 800
rect 49238 0 49294 800
rect 50158 0 50214 800
rect 51170 0 51226 800
rect 52090 0 52146 800
rect 53102 0 53158 800
rect 54022 0 54078 800
rect 54942 0 54998 800
rect 55954 0 56010 800
rect 56874 0 56930 800
rect 57886 0 57942 800
rect 58806 0 58862 800
rect 59726 0 59782 800
rect 60738 0 60794 800
rect 61658 0 61714 800
rect 62670 0 62726 800
rect 63590 0 63646 800
rect 64510 0 64566 800
rect 65522 0 65578 800
rect 66442 0 66498 800
rect 67454 0 67510 800
rect 68374 0 68430 800
rect 69294 0 69350 800
rect 70306 0 70362 800
rect 71226 0 71282 800
rect 72238 0 72294 800
rect 73158 0 73214 800
rect 74078 0 74134 800
rect 75090 0 75146 800
rect 76010 0 76066 800
rect 77022 0 77078 800
rect 77942 0 77998 800
rect 78862 0 78918 800
rect 79874 0 79930 800
rect 80794 0 80850 800
rect 81806 0 81862 800
rect 82726 0 82782 800
rect 83646 0 83702 800
rect 84658 0 84714 800
rect 85578 0 85634 800
rect 86590 0 86646 800
rect 87510 0 87566 800
rect 88430 0 88486 800
rect 89442 0 89498 800
rect 90362 0 90418 800
rect 91374 0 91430 800
rect 92294 0 92350 800
rect 93214 0 93270 800
rect 94226 0 94282 800
rect 95146 0 95202 800
rect 96158 0 96214 800
rect 97078 0 97134 800
rect 97998 0 98054 800
rect 99010 0 99066 800
rect 99930 0 99986 800
rect 100942 0 100998 800
rect 101862 0 101918 800
rect 102782 0 102838 800
rect 103794 0 103850 800
rect 104714 0 104770 800
rect 105726 0 105782 800
rect 106646 0 106702 800
rect 107566 0 107622 800
rect 108578 0 108634 800
rect 109498 0 109554 800
rect 110510 0 110566 800
rect 111430 0 111486 800
rect 112350 0 112406 800
rect 113362 0 113418 800
rect 114282 0 114338 800
rect 115294 0 115350 800
rect 116214 0 116270 800
rect 117134 0 117190 800
rect 118146 0 118202 800
rect 119066 0 119122 800
rect 120078 0 120134 800
rect 120998 0 121054 800
rect 121918 0 121974 800
rect 122930 0 122986 800
rect 123850 0 123906 800
rect 124862 0 124918 800
rect 125782 0 125838 800
rect 126702 0 126758 800
rect 127714 0 127770 800
rect 128634 0 128690 800
rect 129646 0 129702 800
rect 130566 0 130622 800
rect 131486 0 131542 800
rect 132498 0 132554 800
rect 133418 0 133474 800
rect 134430 0 134486 800
rect 135350 0 135406 800
rect 136270 0 136326 800
rect 137282 0 137338 800
rect 138202 0 138258 800
rect 139214 0 139270 800
rect 140134 0 140190 800
rect 141054 0 141110 800
rect 142066 0 142122 800
rect 142986 0 143042 800
rect 143998 0 144054 800
rect 144918 0 144974 800
rect 145838 0 145894 800
rect 146850 0 146906 800
rect 147770 0 147826 800
rect 148782 0 148838 800
rect 149702 0 149758 800
rect 150622 0 150678 800
rect 151634 0 151690 800
rect 152554 0 152610 800
rect 153566 0 153622 800
rect 154486 0 154542 800
rect 155406 0 155462 800
rect 156418 0 156474 800
rect 157338 0 157394 800
rect 158350 0 158406 800
rect 159270 0 159326 800
rect 160190 0 160246 800
rect 161202 0 161258 800
rect 162122 0 162178 800
rect 163134 0 163190 800
rect 164054 0 164110 800
<< obsm2 >>
rect 20 165901 422 166002
rect 590 165901 1342 166002
rect 1510 165901 2262 166002
rect 2430 165901 3182 166002
rect 3350 165901 4194 166002
rect 4362 165901 5114 166002
rect 5282 165901 6034 166002
rect 6202 165901 6954 166002
rect 7122 165901 7966 166002
rect 8134 165901 8886 166002
rect 9054 165901 9806 166002
rect 9974 165901 10818 166002
rect 10986 165901 11738 166002
rect 11906 165901 12658 166002
rect 12826 165901 13578 166002
rect 13746 165901 14590 166002
rect 14758 165901 15510 166002
rect 15678 165901 16430 166002
rect 16598 165901 17442 166002
rect 17610 165901 18362 166002
rect 18530 165901 19282 166002
rect 19450 165901 20202 166002
rect 20370 165901 21214 166002
rect 21382 165901 22134 166002
rect 22302 165901 23054 166002
rect 23222 165901 24066 166002
rect 24234 165901 24986 166002
rect 25154 165901 25906 166002
rect 26074 165901 26826 166002
rect 26994 165901 27838 166002
rect 28006 165901 28758 166002
rect 28926 165901 29678 166002
rect 29846 165901 30690 166002
rect 30858 165901 31610 166002
rect 31778 165901 32530 166002
rect 32698 165901 33450 166002
rect 33618 165901 34462 166002
rect 34630 165901 35382 166002
rect 35550 165901 36302 166002
rect 36470 165901 37222 166002
rect 37390 165901 38234 166002
rect 38402 165901 39154 166002
rect 39322 165901 40074 166002
rect 40242 165901 41086 166002
rect 41254 165901 42006 166002
rect 42174 165901 42926 166002
rect 43094 165901 43846 166002
rect 44014 165901 44858 166002
rect 45026 165901 45778 166002
rect 45946 165901 46698 166002
rect 46866 165901 47710 166002
rect 47878 165901 48630 166002
rect 48798 165901 49550 166002
rect 49718 165901 50470 166002
rect 50638 165901 51482 166002
rect 51650 165901 52402 166002
rect 52570 165901 53322 166002
rect 53490 165901 54334 166002
rect 54502 165901 55254 166002
rect 55422 165901 56174 166002
rect 56342 165901 57094 166002
rect 57262 165901 58106 166002
rect 58274 165901 59026 166002
rect 59194 165901 59946 166002
rect 60114 165901 60958 166002
rect 61126 165901 61878 166002
rect 62046 165901 62798 166002
rect 62966 165901 63718 166002
rect 63886 165901 64730 166002
rect 64898 165901 65650 166002
rect 65818 165901 66570 166002
rect 66738 165901 67490 166002
rect 67658 165901 68502 166002
rect 68670 165901 69422 166002
rect 69590 165901 70342 166002
rect 70510 165901 71354 166002
rect 71522 165901 72274 166002
rect 72442 165901 73194 166002
rect 73362 165901 74114 166002
rect 74282 165901 75126 166002
rect 75294 165901 76046 166002
rect 76214 165901 76966 166002
rect 77134 165901 77978 166002
rect 78146 165901 78898 166002
rect 79066 165901 79818 166002
rect 79986 165901 80738 166002
rect 80906 165901 81750 166002
rect 81918 165901 82670 166002
rect 82838 165901 83590 166002
rect 83758 165901 84602 166002
rect 84770 165901 85522 166002
rect 85690 165901 86442 166002
rect 86610 165901 87362 166002
rect 87530 165901 88374 166002
rect 88542 165901 89294 166002
rect 89462 165901 90214 166002
rect 90382 165901 91226 166002
rect 91394 165901 92146 166002
rect 92314 165901 93066 166002
rect 93234 165901 93986 166002
rect 94154 165901 94998 166002
rect 95166 165901 95918 166002
rect 96086 165901 96838 166002
rect 97006 165901 97850 166002
rect 98018 165901 98770 166002
rect 98938 165901 99690 166002
rect 99858 165901 100610 166002
rect 100778 165901 101622 166002
rect 101790 165901 102542 166002
rect 102710 165901 103462 166002
rect 103630 165901 104382 166002
rect 104550 165901 105394 166002
rect 105562 165901 106314 166002
rect 106482 165901 107234 166002
rect 107402 165901 108246 166002
rect 108414 165901 109166 166002
rect 109334 165901 110086 166002
rect 110254 165901 111006 166002
rect 111174 165901 112018 166002
rect 112186 165901 112938 166002
rect 113106 165901 113858 166002
rect 114026 165901 114870 166002
rect 115038 165901 115790 166002
rect 115958 165901 116710 166002
rect 116878 165901 117630 166002
rect 117798 165901 118642 166002
rect 118810 165901 119562 166002
rect 119730 165901 120482 166002
rect 120650 165901 121494 166002
rect 121662 165901 122414 166002
rect 122582 165901 123334 166002
rect 123502 165901 124254 166002
rect 124422 165901 125266 166002
rect 125434 165901 126186 166002
rect 126354 165901 127106 166002
rect 127274 165901 128118 166002
rect 128286 165901 129038 166002
rect 129206 165901 129958 166002
rect 130126 165901 130878 166002
rect 131046 165901 131890 166002
rect 132058 165901 132810 166002
rect 132978 165901 133730 166002
rect 133898 165901 134650 166002
rect 134818 165901 135662 166002
rect 135830 165901 136582 166002
rect 136750 165901 137502 166002
rect 137670 165901 138514 166002
rect 138682 165901 139434 166002
rect 139602 165901 140354 166002
rect 140522 165901 141274 166002
rect 141442 165901 142286 166002
rect 142454 165901 143206 166002
rect 143374 165901 144126 166002
rect 144294 165901 145138 166002
rect 145306 165901 146058 166002
rect 146226 165901 146978 166002
rect 147146 165901 147898 166002
rect 148066 165901 148910 166002
rect 149078 165901 149830 166002
rect 149998 165901 150750 166002
rect 150918 165901 151762 166002
rect 151930 165901 152682 166002
rect 152850 165901 153602 166002
rect 153770 165901 154522 166002
rect 154690 165901 155534 166002
rect 155702 165901 156454 166002
rect 156622 165901 157374 166002
rect 157542 165901 158386 166002
rect 158554 165901 159306 166002
rect 159474 165901 160226 166002
rect 160394 165901 161146 166002
rect 161314 165901 162158 166002
rect 162326 165901 163078 166002
rect 163246 165901 163998 166002
rect 164166 165901 164570 166002
rect 20 856 164570 165901
rect 20 575 422 856
rect 590 575 1342 856
rect 1510 575 2262 856
rect 2430 575 3274 856
rect 3442 575 4194 856
rect 4362 575 5206 856
rect 5374 575 6126 856
rect 6294 575 7046 856
rect 7214 575 8058 856
rect 8226 575 8978 856
rect 9146 575 9990 856
rect 10158 575 10910 856
rect 11078 575 11830 856
rect 11998 575 12842 856
rect 13010 575 13762 856
rect 13930 575 14774 856
rect 14942 575 15694 856
rect 15862 575 16614 856
rect 16782 575 17626 856
rect 17794 575 18546 856
rect 18714 575 19558 856
rect 19726 575 20478 856
rect 20646 575 21398 856
rect 21566 575 22410 856
rect 22578 575 23330 856
rect 23498 575 24342 856
rect 24510 575 25262 856
rect 25430 575 26182 856
rect 26350 575 27194 856
rect 27362 575 28114 856
rect 28282 575 29126 856
rect 29294 575 30046 856
rect 30214 575 30966 856
rect 31134 575 31978 856
rect 32146 575 32898 856
rect 33066 575 33910 856
rect 34078 575 34830 856
rect 34998 575 35750 856
rect 35918 575 36762 856
rect 36930 575 37682 856
rect 37850 575 38694 856
rect 38862 575 39614 856
rect 39782 575 40534 856
rect 40702 575 41546 856
rect 41714 575 42466 856
rect 42634 575 43478 856
rect 43646 575 44398 856
rect 44566 575 45318 856
rect 45486 575 46330 856
rect 46498 575 47250 856
rect 47418 575 48262 856
rect 48430 575 49182 856
rect 49350 575 50102 856
rect 50270 575 51114 856
rect 51282 575 52034 856
rect 52202 575 53046 856
rect 53214 575 53966 856
rect 54134 575 54886 856
rect 55054 575 55898 856
rect 56066 575 56818 856
rect 56986 575 57830 856
rect 57998 575 58750 856
rect 58918 575 59670 856
rect 59838 575 60682 856
rect 60850 575 61602 856
rect 61770 575 62614 856
rect 62782 575 63534 856
rect 63702 575 64454 856
rect 64622 575 65466 856
rect 65634 575 66386 856
rect 66554 575 67398 856
rect 67566 575 68318 856
rect 68486 575 69238 856
rect 69406 575 70250 856
rect 70418 575 71170 856
rect 71338 575 72182 856
rect 72350 575 73102 856
rect 73270 575 74022 856
rect 74190 575 75034 856
rect 75202 575 75954 856
rect 76122 575 76966 856
rect 77134 575 77886 856
rect 78054 575 78806 856
rect 78974 575 79818 856
rect 79986 575 80738 856
rect 80906 575 81750 856
rect 81918 575 82670 856
rect 82838 575 83590 856
rect 83758 575 84602 856
rect 84770 575 85522 856
rect 85690 575 86534 856
rect 86702 575 87454 856
rect 87622 575 88374 856
rect 88542 575 89386 856
rect 89554 575 90306 856
rect 90474 575 91318 856
rect 91486 575 92238 856
rect 92406 575 93158 856
rect 93326 575 94170 856
rect 94338 575 95090 856
rect 95258 575 96102 856
rect 96270 575 97022 856
rect 97190 575 97942 856
rect 98110 575 98954 856
rect 99122 575 99874 856
rect 100042 575 100886 856
rect 101054 575 101806 856
rect 101974 575 102726 856
rect 102894 575 103738 856
rect 103906 575 104658 856
rect 104826 575 105670 856
rect 105838 575 106590 856
rect 106758 575 107510 856
rect 107678 575 108522 856
rect 108690 575 109442 856
rect 109610 575 110454 856
rect 110622 575 111374 856
rect 111542 575 112294 856
rect 112462 575 113306 856
rect 113474 575 114226 856
rect 114394 575 115238 856
rect 115406 575 116158 856
rect 116326 575 117078 856
rect 117246 575 118090 856
rect 118258 575 119010 856
rect 119178 575 120022 856
rect 120190 575 120942 856
rect 121110 575 121862 856
rect 122030 575 122874 856
rect 123042 575 123794 856
rect 123962 575 124806 856
rect 124974 575 125726 856
rect 125894 575 126646 856
rect 126814 575 127658 856
rect 127826 575 128578 856
rect 128746 575 129590 856
rect 129758 575 130510 856
rect 130678 575 131430 856
rect 131598 575 132442 856
rect 132610 575 133362 856
rect 133530 575 134374 856
rect 134542 575 135294 856
rect 135462 575 136214 856
rect 136382 575 137226 856
rect 137394 575 138146 856
rect 138314 575 139158 856
rect 139326 575 140078 856
rect 140246 575 140998 856
rect 141166 575 142010 856
rect 142178 575 142930 856
rect 143098 575 143942 856
rect 144110 575 144862 856
rect 145030 575 145782 856
rect 145950 575 146794 856
rect 146962 575 147714 856
rect 147882 575 148726 856
rect 148894 575 149646 856
rect 149814 575 150566 856
rect 150734 575 151578 856
rect 151746 575 152498 856
rect 152666 575 153510 856
rect 153678 575 154430 856
rect 154598 575 155350 856
rect 155518 575 156362 856
rect 156530 575 157282 856
rect 157450 575 158294 856
rect 158462 575 159214 856
rect 159382 575 160134 856
rect 160302 575 161146 856
rect 161314 575 162066 856
rect 162234 575 163078 856
rect 163246 575 163998 856
rect 164166 575 164570 856
<< metal3 >>
rect 0 165112 800 165232
rect 163813 165248 164613 165368
rect 163813 162664 164613 162784
rect 0 162120 800 162240
rect 163813 160080 164613 160200
rect 0 159128 800 159248
rect 163813 157496 164613 157616
rect 0 156000 800 156120
rect 163813 154912 164613 155032
rect 0 153008 800 153128
rect 163813 152328 164613 152448
rect 0 150016 800 150136
rect 163813 149608 164613 149728
rect 0 146888 800 147008
rect 163813 147024 164613 147144
rect 163813 144440 164613 144560
rect 0 143896 800 144016
rect 163813 141856 164613 141976
rect 0 140904 800 141024
rect 163813 139272 164613 139392
rect 0 137912 800 138032
rect 163813 136688 164613 136808
rect 0 134784 800 134904
rect 163813 133968 164613 134088
rect 0 131792 800 131912
rect 163813 131384 164613 131504
rect 0 128800 800 128920
rect 163813 128800 164613 128920
rect 163813 126216 164613 126336
rect 0 125672 800 125792
rect 163813 123632 164613 123752
rect 0 122680 800 122800
rect 163813 121048 164613 121168
rect 0 119688 800 119808
rect 163813 118464 164613 118584
rect 0 116696 800 116816
rect 163813 115744 164613 115864
rect 0 113568 800 113688
rect 163813 113160 164613 113280
rect 0 110576 800 110696
rect 163813 110576 164613 110696
rect 163813 107992 164613 108112
rect 0 107584 800 107704
rect 163813 105408 164613 105528
rect 0 104456 800 104576
rect 163813 102824 164613 102944
rect 0 101464 800 101584
rect 163813 100104 164613 100224
rect 0 98472 800 98592
rect 163813 97520 164613 97640
rect 0 95480 800 95600
rect 163813 94936 164613 95056
rect 0 92352 800 92472
rect 163813 92352 164613 92472
rect 163813 89768 164613 89888
rect 0 89360 800 89480
rect 163813 87184 164613 87304
rect 0 86368 800 86488
rect 163813 84600 164613 84720
rect 0 83240 800 83360
rect 163813 81880 164613 82000
rect 0 80248 800 80368
rect 163813 79296 164613 79416
rect 0 77256 800 77376
rect 163813 76712 164613 76832
rect 0 74128 800 74248
rect 163813 74128 164613 74248
rect 163813 71544 164613 71664
rect 0 71136 800 71256
rect 163813 68960 164613 69080
rect 0 68144 800 68264
rect 163813 66240 164613 66360
rect 0 65152 800 65272
rect 163813 63656 164613 63776
rect 0 62024 800 62144
rect 163813 61072 164613 61192
rect 0 59032 800 59152
rect 163813 58488 164613 58608
rect 0 56040 800 56160
rect 163813 55904 164613 56024
rect 163813 53320 164613 53440
rect 0 52912 800 53032
rect 163813 50600 164613 50720
rect 0 49920 800 50040
rect 163813 48016 164613 48136
rect 0 46928 800 47048
rect 163813 45432 164613 45552
rect 0 43936 800 44056
rect 163813 42848 164613 42968
rect 0 40808 800 40928
rect 163813 40264 164613 40384
rect 0 37816 800 37936
rect 163813 37680 164613 37800
rect 163813 35096 164613 35216
rect 0 34824 800 34944
rect 163813 32376 164613 32496
rect 0 31696 800 31816
rect 163813 29792 164613 29912
rect 0 28704 800 28824
rect 163813 27208 164613 27328
rect 0 25712 800 25832
rect 163813 24624 164613 24744
rect 0 22720 800 22840
rect 163813 22040 164613 22160
rect 0 19592 800 19712
rect 163813 19456 164613 19576
rect 0 16600 800 16720
rect 163813 16736 164613 16856
rect 163813 14152 164613 14272
rect 0 13608 800 13728
rect 163813 11568 164613 11688
rect 0 10480 800 10600
rect 163813 8984 164613 9104
rect 0 7488 800 7608
rect 163813 6400 164613 6520
rect 0 4496 800 4616
rect 163813 3816 164613 3936
rect 0 1504 800 1624
rect 163813 1232 164613 1352
<< obsm3 >>
rect 800 165312 163733 165341
rect 880 165168 163733 165312
rect 880 165032 164580 165168
rect 800 162864 164580 165032
rect 800 162584 163733 162864
rect 800 162320 164580 162584
rect 880 162040 164580 162320
rect 800 160280 164580 162040
rect 800 160000 163733 160280
rect 800 159328 164580 160000
rect 880 159048 164580 159328
rect 800 157696 164580 159048
rect 800 157416 163733 157696
rect 800 156200 164580 157416
rect 880 155920 164580 156200
rect 800 155112 164580 155920
rect 800 154832 163733 155112
rect 800 153208 164580 154832
rect 880 152928 164580 153208
rect 800 152528 164580 152928
rect 800 152248 163733 152528
rect 800 150216 164580 152248
rect 880 149936 164580 150216
rect 800 149808 164580 149936
rect 800 149528 163733 149808
rect 800 147224 164580 149528
rect 800 147088 163733 147224
rect 880 146944 163733 147088
rect 880 146808 164580 146944
rect 800 144640 164580 146808
rect 800 144360 163733 144640
rect 800 144096 164580 144360
rect 880 143816 164580 144096
rect 800 142056 164580 143816
rect 800 141776 163733 142056
rect 800 141104 164580 141776
rect 880 140824 164580 141104
rect 800 139472 164580 140824
rect 800 139192 163733 139472
rect 800 138112 164580 139192
rect 880 137832 164580 138112
rect 800 136888 164580 137832
rect 800 136608 163733 136888
rect 800 134984 164580 136608
rect 880 134704 164580 134984
rect 800 134168 164580 134704
rect 800 133888 163733 134168
rect 800 131992 164580 133888
rect 880 131712 164580 131992
rect 800 131584 164580 131712
rect 800 131304 163733 131584
rect 800 129000 164580 131304
rect 880 128720 163733 129000
rect 800 126416 164580 128720
rect 800 126136 163733 126416
rect 800 125872 164580 126136
rect 880 125592 164580 125872
rect 800 123832 164580 125592
rect 800 123552 163733 123832
rect 800 122880 164580 123552
rect 880 122600 164580 122880
rect 800 121248 164580 122600
rect 800 120968 163733 121248
rect 800 119888 164580 120968
rect 880 119608 164580 119888
rect 800 118664 164580 119608
rect 800 118384 163733 118664
rect 800 116896 164580 118384
rect 880 116616 164580 116896
rect 800 115944 164580 116616
rect 800 115664 163733 115944
rect 800 113768 164580 115664
rect 880 113488 164580 113768
rect 800 113360 164580 113488
rect 800 113080 163733 113360
rect 800 110776 164580 113080
rect 880 110496 163733 110776
rect 800 108192 164580 110496
rect 800 107912 163733 108192
rect 800 107784 164580 107912
rect 880 107504 164580 107784
rect 800 105608 164580 107504
rect 800 105328 163733 105608
rect 800 104656 164580 105328
rect 880 104376 164580 104656
rect 800 103024 164580 104376
rect 800 102744 163733 103024
rect 800 101664 164580 102744
rect 880 101384 164580 101664
rect 800 100304 164580 101384
rect 800 100024 163733 100304
rect 800 98672 164580 100024
rect 880 98392 164580 98672
rect 800 97720 164580 98392
rect 800 97440 163733 97720
rect 800 95680 164580 97440
rect 880 95400 164580 95680
rect 800 95136 164580 95400
rect 800 94856 163733 95136
rect 800 92552 164580 94856
rect 880 92272 163733 92552
rect 800 89968 164580 92272
rect 800 89688 163733 89968
rect 800 89560 164580 89688
rect 880 89280 164580 89560
rect 800 87384 164580 89280
rect 800 87104 163733 87384
rect 800 86568 164580 87104
rect 880 86288 164580 86568
rect 800 84800 164580 86288
rect 800 84520 163733 84800
rect 800 83440 164580 84520
rect 880 83160 164580 83440
rect 800 82080 164580 83160
rect 800 81800 163733 82080
rect 800 80448 164580 81800
rect 880 80168 164580 80448
rect 800 79496 164580 80168
rect 800 79216 163733 79496
rect 800 77456 164580 79216
rect 880 77176 164580 77456
rect 800 76912 164580 77176
rect 800 76632 163733 76912
rect 800 74328 164580 76632
rect 880 74048 163733 74328
rect 800 71744 164580 74048
rect 800 71464 163733 71744
rect 800 71336 164580 71464
rect 880 71056 164580 71336
rect 800 69160 164580 71056
rect 800 68880 163733 69160
rect 800 68344 164580 68880
rect 880 68064 164580 68344
rect 800 66440 164580 68064
rect 800 66160 163733 66440
rect 800 65352 164580 66160
rect 880 65072 164580 65352
rect 800 63856 164580 65072
rect 800 63576 163733 63856
rect 800 62224 164580 63576
rect 880 61944 164580 62224
rect 800 61272 164580 61944
rect 800 60992 163733 61272
rect 800 59232 164580 60992
rect 880 58952 164580 59232
rect 800 58688 164580 58952
rect 800 58408 163733 58688
rect 800 56240 164580 58408
rect 880 56104 164580 56240
rect 880 55960 163733 56104
rect 800 55824 163733 55960
rect 800 53520 164580 55824
rect 800 53240 163733 53520
rect 800 53112 164580 53240
rect 880 52832 164580 53112
rect 800 50800 164580 52832
rect 800 50520 163733 50800
rect 800 50120 164580 50520
rect 880 49840 164580 50120
rect 800 48216 164580 49840
rect 800 47936 163733 48216
rect 800 47128 164580 47936
rect 880 46848 164580 47128
rect 800 45632 164580 46848
rect 800 45352 163733 45632
rect 800 44136 164580 45352
rect 880 43856 164580 44136
rect 800 43048 164580 43856
rect 800 42768 163733 43048
rect 800 41008 164580 42768
rect 880 40728 164580 41008
rect 800 40464 164580 40728
rect 800 40184 163733 40464
rect 800 38016 164580 40184
rect 880 37880 164580 38016
rect 880 37736 163733 37880
rect 800 37600 163733 37736
rect 800 35296 164580 37600
rect 800 35024 163733 35296
rect 880 35016 163733 35024
rect 880 34744 164580 35016
rect 800 32576 164580 34744
rect 800 32296 163733 32576
rect 800 31896 164580 32296
rect 880 31616 164580 31896
rect 800 29992 164580 31616
rect 800 29712 163733 29992
rect 800 28904 164580 29712
rect 880 28624 164580 28904
rect 800 27408 164580 28624
rect 800 27128 163733 27408
rect 800 25912 164580 27128
rect 880 25632 164580 25912
rect 800 24824 164580 25632
rect 800 24544 163733 24824
rect 800 22920 164580 24544
rect 880 22640 164580 22920
rect 800 22240 164580 22640
rect 800 21960 163733 22240
rect 800 19792 164580 21960
rect 880 19656 164580 19792
rect 880 19512 163733 19656
rect 800 19376 163733 19512
rect 800 16936 164580 19376
rect 800 16800 163733 16936
rect 880 16656 163733 16800
rect 880 16520 164580 16656
rect 800 14352 164580 16520
rect 800 14072 163733 14352
rect 800 13808 164580 14072
rect 880 13528 164580 13808
rect 800 11768 164580 13528
rect 800 11488 163733 11768
rect 800 10680 164580 11488
rect 880 10400 164580 10680
rect 800 9184 164580 10400
rect 800 8904 163733 9184
rect 800 7688 164580 8904
rect 880 7408 164580 7688
rect 800 6600 164580 7408
rect 800 6320 163733 6600
rect 800 4696 164580 6320
rect 880 4416 164580 4696
rect 800 4016 164580 4416
rect 800 3736 163733 4016
rect 800 1704 164580 3736
rect 880 1432 164580 1704
rect 880 1424 163733 1432
rect 800 1152 163733 1424
rect 800 579 164580 1152
<< metal4 >>
rect 4208 2128 4528 164336
rect 19568 2128 19888 164336
rect 34928 2128 35248 164336
rect 50288 2128 50608 164336
rect 65648 2128 65968 164336
rect 81008 2128 81328 164336
rect 96368 2128 96688 164336
rect 111728 2128 112048 164336
rect 127088 2128 127408 164336
rect 142448 2128 142768 164336
rect 157808 2128 158128 164336
<< obsm4 >>
rect 18459 2048 19488 163981
rect 19968 2048 34848 163981
rect 35328 2048 50208 163981
rect 50688 2048 65568 163981
rect 66048 2048 80928 163981
rect 81408 2048 96288 163981
rect 96768 2048 111648 163981
rect 112128 2048 127008 163981
rect 127488 2048 142368 163981
rect 142848 2048 157728 163981
rect 158208 63610 164613 163981
rect 158208 51854 164618 63610
rect 158208 2048 164613 51854
rect 18459 579 164613 2048
<< labels >>
rlabel metal3 s 163813 6400 164613 6520 6 i_dout0[0]
port 1 nsew signal input
rlabel metal3 s 0 89360 800 89480 6 i_dout0[10]
port 2 nsew signal input
rlabel metal3 s 163813 79296 164613 79416 6 i_dout0[11]
port 3 nsew signal input
rlabel metal2 s 137282 0 137338 800 6 i_dout0[12]
port 4 nsew signal input
rlabel metal3 s 0 92352 800 92472 6 i_dout0[13]
port 5 nsew signal input
rlabel metal3 s 0 101464 800 101584 6 i_dout0[14]
port 6 nsew signal input
rlabel metal3 s 0 110576 800 110696 6 i_dout0[15]
port 7 nsew signal input
rlabel metal2 s 140410 165957 140466 166757 6 i_dout0[16]
port 8 nsew signal input
rlabel metal2 s 142066 0 142122 800 6 i_dout0[17]
port 9 nsew signal input
rlabel metal3 s 163813 110576 164613 110696 6 i_dout0[18]
port 10 nsew signal input
rlabel metal3 s 0 122680 800 122800 6 i_dout0[19]
port 11 nsew signal input
rlabel metal2 s 109498 0 109554 800 6 i_dout0[1]
port 12 nsew signal input
rlabel metal3 s 0 128800 800 128920 6 i_dout0[20]
port 13 nsew signal input
rlabel metal2 s 147770 0 147826 800 6 i_dout0[21]
port 14 nsew signal input
rlabel metal3 s 163813 118464 164613 118584 6 i_dout0[22]
port 15 nsew signal input
rlabel metal3 s 163813 121048 164613 121168 6 i_dout0[23]
port 16 nsew signal input
rlabel metal2 s 156510 165957 156566 166757 6 i_dout0[24]
port 17 nsew signal input
rlabel metal2 s 152554 0 152610 800 6 i_dout0[25]
port 18 nsew signal input
rlabel metal3 s 163813 141856 164613 141976 6 i_dout0[26]
port 19 nsew signal input
rlabel metal3 s 163813 149608 164613 149728 6 i_dout0[27]
port 20 nsew signal input
rlabel metal3 s 163813 154912 164613 155032 6 i_dout0[28]
port 21 nsew signal input
rlabel metal3 s 0 150016 800 150136 6 i_dout0[29]
port 22 nsew signal input
rlabel metal2 s 113362 0 113418 800 6 i_dout0[2]
port 23 nsew signal input
rlabel metal2 s 163134 165957 163190 166757 6 i_dout0[30]
port 24 nsew signal input
rlabel metal3 s 0 165112 800 165232 6 i_dout0[31]
port 25 nsew signal input
rlabel metal3 s 0 37816 800 37936 6 i_dout0[3]
port 26 nsew signal input
rlabel metal3 s 163813 37680 164613 37800 6 i_dout0[4]
port 27 nsew signal input
rlabel metal3 s 0 49920 800 50040 6 i_dout0[5]
port 28 nsew signal input
rlabel metal2 s 124862 0 124918 800 6 i_dout0[6]
port 29 nsew signal input
rlabel metal3 s 163813 50600 164613 50720 6 i_dout0[7]
port 30 nsew signal input
rlabel metal2 s 129646 0 129702 800 6 i_dout0[8]
port 31 nsew signal input
rlabel metal2 s 127162 165957 127218 166757 6 i_dout0[9]
port 32 nsew signal input
rlabel metal3 s 163813 8984 164613 9104 6 i_dout0_1[0]
port 33 nsew signal input
rlabel metal2 s 129094 165957 129150 166757 6 i_dout0_1[10]
port 34 nsew signal input
rlabel metal2 s 131946 165957 132002 166757 6 i_dout0_1[11]
port 35 nsew signal input
rlabel metal2 s 133786 165957 133842 166757 6 i_dout0_1[12]
port 36 nsew signal input
rlabel metal2 s 135718 165957 135774 166757 6 i_dout0_1[13]
port 37 nsew signal input
rlabel metal3 s 0 95480 800 95600 6 i_dout0_1[14]
port 38 nsew signal input
rlabel metal3 s 163813 89768 164613 89888 6 i_dout0_1[15]
port 39 nsew signal input
rlabel metal2 s 139490 165957 139546 166757 6 i_dout0_1[16]
port 40 nsew signal input
rlabel metal2 s 141054 0 141110 800 6 i_dout0_1[17]
port 41 nsew signal input
rlabel metal2 s 144182 165957 144238 166757 6 i_dout0_1[18]
port 42 nsew signal input
rlabel metal2 s 146114 165957 146170 166757 6 i_dout0_1[19]
port 43 nsew signal input
rlabel metal3 s 0 22720 800 22840 6 i_dout0_1[1]
port 44 nsew signal input
rlabel metal3 s 0 125672 800 125792 6 i_dout0_1[20]
port 45 nsew signal input
rlabel metal3 s 163813 115744 164613 115864 6 i_dout0_1[21]
port 46 nsew signal input
rlabel metal3 s 0 134784 800 134904 6 i_dout0_1[22]
port 47 nsew signal input
rlabel metal2 s 153658 165957 153714 166757 6 i_dout0_1[23]
port 48 nsew signal input
rlabel metal3 s 163813 126216 164613 126336 6 i_dout0_1[24]
port 49 nsew signal input
rlabel metal3 s 163813 131384 164613 131504 6 i_dout0_1[25]
port 50 nsew signal input
rlabel metal2 s 153566 0 153622 800 6 i_dout0_1[26]
port 51 nsew signal input
rlabel metal2 s 154486 0 154542 800 6 i_dout0_1[27]
port 52 nsew signal input
rlabel metal2 s 161202 165957 161258 166757 6 i_dout0_1[28]
port 53 nsew signal input
rlabel metal2 s 159270 0 159326 800 6 i_dout0_1[29]
port 54 nsew signal input
rlabel metal3 s 163813 16736 164613 16856 6 i_dout0_1[2]
port 55 nsew signal input
rlabel metal2 s 162214 165957 162270 166757 6 i_dout0_1[30]
port 56 nsew signal input
rlabel metal2 s 162122 0 162178 800 6 i_dout0_1[31]
port 57 nsew signal input
rlabel metal3 s 0 34824 800 34944 6 i_dout0_1[3]
port 58 nsew signal input
rlabel metal2 s 117134 0 117190 800 6 i_dout0_1[4]
port 59 nsew signal input
rlabel metal3 s 0 43936 800 44056 6 i_dout0_1[5]
port 60 nsew signal input
rlabel metal2 s 123850 0 123906 800 6 i_dout0_1[6]
port 61 nsew signal input
rlabel metal3 s 163813 48016 164613 48136 6 i_dout0_1[7]
port 62 nsew signal input
rlabel metal3 s 163813 61072 164613 61192 6 i_dout0_1[8]
port 63 nsew signal input
rlabel metal3 s 163813 74128 164613 74248 6 i_dout0_1[9]
port 64 nsew signal input
rlabel metal2 s 104714 0 104770 800 6 i_dout1[0]
port 65 nsew signal input
rlabel metal2 s 130014 165957 130070 166757 6 i_dout1[10]
port 66 nsew signal input
rlabel metal3 s 163813 81880 164613 82000 6 i_dout1[11]
port 67 nsew signal input
rlabel metal2 s 138202 0 138258 800 6 i_dout1[12]
port 68 nsew signal input
rlabel metal2 s 137558 165957 137614 166757 6 i_dout1[13]
port 69 nsew signal input
rlabel metal3 s 0 104456 800 104576 6 i_dout1[14]
port 70 nsew signal input
rlabel metal3 s 163813 94936 164613 95056 6 i_dout1[15]
port 71 nsew signal input
rlabel metal2 s 141330 165957 141386 166757 6 i_dout1[16]
port 72 nsew signal input
rlabel metal3 s 163813 107992 164613 108112 6 i_dout1[17]
port 73 nsew signal input
rlabel metal3 s 0 116696 800 116816 6 i_dout1[18]
port 74 nsew signal input
rlabel metal2 s 147954 165957 148010 166757 6 i_dout1[19]
port 75 nsew signal input
rlabel metal2 s 110142 165957 110198 166757 6 i_dout1[1]
port 76 nsew signal input
rlabel metal2 s 144918 0 144974 800 6 i_dout1[20]
port 77 nsew signal input
rlabel metal2 s 149886 165957 149942 166757 6 i_dout1[21]
port 78 nsew signal input
rlabel metal2 s 149702 0 149758 800 6 i_dout1[22]
port 79 nsew signal input
rlabel metal2 s 155590 165957 155646 166757 6 i_dout1[23]
port 80 nsew signal input
rlabel metal3 s 163813 128800 164613 128920 6 i_dout1[24]
port 81 nsew signal input
rlabel metal3 s 163813 136688 164613 136808 6 i_dout1[25]
port 82 nsew signal input
rlabel metal3 s 0 140904 800 141024 6 i_dout1[26]
port 83 nsew signal input
rlabel metal3 s 0 143896 800 144016 6 i_dout1[27]
port 84 nsew signal input
rlabel metal3 s 163813 157496 164613 157616 6 i_dout1[28]
port 85 nsew signal input
rlabel metal3 s 0 153008 800 153128 6 i_dout1[29]
port 86 nsew signal input
rlabel metal2 s 114282 0 114338 800 6 i_dout1[2]
port 87 nsew signal input
rlabel metal3 s 0 159128 800 159248 6 i_dout1[30]
port 88 nsew signal input
rlabel metal2 s 164054 165957 164110 166757 6 i_dout1[31]
port 89 nsew signal input
rlabel metal2 s 117686 165957 117742 166757 6 i_dout1[3]
port 90 nsew signal input
rlabel metal2 s 121550 165957 121606 166757 6 i_dout1[4]
port 91 nsew signal input
rlabel metal3 s 163813 45432 164613 45552 6 i_dout1[5]
port 92 nsew signal input
rlabel metal2 s 125782 0 125838 800 6 i_dout1[6]
port 93 nsew signal input
rlabel metal2 s 127714 0 127770 800 6 i_dout1[7]
port 94 nsew signal input
rlabel metal2 s 126242 165957 126298 166757 6 i_dout1[8]
port 95 nsew signal input
rlabel metal2 s 131486 0 131542 800 6 i_dout1[9]
port 96 nsew signal input
rlabel metal2 s 108302 165957 108358 166757 6 i_dout1_1[0]
port 97 nsew signal input
rlabel metal2 s 132498 0 132554 800 6 i_dout1_1[10]
port 98 nsew signal input
rlabel metal2 s 134430 0 134486 800 6 i_dout1_1[11]
port 99 nsew signal input
rlabel metal2 s 136270 0 136326 800 6 i_dout1_1[12]
port 100 nsew signal input
rlabel metal2 s 136638 165957 136694 166757 6 i_dout1_1[13]
port 101 nsew signal input
rlabel metal3 s 0 98472 800 98592 6 i_dout1_1[14]
port 102 nsew signal input
rlabel metal3 s 163813 92352 164613 92472 6 i_dout1_1[15]
port 103 nsew signal input
rlabel metal3 s 163813 100104 164613 100224 6 i_dout1_1[16]
port 104 nsew signal input
rlabel metal3 s 163813 105408 164613 105528 6 i_dout1_1[17]
port 105 nsew signal input
rlabel metal3 s 0 113568 800 113688 6 i_dout1_1[18]
port 106 nsew signal input
rlabel metal2 s 147034 165957 147090 166757 6 i_dout1_1[19]
port 107 nsew signal input
rlabel metal3 s 0 25712 800 25832 6 i_dout1_1[1]
port 108 nsew signal input
rlabel metal2 s 143998 0 144054 800 6 i_dout1_1[20]
port 109 nsew signal input
rlabel metal3 s 0 131792 800 131912 6 i_dout1_1[21]
port 110 nsew signal input
rlabel metal2 s 151818 165957 151874 166757 6 i_dout1_1[22]
port 111 nsew signal input
rlabel metal2 s 154578 165957 154634 166757 6 i_dout1_1[23]
port 112 nsew signal input
rlabel metal3 s 0 137912 800 138032 6 i_dout1_1[24]
port 113 nsew signal input
rlabel metal3 s 163813 133968 164613 134088 6 i_dout1_1[25]
port 114 nsew signal input
rlabel metal2 s 160282 165957 160338 166757 6 i_dout1_1[26]
port 115 nsew signal input
rlabel metal2 s 155406 0 155462 800 6 i_dout1_1[27]
port 116 nsew signal input
rlabel metal3 s 0 146888 800 147008 6 i_dout1_1[28]
port 117 nsew signal input
rlabel metal2 s 160190 0 160246 800 6 i_dout1_1[29]
port 118 nsew signal input
rlabel metal3 s 163813 19456 164613 19576 6 i_dout1_1[2]
port 119 nsew signal input
rlabel metal3 s 163813 160080 164613 160200 6 i_dout1_1[30]
port 120 nsew signal input
rlabel metal2 s 163134 0 163190 800 6 i_dout1_1[31]
port 121 nsew signal input
rlabel metal2 s 115294 0 115350 800 6 i_dout1_1[3]
port 122 nsew signal input
rlabel metal3 s 163813 35096 164613 35216 6 i_dout1_1[4]
port 123 nsew signal input
rlabel metal3 s 0 46928 800 47048 6 i_dout1_1[5]
port 124 nsew signal input
rlabel metal3 s 0 52912 800 53032 6 i_dout1_1[6]
port 125 nsew signal input
rlabel metal3 s 0 71136 800 71256 6 i_dout1_1[7]
port 126 nsew signal input
rlabel metal3 s 163813 63656 164613 63776 6 i_dout1_1[8]
port 127 nsew signal input
rlabel metal3 s 163813 76712 164613 76832 6 i_dout1_1[9]
port 128 nsew signal input
rlabel metal2 s 478 165957 534 166757 6 io_in[0]
port 129 nsew signal input
rlabel metal2 s 28814 165957 28870 166757 6 io_in[10]
port 130 nsew signal input
rlabel metal2 s 31666 165957 31722 166757 6 io_in[11]
port 131 nsew signal input
rlabel metal2 s 34518 165957 34574 166757 6 io_in[12]
port 132 nsew signal input
rlabel metal2 s 37278 165957 37334 166757 6 io_in[13]
port 133 nsew signal input
rlabel metal2 s 40130 165957 40186 166757 6 io_in[14]
port 134 nsew signal input
rlabel metal2 s 42982 165957 43038 166757 6 io_in[15]
port 135 nsew signal input
rlabel metal2 s 45834 165957 45890 166757 6 io_in[16]
port 136 nsew signal input
rlabel metal2 s 48686 165957 48742 166757 6 io_in[17]
port 137 nsew signal input
rlabel metal2 s 51538 165957 51594 166757 6 io_in[18]
port 138 nsew signal input
rlabel metal2 s 54390 165957 54446 166757 6 io_in[19]
port 139 nsew signal input
rlabel metal2 s 3238 165957 3294 166757 6 io_in[1]
port 140 nsew signal input
rlabel metal2 s 57150 165957 57206 166757 6 io_in[20]
port 141 nsew signal input
rlabel metal2 s 60002 165957 60058 166757 6 io_in[21]
port 142 nsew signal input
rlabel metal2 s 62854 165957 62910 166757 6 io_in[22]
port 143 nsew signal input
rlabel metal2 s 65706 165957 65762 166757 6 io_in[23]
port 144 nsew signal input
rlabel metal2 s 68558 165957 68614 166757 6 io_in[24]
port 145 nsew signal input
rlabel metal2 s 71410 165957 71466 166757 6 io_in[25]
port 146 nsew signal input
rlabel metal2 s 74170 165957 74226 166757 6 io_in[26]
port 147 nsew signal input
rlabel metal2 s 77022 165957 77078 166757 6 io_in[27]
port 148 nsew signal input
rlabel metal2 s 79874 165957 79930 166757 6 io_in[28]
port 149 nsew signal input
rlabel metal2 s 82726 165957 82782 166757 6 io_in[29]
port 150 nsew signal input
rlabel metal2 s 6090 165957 6146 166757 6 io_in[2]
port 151 nsew signal input
rlabel metal2 s 85578 165957 85634 166757 6 io_in[30]
port 152 nsew signal input
rlabel metal2 s 88430 165957 88486 166757 6 io_in[31]
port 153 nsew signal input
rlabel metal2 s 91282 165957 91338 166757 6 io_in[32]
port 154 nsew signal input
rlabel metal2 s 94042 165957 94098 166757 6 io_in[33]
port 155 nsew signal input
rlabel metal2 s 96894 165957 96950 166757 6 io_in[34]
port 156 nsew signal input
rlabel metal2 s 99746 165957 99802 166757 6 io_in[35]
port 157 nsew signal input
rlabel metal2 s 102598 165957 102654 166757 6 io_in[36]
port 158 nsew signal input
rlabel metal2 s 105450 165957 105506 166757 6 io_in[37]
port 159 nsew signal input
rlabel metal2 s 8942 165957 8998 166757 6 io_in[3]
port 160 nsew signal input
rlabel metal2 s 11794 165957 11850 166757 6 io_in[4]
port 161 nsew signal input
rlabel metal2 s 14646 165957 14702 166757 6 io_in[5]
port 162 nsew signal input
rlabel metal2 s 17498 165957 17554 166757 6 io_in[6]
port 163 nsew signal input
rlabel metal2 s 20258 165957 20314 166757 6 io_in[7]
port 164 nsew signal input
rlabel metal2 s 23110 165957 23166 166757 6 io_in[8]
port 165 nsew signal input
rlabel metal2 s 25962 165957 26018 166757 6 io_in[9]
port 166 nsew signal input
rlabel metal2 s 1398 165957 1454 166757 6 io_oeb[0]
port 167 nsew signal output
rlabel metal2 s 29734 165957 29790 166757 6 io_oeb[10]
port 168 nsew signal output
rlabel metal2 s 32586 165957 32642 166757 6 io_oeb[11]
port 169 nsew signal output
rlabel metal2 s 35438 165957 35494 166757 6 io_oeb[12]
port 170 nsew signal output
rlabel metal2 s 38290 165957 38346 166757 6 io_oeb[13]
port 171 nsew signal output
rlabel metal2 s 41142 165957 41198 166757 6 io_oeb[14]
port 172 nsew signal output
rlabel metal2 s 43902 165957 43958 166757 6 io_oeb[15]
port 173 nsew signal output
rlabel metal2 s 46754 165957 46810 166757 6 io_oeb[16]
port 174 nsew signal output
rlabel metal2 s 49606 165957 49662 166757 6 io_oeb[17]
port 175 nsew signal output
rlabel metal2 s 52458 165957 52514 166757 6 io_oeb[18]
port 176 nsew signal output
rlabel metal2 s 55310 165957 55366 166757 6 io_oeb[19]
port 177 nsew signal output
rlabel metal2 s 4250 165957 4306 166757 6 io_oeb[1]
port 178 nsew signal output
rlabel metal2 s 58162 165957 58218 166757 6 io_oeb[20]
port 179 nsew signal output
rlabel metal2 s 61014 165957 61070 166757 6 io_oeb[21]
port 180 nsew signal output
rlabel metal2 s 63774 165957 63830 166757 6 io_oeb[22]
port 181 nsew signal output
rlabel metal2 s 66626 165957 66682 166757 6 io_oeb[23]
port 182 nsew signal output
rlabel metal2 s 69478 165957 69534 166757 6 io_oeb[24]
port 183 nsew signal output
rlabel metal2 s 72330 165957 72386 166757 6 io_oeb[25]
port 184 nsew signal output
rlabel metal2 s 75182 165957 75238 166757 6 io_oeb[26]
port 185 nsew signal output
rlabel metal2 s 78034 165957 78090 166757 6 io_oeb[27]
port 186 nsew signal output
rlabel metal2 s 80794 165957 80850 166757 6 io_oeb[28]
port 187 nsew signal output
rlabel metal2 s 83646 165957 83702 166757 6 io_oeb[29]
port 188 nsew signal output
rlabel metal2 s 7010 165957 7066 166757 6 io_oeb[2]
port 189 nsew signal output
rlabel metal2 s 86498 165957 86554 166757 6 io_oeb[30]
port 190 nsew signal output
rlabel metal2 s 89350 165957 89406 166757 6 io_oeb[31]
port 191 nsew signal output
rlabel metal2 s 92202 165957 92258 166757 6 io_oeb[32]
port 192 nsew signal output
rlabel metal2 s 95054 165957 95110 166757 6 io_oeb[33]
port 193 nsew signal output
rlabel metal2 s 97906 165957 97962 166757 6 io_oeb[34]
port 194 nsew signal output
rlabel metal2 s 100666 165957 100722 166757 6 io_oeb[35]
port 195 nsew signal output
rlabel metal2 s 103518 165957 103574 166757 6 io_oeb[36]
port 196 nsew signal output
rlabel metal2 s 106370 165957 106426 166757 6 io_oeb[37]
port 197 nsew signal output
rlabel metal2 s 9862 165957 9918 166757 6 io_oeb[3]
port 198 nsew signal output
rlabel metal2 s 12714 165957 12770 166757 6 io_oeb[4]
port 199 nsew signal output
rlabel metal2 s 15566 165957 15622 166757 6 io_oeb[5]
port 200 nsew signal output
rlabel metal2 s 18418 165957 18474 166757 6 io_oeb[6]
port 201 nsew signal output
rlabel metal2 s 21270 165957 21326 166757 6 io_oeb[7]
port 202 nsew signal output
rlabel metal2 s 24122 165957 24178 166757 6 io_oeb[8]
port 203 nsew signal output
rlabel metal2 s 26882 165957 26938 166757 6 io_oeb[9]
port 204 nsew signal output
rlabel metal2 s 2318 165957 2374 166757 6 io_out[0]
port 205 nsew signal output
rlabel metal2 s 30746 165957 30802 166757 6 io_out[10]
port 206 nsew signal output
rlabel metal2 s 33506 165957 33562 166757 6 io_out[11]
port 207 nsew signal output
rlabel metal2 s 36358 165957 36414 166757 6 io_out[12]
port 208 nsew signal output
rlabel metal2 s 39210 165957 39266 166757 6 io_out[13]
port 209 nsew signal output
rlabel metal2 s 42062 165957 42118 166757 6 io_out[14]
port 210 nsew signal output
rlabel metal2 s 44914 165957 44970 166757 6 io_out[15]
port 211 nsew signal output
rlabel metal2 s 47766 165957 47822 166757 6 io_out[16]
port 212 nsew signal output
rlabel metal2 s 50526 165957 50582 166757 6 io_out[17]
port 213 nsew signal output
rlabel metal2 s 53378 165957 53434 166757 6 io_out[18]
port 214 nsew signal output
rlabel metal2 s 56230 165957 56286 166757 6 io_out[19]
port 215 nsew signal output
rlabel metal2 s 5170 165957 5226 166757 6 io_out[1]
port 216 nsew signal output
rlabel metal2 s 59082 165957 59138 166757 6 io_out[20]
port 217 nsew signal output
rlabel metal2 s 61934 165957 61990 166757 6 io_out[21]
port 218 nsew signal output
rlabel metal2 s 64786 165957 64842 166757 6 io_out[22]
port 219 nsew signal output
rlabel metal2 s 67546 165957 67602 166757 6 io_out[23]
port 220 nsew signal output
rlabel metal2 s 70398 165957 70454 166757 6 io_out[24]
port 221 nsew signal output
rlabel metal2 s 73250 165957 73306 166757 6 io_out[25]
port 222 nsew signal output
rlabel metal2 s 76102 165957 76158 166757 6 io_out[26]
port 223 nsew signal output
rlabel metal2 s 78954 165957 79010 166757 6 io_out[27]
port 224 nsew signal output
rlabel metal2 s 81806 165957 81862 166757 6 io_out[28]
port 225 nsew signal output
rlabel metal2 s 84658 165957 84714 166757 6 io_out[29]
port 226 nsew signal output
rlabel metal2 s 8022 165957 8078 166757 6 io_out[2]
port 227 nsew signal output
rlabel metal2 s 87418 165957 87474 166757 6 io_out[30]
port 228 nsew signal output
rlabel metal2 s 90270 165957 90326 166757 6 io_out[31]
port 229 nsew signal output
rlabel metal2 s 93122 165957 93178 166757 6 io_out[32]
port 230 nsew signal output
rlabel metal2 s 95974 165957 96030 166757 6 io_out[33]
port 231 nsew signal output
rlabel metal2 s 98826 165957 98882 166757 6 io_out[34]
port 232 nsew signal output
rlabel metal2 s 101678 165957 101734 166757 6 io_out[35]
port 233 nsew signal output
rlabel metal2 s 104438 165957 104494 166757 6 io_out[36]
port 234 nsew signal output
rlabel metal2 s 107290 165957 107346 166757 6 io_out[37]
port 235 nsew signal output
rlabel metal2 s 10874 165957 10930 166757 6 io_out[3]
port 236 nsew signal output
rlabel metal2 s 13634 165957 13690 166757 6 io_out[4]
port 237 nsew signal output
rlabel metal2 s 16486 165957 16542 166757 6 io_out[5]
port 238 nsew signal output
rlabel metal2 s 19338 165957 19394 166757 6 io_out[6]
port 239 nsew signal output
rlabel metal2 s 22190 165957 22246 166757 6 io_out[7]
port 240 nsew signal output
rlabel metal2 s 25042 165957 25098 166757 6 io_out[8]
port 241 nsew signal output
rlabel metal2 s 27894 165957 27950 166757 6 io_out[9]
port 242 nsew signal output
rlabel metal2 s 101862 0 101918 800 6 irq[0]
port 243 nsew signal output
rlabel metal2 s 102782 0 102838 800 6 irq[1]
port 244 nsew signal output
rlabel metal2 s 103794 0 103850 800 6 irq[2]
port 245 nsew signal output
rlabel metal2 s 105726 0 105782 800 6 o_addr1[0]
port 246 nsew signal output
rlabel metal2 s 110510 0 110566 800 6 o_addr1[1]
port 247 nsew signal output
rlabel metal3 s 163813 22040 164613 22160 6 o_addr1[2]
port 248 nsew signal output
rlabel metal3 s 163813 27208 164613 27328 6 o_addr1[3]
port 249 nsew signal output
rlabel metal3 s 163813 40264 164613 40384 6 o_addr1[4]
port 250 nsew signal output
rlabel metal2 s 122930 0 122986 800 6 o_addr1[5]
port 251 nsew signal output
rlabel metal3 s 0 59032 800 59152 6 o_addr1[6]
port 252 nsew signal output
rlabel metal2 s 128634 0 128690 800 6 o_addr1[7]
port 253 nsew signal output
rlabel metal2 s 130566 0 130622 800 6 o_addr1[8]
port 254 nsew signal output
rlabel metal3 s 0 13608 800 13728 6 o_addr1_1[0]
port 255 nsew signal output
rlabel metal3 s 163813 11568 164613 11688 6 o_addr1_1[1]
port 256 nsew signal output
rlabel metal2 s 112994 165957 113050 166757 6 o_addr1_1[2]
port 257 nsew signal output
rlabel metal2 s 116214 0 116270 800 6 o_addr1_1[3]
port 258 nsew signal output
rlabel metal2 s 118146 0 118202 800 6 o_addr1_1[4]
port 259 nsew signal output
rlabel metal2 s 121918 0 121974 800 6 o_addr1_1[5]
port 260 nsew signal output
rlabel metal3 s 0 56040 800 56160 6 o_addr1_1[6]
port 261 nsew signal output
rlabel metal3 s 0 74128 800 74248 6 o_addr1_1[7]
port 262 nsew signal output
rlabel metal3 s 0 80248 800 80368 6 o_addr1_1[8]
port 263 nsew signal output
rlabel metal3 s 0 1504 800 1624 6 o_csb0
port 264 nsew signal output
rlabel metal3 s 0 4496 800 4616 6 o_csb0_1
port 265 nsew signal output
rlabel metal3 s 0 7488 800 7608 6 o_csb1
port 266 nsew signal output
rlabel metal3 s 0 10480 800 10600 6 o_csb1_1
port 267 nsew signal output
rlabel metal2 s 106646 0 106702 800 6 o_din0[0]
port 268 nsew signal output
rlabel metal2 s 133418 0 133474 800 6 o_din0[10]
port 269 nsew signal output
rlabel metal2 s 132866 165957 132922 166757 6 o_din0[11]
port 270 nsew signal output
rlabel metal2 s 134706 165957 134762 166757 6 o_din0[12]
port 271 nsew signal output
rlabel metal3 s 163813 87184 164613 87304 6 o_din0[13]
port 272 nsew signal output
rlabel metal2 s 138570 165957 138626 166757 6 o_din0[14]
port 273 nsew signal output
rlabel metal2 s 140134 0 140190 800 6 o_din0[15]
port 274 nsew signal output
rlabel metal2 s 142342 165957 142398 166757 6 o_din0[16]
port 275 nsew signal output
rlabel metal2 s 142986 0 143042 800 6 o_din0[17]
port 276 nsew signal output
rlabel metal3 s 0 119688 800 119808 6 o_din0[18]
port 277 nsew signal output
rlabel metal2 s 148966 165957 149022 166757 6 o_din0[19]
port 278 nsew signal output
rlabel metal2 s 111062 165957 111118 166757 6 o_din0[1]
port 279 nsew signal output
rlabel metal2 s 146850 0 146906 800 6 o_din0[20]
port 280 nsew signal output
rlabel metal2 s 148782 0 148838 800 6 o_din0[21]
port 281 nsew signal output
rlabel metal2 s 152738 165957 152794 166757 6 o_din0[22]
port 282 nsew signal output
rlabel metal2 s 151634 0 151690 800 6 o_din0[23]
port 283 nsew signal output
rlabel metal2 s 158442 165957 158498 166757 6 o_din0[24]
port 284 nsew signal output
rlabel metal3 s 163813 139272 164613 139392 6 o_din0[25]
port 285 nsew signal output
rlabel metal3 s 163813 147024 164613 147144 6 o_din0[26]
port 286 nsew signal output
rlabel metal3 s 163813 152328 164613 152448 6 o_din0[27]
port 287 nsew signal output
rlabel metal2 s 158350 0 158406 800 6 o_din0[28]
port 288 nsew signal output
rlabel metal3 s 0 156000 800 156120 6 o_din0[29]
port 289 nsew signal output
rlabel metal2 s 114926 165957 114982 166757 6 o_din0[2]
port 290 nsew signal output
rlabel metal3 s 0 162120 800 162240 6 o_din0[30]
port 291 nsew signal output
rlabel metal2 s 164054 0 164110 800 6 o_din0[31]
port 292 nsew signal output
rlabel metal3 s 0 40808 800 40928 6 o_din0[3]
port 293 nsew signal output
rlabel metal2 s 120078 0 120134 800 6 o_din0[4]
port 294 nsew signal output
rlabel metal2 s 123390 165957 123446 166757 6 o_din0[5]
port 295 nsew signal output
rlabel metal3 s 0 65152 800 65272 6 o_din0[6]
port 296 nsew signal output
rlabel metal3 s 163813 55904 164613 56024 6 o_din0[7]
port 297 nsew signal output
rlabel metal3 s 163813 68960 164613 69080 6 o_din0[8]
port 298 nsew signal output
rlabel metal2 s 128174 165957 128230 166757 6 o_din0[9]
port 299 nsew signal output
rlabel metal2 s 107566 0 107622 800 6 o_din0_1[0]
port 300 nsew signal output
rlabel metal2 s 130934 165957 130990 166757 6 o_din0_1[10]
port 301 nsew signal output
rlabel metal2 s 135350 0 135406 800 6 o_din0_1[11]
port 302 nsew signal output
rlabel metal2 s 139214 0 139270 800 6 o_din0_1[12]
port 303 nsew signal output
rlabel metal3 s 163813 84600 164613 84720 6 o_din0_1[13]
port 304 nsew signal output
rlabel metal3 s 0 107584 800 107704 6 o_din0_1[14]
port 305 nsew signal output
rlabel metal3 s 163813 97520 164613 97640 6 o_din0_1[15]
port 306 nsew signal output
rlabel metal3 s 163813 102824 164613 102944 6 o_din0_1[16]
port 307 nsew signal output
rlabel metal2 s 143262 165957 143318 166757 6 o_din0_1[17]
port 308 nsew signal output
rlabel metal2 s 145194 165957 145250 166757 6 o_din0_1[18]
port 309 nsew signal output
rlabel metal3 s 163813 113160 164613 113280 6 o_din0_1[19]
port 310 nsew signal output
rlabel metal3 s 0 28704 800 28824 6 o_din0_1[1]
port 311 nsew signal output
rlabel metal2 s 145838 0 145894 800 6 o_din0_1[20]
port 312 nsew signal output
rlabel metal2 s 150806 165957 150862 166757 6 o_din0_1[21]
port 313 nsew signal output
rlabel metal2 s 150622 0 150678 800 6 o_din0_1[22]
port 314 nsew signal output
rlabel metal3 s 163813 123632 164613 123752 6 o_din0_1[23]
port 315 nsew signal output
rlabel metal2 s 157430 165957 157486 166757 6 o_din0_1[24]
port 316 nsew signal output
rlabel metal2 s 159362 165957 159418 166757 6 o_din0_1[25]
port 317 nsew signal output
rlabel metal3 s 163813 144440 164613 144560 6 o_din0_1[26]
port 318 nsew signal output
rlabel metal2 s 156418 0 156474 800 6 o_din0_1[27]
port 319 nsew signal output
rlabel metal2 s 157338 0 157394 800 6 o_din0_1[28]
port 320 nsew signal output
rlabel metal2 s 161202 0 161258 800 6 o_din0_1[29]
port 321 nsew signal output
rlabel metal2 s 113914 165957 113970 166757 6 o_din0_1[2]
port 322 nsew signal output
rlabel metal3 s 163813 162664 164613 162784 6 o_din0_1[30]
port 323 nsew signal output
rlabel metal3 s 163813 165248 164613 165368 6 o_din0_1[31]
port 324 nsew signal output
rlabel metal3 s 163813 29792 164613 29912 6 o_din0_1[3]
port 325 nsew signal output
rlabel metal2 s 119066 0 119122 800 6 o_din0_1[4]
port 326 nsew signal output
rlabel metal2 s 122470 165957 122526 166757 6 o_din0_1[5]
port 327 nsew signal output
rlabel metal3 s 0 62024 800 62144 6 o_din0_1[6]
port 328 nsew signal output
rlabel metal3 s 163813 53320 164613 53440 6 o_din0_1[7]
port 329 nsew signal output
rlabel metal3 s 163813 66240 164613 66360 6 o_din0_1[8]
port 330 nsew signal output
rlabel metal3 s 0 86368 800 86488 6 o_din0_1[9]
port 331 nsew signal output
rlabel metal2 s 109222 165957 109278 166757 6 o_waddr0[0]
port 332 nsew signal output
rlabel metal3 s 163813 14152 164613 14272 6 o_waddr0[1]
port 333 nsew signal output
rlabel metal3 s 163813 24624 164613 24744 6 o_waddr0[2]
port 334 nsew signal output
rlabel metal2 s 119618 165957 119674 166757 6 o_waddr0[3]
port 335 nsew signal output
rlabel metal2 s 120998 0 121054 800 6 o_waddr0[4]
port 336 nsew signal output
rlabel metal2 s 125322 165957 125378 166757 6 o_waddr0[5]
port 337 nsew signal output
rlabel metal3 s 0 68144 800 68264 6 o_waddr0[6]
port 338 nsew signal output
rlabel metal3 s 0 77256 800 77376 6 o_waddr0[7]
port 339 nsew signal output
rlabel metal3 s 0 83240 800 83360 6 o_waddr0[8]
port 340 nsew signal output
rlabel metal2 s 108578 0 108634 800 6 o_waddr0_1[0]
port 341 nsew signal output
rlabel metal2 s 112074 165957 112130 166757 6 o_waddr0_1[1]
port 342 nsew signal output
rlabel metal2 s 115846 165957 115902 166757 6 o_waddr0_1[2]
port 343 nsew signal output
rlabel metal2 s 118698 165957 118754 166757 6 o_waddr0_1[3]
port 344 nsew signal output
rlabel metal3 s 163813 42848 164613 42968 6 o_waddr0_1[4]
port 345 nsew signal output
rlabel metal2 s 124310 165957 124366 166757 6 o_waddr0_1[5]
port 346 nsew signal output
rlabel metal2 s 126702 0 126758 800 6 o_waddr0_1[6]
port 347 nsew signal output
rlabel metal3 s 163813 58488 164613 58608 6 o_waddr0_1[7]
port 348 nsew signal output
rlabel metal3 s 163813 71544 164613 71664 6 o_waddr0_1[8]
port 349 nsew signal output
rlabel metal3 s 163813 1232 164613 1352 6 o_web0
port 350 nsew signal output
rlabel metal3 s 163813 3816 164613 3936 6 o_web0_1
port 351 nsew signal output
rlabel metal3 s 0 16600 800 16720 6 o_wmask0[0]
port 352 nsew signal output
rlabel metal2 s 112350 0 112406 800 6 o_wmask0[1]
port 353 nsew signal output
rlabel metal2 s 116766 165957 116822 166757 6 o_wmask0[2]
port 354 nsew signal output
rlabel metal3 s 163813 32376 164613 32496 6 o_wmask0[3]
port 355 nsew signal output
rlabel metal3 s 0 19592 800 19712 6 o_wmask0_1[0]
port 356 nsew signal output
rlabel metal2 s 111430 0 111486 800 6 o_wmask0_1[1]
port 357 nsew signal output
rlabel metal3 s 0 31696 800 31816 6 o_wmask0_1[2]
port 358 nsew signal output
rlabel metal2 s 120538 165957 120594 166757 6 o_wmask0_1[3]
port 359 nsew signal output
rlabel metal4 s 4208 2128 4528 164336 6 vccd1
port 360 nsew power input
rlabel metal4 s 34928 2128 35248 164336 6 vccd1
port 360 nsew power input
rlabel metal4 s 65648 2128 65968 164336 6 vccd1
port 360 nsew power input
rlabel metal4 s 96368 2128 96688 164336 6 vccd1
port 360 nsew power input
rlabel metal4 s 127088 2128 127408 164336 6 vccd1
port 360 nsew power input
rlabel metal4 s 157808 2128 158128 164336 6 vccd1
port 360 nsew power input
rlabel metal4 s 19568 2128 19888 164336 6 vssd1
port 361 nsew ground input
rlabel metal4 s 50288 2128 50608 164336 6 vssd1
port 361 nsew ground input
rlabel metal4 s 81008 2128 81328 164336 6 vssd1
port 361 nsew ground input
rlabel metal4 s 111728 2128 112048 164336 6 vssd1
port 361 nsew ground input
rlabel metal4 s 142448 2128 142768 164336 6 vssd1
port 361 nsew ground input
rlabel metal2 s 478 0 534 800 6 wb_clk_i
port 362 nsew signal input
rlabel metal2 s 1398 0 1454 800 6 wb_rst_i
port 363 nsew signal input
rlabel metal2 s 2318 0 2374 800 6 wbs_ack_o
port 364 nsew signal output
rlabel metal2 s 6182 0 6238 800 6 wbs_adr_i[0]
port 365 nsew signal input
rlabel metal2 s 38750 0 38806 800 6 wbs_adr_i[10]
port 366 nsew signal input
rlabel metal2 s 41602 0 41658 800 6 wbs_adr_i[11]
port 367 nsew signal input
rlabel metal2 s 44454 0 44510 800 6 wbs_adr_i[12]
port 368 nsew signal input
rlabel metal2 s 47306 0 47362 800 6 wbs_adr_i[13]
port 369 nsew signal input
rlabel metal2 s 50158 0 50214 800 6 wbs_adr_i[14]
port 370 nsew signal input
rlabel metal2 s 53102 0 53158 800 6 wbs_adr_i[15]
port 371 nsew signal input
rlabel metal2 s 55954 0 56010 800 6 wbs_adr_i[16]
port 372 nsew signal input
rlabel metal2 s 58806 0 58862 800 6 wbs_adr_i[17]
port 373 nsew signal input
rlabel metal2 s 61658 0 61714 800 6 wbs_adr_i[18]
port 374 nsew signal input
rlabel metal2 s 64510 0 64566 800 6 wbs_adr_i[19]
port 375 nsew signal input
rlabel metal2 s 10046 0 10102 800 6 wbs_adr_i[1]
port 376 nsew signal input
rlabel metal2 s 67454 0 67510 800 6 wbs_adr_i[20]
port 377 nsew signal input
rlabel metal2 s 70306 0 70362 800 6 wbs_adr_i[21]
port 378 nsew signal input
rlabel metal2 s 73158 0 73214 800 6 wbs_adr_i[22]
port 379 nsew signal input
rlabel metal2 s 76010 0 76066 800 6 wbs_adr_i[23]
port 380 nsew signal input
rlabel metal2 s 78862 0 78918 800 6 wbs_adr_i[24]
port 381 nsew signal input
rlabel metal2 s 81806 0 81862 800 6 wbs_adr_i[25]
port 382 nsew signal input
rlabel metal2 s 84658 0 84714 800 6 wbs_adr_i[26]
port 383 nsew signal input
rlabel metal2 s 87510 0 87566 800 6 wbs_adr_i[27]
port 384 nsew signal input
rlabel metal2 s 90362 0 90418 800 6 wbs_adr_i[28]
port 385 nsew signal input
rlabel metal2 s 93214 0 93270 800 6 wbs_adr_i[29]
port 386 nsew signal input
rlabel metal2 s 13818 0 13874 800 6 wbs_adr_i[2]
port 387 nsew signal input
rlabel metal2 s 96158 0 96214 800 6 wbs_adr_i[30]
port 388 nsew signal input
rlabel metal2 s 99010 0 99066 800 6 wbs_adr_i[31]
port 389 nsew signal input
rlabel metal2 s 17682 0 17738 800 6 wbs_adr_i[3]
port 390 nsew signal input
rlabel metal2 s 21454 0 21510 800 6 wbs_adr_i[4]
port 391 nsew signal input
rlabel metal2 s 24398 0 24454 800 6 wbs_adr_i[5]
port 392 nsew signal input
rlabel metal2 s 27250 0 27306 800 6 wbs_adr_i[6]
port 393 nsew signal input
rlabel metal2 s 30102 0 30158 800 6 wbs_adr_i[7]
port 394 nsew signal input
rlabel metal2 s 32954 0 33010 800 6 wbs_adr_i[8]
port 395 nsew signal input
rlabel metal2 s 35806 0 35862 800 6 wbs_adr_i[9]
port 396 nsew signal input
rlabel metal2 s 3330 0 3386 800 6 wbs_cyc_i
port 397 nsew signal input
rlabel metal2 s 7102 0 7158 800 6 wbs_dat_i[0]
port 398 nsew signal input
rlabel metal2 s 39670 0 39726 800 6 wbs_dat_i[10]
port 399 nsew signal input
rlabel metal2 s 42522 0 42578 800 6 wbs_dat_i[11]
port 400 nsew signal input
rlabel metal2 s 45374 0 45430 800 6 wbs_dat_i[12]
port 401 nsew signal input
rlabel metal2 s 48318 0 48374 800 6 wbs_dat_i[13]
port 402 nsew signal input
rlabel metal2 s 51170 0 51226 800 6 wbs_dat_i[14]
port 403 nsew signal input
rlabel metal2 s 54022 0 54078 800 6 wbs_dat_i[15]
port 404 nsew signal input
rlabel metal2 s 56874 0 56930 800 6 wbs_dat_i[16]
port 405 nsew signal input
rlabel metal2 s 59726 0 59782 800 6 wbs_dat_i[17]
port 406 nsew signal input
rlabel metal2 s 62670 0 62726 800 6 wbs_dat_i[18]
port 407 nsew signal input
rlabel metal2 s 65522 0 65578 800 6 wbs_dat_i[19]
port 408 nsew signal input
rlabel metal2 s 10966 0 11022 800 6 wbs_dat_i[1]
port 409 nsew signal input
rlabel metal2 s 68374 0 68430 800 6 wbs_dat_i[20]
port 410 nsew signal input
rlabel metal2 s 71226 0 71282 800 6 wbs_dat_i[21]
port 411 nsew signal input
rlabel metal2 s 74078 0 74134 800 6 wbs_dat_i[22]
port 412 nsew signal input
rlabel metal2 s 77022 0 77078 800 6 wbs_dat_i[23]
port 413 nsew signal input
rlabel metal2 s 79874 0 79930 800 6 wbs_dat_i[24]
port 414 nsew signal input
rlabel metal2 s 82726 0 82782 800 6 wbs_dat_i[25]
port 415 nsew signal input
rlabel metal2 s 85578 0 85634 800 6 wbs_dat_i[26]
port 416 nsew signal input
rlabel metal2 s 88430 0 88486 800 6 wbs_dat_i[27]
port 417 nsew signal input
rlabel metal2 s 91374 0 91430 800 6 wbs_dat_i[28]
port 418 nsew signal input
rlabel metal2 s 94226 0 94282 800 6 wbs_dat_i[29]
port 419 nsew signal input
rlabel metal2 s 14830 0 14886 800 6 wbs_dat_i[2]
port 420 nsew signal input
rlabel metal2 s 97078 0 97134 800 6 wbs_dat_i[30]
port 421 nsew signal input
rlabel metal2 s 99930 0 99986 800 6 wbs_dat_i[31]
port 422 nsew signal input
rlabel metal2 s 18602 0 18658 800 6 wbs_dat_i[3]
port 423 nsew signal input
rlabel metal2 s 22466 0 22522 800 6 wbs_dat_i[4]
port 424 nsew signal input
rlabel metal2 s 25318 0 25374 800 6 wbs_dat_i[5]
port 425 nsew signal input
rlabel metal2 s 28170 0 28226 800 6 wbs_dat_i[6]
port 426 nsew signal input
rlabel metal2 s 31022 0 31078 800 6 wbs_dat_i[7]
port 427 nsew signal input
rlabel metal2 s 33966 0 34022 800 6 wbs_dat_i[8]
port 428 nsew signal input
rlabel metal2 s 36818 0 36874 800 6 wbs_dat_i[9]
port 429 nsew signal input
rlabel metal2 s 8114 0 8170 800 6 wbs_dat_o[0]
port 430 nsew signal output
rlabel metal2 s 40590 0 40646 800 6 wbs_dat_o[10]
port 431 nsew signal output
rlabel metal2 s 43534 0 43590 800 6 wbs_dat_o[11]
port 432 nsew signal output
rlabel metal2 s 46386 0 46442 800 6 wbs_dat_o[12]
port 433 nsew signal output
rlabel metal2 s 49238 0 49294 800 6 wbs_dat_o[13]
port 434 nsew signal output
rlabel metal2 s 52090 0 52146 800 6 wbs_dat_o[14]
port 435 nsew signal output
rlabel metal2 s 54942 0 54998 800 6 wbs_dat_o[15]
port 436 nsew signal output
rlabel metal2 s 57886 0 57942 800 6 wbs_dat_o[16]
port 437 nsew signal output
rlabel metal2 s 60738 0 60794 800 6 wbs_dat_o[17]
port 438 nsew signal output
rlabel metal2 s 63590 0 63646 800 6 wbs_dat_o[18]
port 439 nsew signal output
rlabel metal2 s 66442 0 66498 800 6 wbs_dat_o[19]
port 440 nsew signal output
rlabel metal2 s 11886 0 11942 800 6 wbs_dat_o[1]
port 441 nsew signal output
rlabel metal2 s 69294 0 69350 800 6 wbs_dat_o[20]
port 442 nsew signal output
rlabel metal2 s 72238 0 72294 800 6 wbs_dat_o[21]
port 443 nsew signal output
rlabel metal2 s 75090 0 75146 800 6 wbs_dat_o[22]
port 444 nsew signal output
rlabel metal2 s 77942 0 77998 800 6 wbs_dat_o[23]
port 445 nsew signal output
rlabel metal2 s 80794 0 80850 800 6 wbs_dat_o[24]
port 446 nsew signal output
rlabel metal2 s 83646 0 83702 800 6 wbs_dat_o[25]
port 447 nsew signal output
rlabel metal2 s 86590 0 86646 800 6 wbs_dat_o[26]
port 448 nsew signal output
rlabel metal2 s 89442 0 89498 800 6 wbs_dat_o[27]
port 449 nsew signal output
rlabel metal2 s 92294 0 92350 800 6 wbs_dat_o[28]
port 450 nsew signal output
rlabel metal2 s 95146 0 95202 800 6 wbs_dat_o[29]
port 451 nsew signal output
rlabel metal2 s 15750 0 15806 800 6 wbs_dat_o[2]
port 452 nsew signal output
rlabel metal2 s 97998 0 98054 800 6 wbs_dat_o[30]
port 453 nsew signal output
rlabel metal2 s 100942 0 100998 800 6 wbs_dat_o[31]
port 454 nsew signal output
rlabel metal2 s 19614 0 19670 800 6 wbs_dat_o[3]
port 455 nsew signal output
rlabel metal2 s 23386 0 23442 800 6 wbs_dat_o[4]
port 456 nsew signal output
rlabel metal2 s 26238 0 26294 800 6 wbs_dat_o[5]
port 457 nsew signal output
rlabel metal2 s 29182 0 29238 800 6 wbs_dat_o[6]
port 458 nsew signal output
rlabel metal2 s 32034 0 32090 800 6 wbs_dat_o[7]
port 459 nsew signal output
rlabel metal2 s 34886 0 34942 800 6 wbs_dat_o[8]
port 460 nsew signal output
rlabel metal2 s 37738 0 37794 800 6 wbs_dat_o[9]
port 461 nsew signal output
rlabel metal2 s 9034 0 9090 800 6 wbs_sel_i[0]
port 462 nsew signal input
rlabel metal2 s 12898 0 12954 800 6 wbs_sel_i[1]
port 463 nsew signal input
rlabel metal2 s 16670 0 16726 800 6 wbs_sel_i[2]
port 464 nsew signal input
rlabel metal2 s 20534 0 20590 800 6 wbs_sel_i[3]
port 465 nsew signal input
rlabel metal2 s 4250 0 4306 800 6 wbs_stb_i
port 466 nsew signal input
rlabel metal2 s 5262 0 5318 800 6 wbs_we_i
port 467 nsew signal input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 164613 166757
string LEFview TRUE
string GDS_FILE /local/caravel_user_project/openlane/user_proj/runs/user_proj/results/magic/user_proj.gds
string GDS_END 80477832
string GDS_START 1360530
<< end >>

